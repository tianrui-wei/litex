
 
 
 
 
 
 
 
module network_input_blk_multi_out 
   #(parameter LOG2_NUMBER_FIFO_ELEMENTS = 2)
(
   input wire clk, 
   input wire reset,
   input wire [64-1:0] data_in, 
   input wire valid_in, 
   input wire thanks_in,
   output wire yummy_out, 
   
   
   output wire [64-1:0] data_val, 
   output wire [64-1:0] data_val1, 
   output wire data_avail 
);
reg [64-1:0] storage_data_f [0:(1<<LOG2_NUMBER_FIFO_ELEMENTS)-1];
reg [LOG2_NUMBER_FIFO_ELEMENTS-1:0] head_ptr_f;
reg [LOG2_NUMBER_FIFO_ELEMENTS-1:0] tail_ptr_f;
reg [LOG2_NUMBER_FIFO_ELEMENTS:0] elements_in_array_f;
reg [LOG2_NUMBER_FIFO_ELEMENTS-1:0] head_ptr_next;
reg [LOG2_NUMBER_FIFO_ELEMENTS-1:0] tail_ptr_next;
reg [LOG2_NUMBER_FIFO_ELEMENTS:0] elements_in_array_next;
reg yummy_out_f;
assign yummy_out = yummy_out_f;
assign data_val = storage_data_f[head_ptr_f];
assign data_val1 = storage_data_f[head_ptr_f];
assign data_avail = elements_in_array_f != 0;
always @ *
begin
   head_ptr_next = head_ptr_f;
   tail_ptr_next = tail_ptr_f;
   elements_in_array_next = elements_in_array_f;
   case({valid_in,thanks_in})
      2'b00:
         begin
            
         end
      2'b01:
         begin
            
            head_ptr_next = head_ptr_f + 1;
            elements_in_array_next = elements_in_array_f - 1;
         end
      2'b10:
         begin
            
            tail_ptr_next = tail_ptr_f + 1;
            elements_in_array_next = elements_in_array_f + 1;
         end
      2'b11:
         begin
            
            head_ptr_next = head_ptr_f + 1;
            tail_ptr_next = tail_ptr_f + 1;
         end
      default:
         begin
            
         end
   endcase
end
always @ (posedge clk)
begin
   if (reset)
   begin
      yummy_out_f <= 0;
      head_ptr_f <= 0;
      tail_ptr_f <= 0;
      elements_in_array_f <= 0;
   end
   else
   begin
      yummy_out_f <= thanks_in; 
      head_ptr_f <= head_ptr_next;
      tail_ptr_f <= tail_ptr_next;
      elements_in_array_f <= elements_in_array_next;
      if(valid_in)
      begin
         storage_data_f[tail_ptr_f] <= data_in;
      end
   end
end
endmodule
module space_avail_top (valid,
		    yummy,
		    spc_avail,
		    clk,
		    reset);
parameter BUFFER_SIZE = 4;
parameter BUFFER_BITS = 3;
   
 
input valid;			
input yummy;			
output spc_avail;		
input clk;
input reset;
reg yummy_f;
reg valid_f;
reg [BUFFER_BITS-1:0] count_f;
reg is_one_f;
reg is_two_or_more_f;
wire [BUFFER_BITS-1:0] count_plus_1;
wire [BUFFER_BITS-1:0] count_minus_1;
wire up;
wire down;
reg [BUFFER_BITS-1:0] count_temp;
assign count_plus_1 = count_f + 1'b1;
assign count_minus_1 = count_f - 1'b1;
assign spc_avail = (is_two_or_more_f | yummy_f | (is_one_f & ~valid_f));
assign up = yummy_f & ~valid_f;
assign down = ~yummy_f & valid_f;
always @ (count_f or count_plus_1 or count_minus_1 or up or down)
begin
	case (count_f)
	0:
		begin
			if(up)
			begin
				count_temp <= count_plus_1;
			end
			else
			begin
				count_temp <= count_f;
			end
		end
	BUFFER_SIZE:
		begin
			if(down)
			begin
				count_temp <= count_minus_1;
			end
			else
			begin
				count_temp <= count_f;
			end
		end
	default:
		begin
			case ({up, down})
				2'b10:	count_temp <= count_plus_1;
				2'b01:	count_temp <= count_minus_1;
				default:	count_temp <= count_f;
			endcase
		end
	endcase
end
wire top_bits_zero_temp = ~| count_temp[BUFFER_BITS-1:1];
always @ (posedge clk)
begin
	if(reset)
	begin
	   count_f <= BUFFER_SIZE;
	   yummy_f <= 1'b0;
	   valid_f <= 1'b0;
	   is_one_f <= (BUFFER_SIZE == 1);
	   is_two_or_more_f <= (BUFFER_SIZE >= 2);
	end
	else
	begin
	   count_f <= count_temp;
	   yummy_f <= yummy;
	   valid_f <= valid;
	   is_one_f         <= top_bits_zero_temp & count_temp[0];
   	   is_two_or_more_f <= ~top_bits_zero_temp;
	end
end
endmodule
      
module bram_map #(parameter MEM_ADDR_WIDTH=64, PHY_ADDR_WIDTH=40, BRAM_ADDR_WIDTH=12)
(
    input       [PHY_ADDR_WIDTH-1:0]    msg_addr,
    
    output      [BRAM_ADDR_WIDTH-1:0]   bram_blk_addr,
    output                              hit_any_section
);
assign bram_blk_addr = {BRAM_ADDR_WIDTH{1'b0}};
assign hit_any_section = 0;
endmodule
 
 
 
 
 
 
 
 
 
  
module ciop_iob (
    input                               chip_clk,
    input                               fpga_clk,
    input                               rst_n,
    
                     
    input                               noc1_in_val,
    input [64-1:0]         noc1_in_data,
    output reg                          noc1_in_rdy,
    output                              noc2_out_val,
    output reg [64-1:0]        noc2_out_data,
    input                               noc2_out_rdy,
    input                               noc3_in_val,
    input [64-1:0]         noc3_in_data,
    output wire                         noc3_in_rdy,
    input                               noc2_in_val,
    input [64-1:0]         noc2_in_data,
    output reg                          noc2_in_rdy,
    output                              noc3_out_val,
    output [64-1:0]        noc3_out_data,
    input                               noc3_out_rdy,
    input                               uart_interrupt,
    input                               net_interrupt
);
   parameter OK_IOB_CNT = 40000; 
wire                    ok_iob;
reg     [31:0]          ok_iob_cnt;
assign noc3_in_rdy = 1'b1;
assign  ok_iob = ok_iob_cnt == OK_IOB_CNT;
always @(posedge chip_clk) begin
    if (~rst_n)
        ok_iob_cnt <= 32'b0;
    else
        ok_iob_cnt <= ok_iob ? ok_iob_cnt : ok_iob_cnt + 1'b1 ;
end
parameter FLIT_TO_SEND = 2;
wire [63:0]         iob_buffer_flit1;
wire [63:0]         iob_buffer_flit2;
reg                 iob_buffer_val;
reg  [1:0]          flit_cnt;
reg  [1:0]          net_flit_cnt;
reg  [1:0]          uart_flit_cnt;
assign iob_buffer_flit1     = 64'h0000_0000_0048_4000;
assign iob_buffer_flit2     = 64'h0000_0000_0001_0001;
reg                 ok_iob_sent;
wire [63:0]         iob_buffer_net_flit2;
reg                 pending_net_interrupt;
reg                 net_interrupt_in_prog;
reg                 prev_net_interrupt;
reg                 buf_prev_net_int;
   
wire [63:0]         iob_buffer_uart_flit2;
reg                 pending_uart_interrupt;
reg                 uart_interrupt_in_prog;
reg                 prev_uart_interrupt;
reg                 buf_prev_uart_int;
   
assign iob_buffer_net_flit2 = 64'h0000_0000_0000_001d;
assign iob_buffer_uart_flit2 = 64'h0000_0000_0000_001c;
   
always @(posedge fpga_clk) begin
    if (~rst_n) begin
        flit_cnt <= 2'b0;
        
        net_flit_cnt <= 2'b0;
        pending_net_interrupt <= 1'b0;
        net_interrupt_in_prog <= 1'b0;
        
        uart_flit_cnt <= 2'b0;
        pending_uart_interrupt <= 1'b0;
        uart_interrupt_in_prog <= 1'b0;
    end
    else if (~ok_iob_sent) begin
        flit_cnt <= noc2_out_val & noc2_out_rdy ? flit_cnt + 1 : flit_cnt;
    end 
    else begin
        flit_cnt <= flit_cnt;
     
     
    end
end
   
always @(posedge fpga_clk) begin
    if (~rst_n) begin
       prev_net_interrupt <= 1'b0;
       buf_prev_net_int <= 1'b0;
       prev_uart_interrupt <= 1'b0;
       buf_prev_uart_int <= 1'b0;
       iob_buffer_val = 1'b0;
    end
    else begin
       prev_net_interrupt <= net_interrupt;
       buf_prev_net_int <= prev_net_interrupt;
       prev_uart_interrupt <= uart_interrupt;
       buf_prev_uart_int <= prev_uart_interrupt;
       iob_buffer_val <= ok_iob;
    end
end
assign noc2_out_val = iob_buffer_val & (((flit_cnt < FLIT_TO_SEND) && !ok_iob_sent)
                    );
always @(*) begin
    if (!ok_iob_sent) begin
        if(flit_cnt == 2'b0) begin
            noc2_out_data = iob_buffer_flit1;
        end else if (flit_cnt == 2'b1) begin
            noc2_out_data = iob_buffer_flit2;
        end 
        else begin
            noc2_out_data =  {64{1'b0}};
        end
    end 
    else begin
        noc2_out_data =  {64{1'b0}};
    end
end
always @(posedge fpga_clk) begin
    if (~rst_n) begin
        ok_iob_sent <= 1'b0;
    end
    else if (flit_cnt == FLIT_TO_SEND) begin
       ok_iob_sent <= 1'b1;
    end
end
assign noc3_out_val     = 1'b0;
assign noc3_out_data    = {64{1'b0}};
endmodule
module eth_top #(
  parameter SWAP_ENDIANESS = 0
) (
    input                                   chipset_clk,
    input                                   rst_n,
    output                                  net_interrupt,
    input                                   noc_in_val,
    input       [64-1:0]       noc_in_data,
    output                                  noc_in_rdy,
    output                                  noc_out_val,
    output      [64-1:0]       noc_out_data,
    input                                   noc_out_rdy,
    input                                   net_axi_clk,
    output                                  net_phy_rst_n,
    input                                   net_phy_tx_clk,
    output                                  net_phy_tx_en,
    output  [3 : 0]                         net_phy_tx_data,
    input                                   net_phy_rx_clk,
    input                                   net_phy_dv,
    input  [3 : 0]                          net_phy_rx_data,
    input                                   net_phy_rx_er,
    inout                                   net_phy_mdio_io,
    output                                  net_phy_mdc
);
   
    assign noc_in_rdy    = 1'b0;
    assign noc_out_val    = 1'b0;
    assign noc_out_data   = {64{1'b0}};
    assign net_phy_tx_en        = 1'b0;
    assign net_phy_mdc          = 1'b0;
  
endmodule
      
 
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
   
    
   
    
       
        
        
    
  
   
     
    
   
   
    
    
module fake_boot_ctrl(
    input wire clk,
    input wire rst_n,
    input wire noc_valid_in,
    input wire [64-1:0] noc_data_in,
    output reg noc_ready_in,
    output reg noc_valid_out,
    output reg [64-1:0] noc_data_out,
    input wire noc_ready_out
);
reg mem_valid_in;
reg [3*64-1:0] mem_header_in;
reg mem_ready_in;
reg [64-1:0] buf_in_mem_f [10:0];
reg [64-1:0] buf_in_mem_next;
reg [8-1:0] buf_in_counter_f;
reg [8-1:0] buf_in_counter_next;
reg [3:0] buf_in_wr_ptr_f;
reg [3:0] buf_in_wr_ptr_next;
always @ *
begin
    noc_ready_in = (buf_in_counter_f == 0) || (buf_in_counter_f < (buf_in_mem_f[0][29:22]+1));
end
always @ *
begin
    if (noc_valid_in && noc_ready_in)
    begin
        buf_in_counter_next = buf_in_counter_f + 1;
    end
    else if (mem_valid_in && mem_ready_in)
    begin
        buf_in_counter_next = 0;
    end
    else
    begin
        buf_in_counter_next = buf_in_counter_f;
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        buf_in_counter_f <= 0;
    end
    else
    begin
        buf_in_counter_f <= buf_in_counter_next;
    end
end
always @ *
begin
    if (mem_valid_in && mem_ready_in)
    begin
        buf_in_wr_ptr_next = 0;
    end
    else if (noc_valid_in && noc_ready_in)
    begin
        buf_in_wr_ptr_next = buf_in_wr_ptr_f + 1;
    end
    else
    begin
        buf_in_wr_ptr_next = buf_in_wr_ptr_f;
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        buf_in_wr_ptr_f <= 0;
    end
    else
    begin
        buf_in_wr_ptr_f <= buf_in_wr_ptr_next;
    end
end
always @ *
begin
    if (noc_valid_in && noc_ready_in)
    begin
        buf_in_mem_next = noc_data_in;
    end
    else
    begin
        buf_in_mem_next = buf_in_mem_f[buf_in_wr_ptr_f];
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        buf_in_mem_f[buf_in_wr_ptr_f] <= 0;
    end
    else
    begin
        buf_in_mem_f[buf_in_wr_ptr_f] <= buf_in_mem_next;
    end
end
always @ *
begin
    mem_valid_in = (buf_in_counter_f != 0) && (buf_in_counter_f == (buf_in_mem_f[0][29:22]+1));
end
always @ *
begin
    mem_header_in = {buf_in_mem_f[2], buf_in_mem_f[1], buf_in_mem_f[0]};
end
wire [8-1:0] msg_type;
wire [8-1:0] msg_mshrid;
wire [3-1:0] msg_data_size;
wire [40-1:0] msg_addr;
wire [14-1:0] msg_src_chipid;
wire [8-1:0] msg_src_x;
wire [8-1:0] msg_src_y;
wire [4-1:0] msg_src_fbits;
reg [64-1:0] msg_send_data [7:0];
reg [64-1:0] mem_temp;
wire [64*3-1:0] msg_send_header;
wire    bram_ce;
wire    bram_rdwen;
l2_decoder decoder(
    .msg_header         (mem_header_in),
    .msg_type           (msg_type),
    .msg_length         (),
    .msg_mshrid         (msg_mshrid),
    .msg_data_size      (msg_data_size),
    .msg_cache_type     (),
    .msg_subline_vector (),
    .msg_mesi           (),
    .msg_l2_miss        (),
    .msg_subline_id     (),
    .msg_last_subline   (),
    .msg_addr           (msg_addr),
    .msg_src_chipid     (msg_src_chipid),
    .msg_src_x          (msg_src_x),
    .msg_src_y          (msg_src_y),
    .msg_src_fbits      (msg_src_fbits),
    .msg_sdid           (),
    .msg_lsid           ()
);
reg [63:0] write_mask;
always @ *
begin
    if (msg_data_size == 3'b001)
    begin
        write_mask = 64'hff00000000000000;
        write_mask = write_mask >> (8*msg_addr[2:0]);
    end
    else if (msg_data_size == 3'b010)
    begin
        write_mask = 64'hffff000000000000;
        write_mask = write_mask >> (16*msg_addr[2:1]);
    end
    else if (msg_data_size == 3'b011)
    begin
        write_mask = 64'hffffffff00000000;
        write_mask = write_mask >> (32*msg_addr[2]);
    end
    else if (msg_data_size == 3'b100)
    begin
        write_mask = 64'hffffffffffffffff;
    end
    else
    begin
        write_mask = 64'h0000000000000000;
    end
end
localparam BRAM_ADDR_WIDTH  =   clogb2(16384);
wire                            bram_r_val;
wire                            bram_r_val_hit;
wire [512-1:0]      bram_data_out;
wire                            bram_w_val;
wire                            bram_w_val_hit;
wire [512-1:0]      bram_w_mask;
wire [512-1:0]      bram_data_in;
wire [BRAM_ADDR_WIDTH-1:0]      bram_addr;    
wire [BRAM_ADDR_WIDTH-1+3:0]    translated_addr; 
wire [64-1:0]      buf_out_mem [8:0];
reg  [64*3-1:0]    msg_send_header_r;
wire [8-1:0]      msg_send_type;
wire [8-1:0]    msg_send_length;
reg  [2-1:0] addr_subline_r;
wire                            hit_bram;
reg                             hit_bram_r;
wire [512-1:0]      read_data;
reg  [64-1:0]      buf_out_mem_r [8:0];
wire                            mem_process_next_val;
reg                             mem_process_next_val_r;
    storage_addr_trans #(
        .STORAGE_ADDR_WIDTH (BRAM_ADDR_WIDTH)
    ) storage_addr_trans (
        .va_byte_addr       (msg_addr       ),
        .storage_addr_out   (translated_addr),
        .hit_any_section    (hit_bram       )
    );
assign bram_addr = translated_addr[BRAM_ADDR_WIDTH-1+3:3];
assign mem_process_next_val = mem_valid_in & mem_ready_in;
assign read_data = hit_bram_r ? bram_data_out : {512{1'b0}};
assign bram_r_val       = mem_valid_in & ((msg_type == 8'd19) | (msg_type == 8'd14));
assign buf_out_mem[0]   = mem_process_next_val_r  ? msg_send_header_r[64-1:0] : buf_out_mem_r[0];
assign {buf_out_mem[8], buf_out_mem[7], buf_out_mem[6], buf_out_mem[5],
        buf_out_mem[4], buf_out_mem[3]}     = mem_process_next_val_r ? read_data[511:128] : 
                                              {buf_out_mem_r[8], buf_out_mem_r[7], buf_out_mem_r[6], buf_out_mem_r[5],
                                               buf_out_mem_r[4], buf_out_mem_r[3]};
assign {buf_out_mem[2], buf_out_mem[1]}     = mem_process_next_val_r ? 
                                             (addr_subline_r == 2'b00 ? read_data[127:0]    :
                                              addr_subline_r == 2'b01 ? read_data[255:128]  :
                                              addr_subline_r == 2'b10 ? read_data[383:256]  : read_data[511:384]) :
                                             {buf_out_mem_r[2], buf_out_mem_r[1]};
assign bram_w_val       = mem_valid_in & ((msg_type == 8'd20) | (msg_type == 8'd15));
assign bram_data_in     = {buf_in_mem_f[10], buf_in_mem_f[9], buf_in_mem_f[8], buf_in_mem_f[7], 
                           buf_in_mem_f[6],  buf_in_mem_f[5], buf_in_mem_f[4], buf_in_mem_f[3]};
assign bram_w_mask      = msg_type == 8'd15 ? write_mask <<  64*(1<<msg_addr[5:3]) : {512{1'b1}};
assign msg_send_type    = {8{mem_valid_in}} &
                         (msg_type == 8'd19        ? 8'd24        :
                          msg_type == 8'd20       ? 8'd25       :
                          msg_type == 8'd14     ? 8'd26     :
                          msg_type == 8'd15    ? 8'd27    : 8'd30);
assign msg_send_length  = {8{1'b1}} & 
                         (msg_type == 8'd19        ? 8'd8  :
                          msg_type == 8'd20       ? 8'd0  :
                          msg_type == 8'd14     ? 8'd2  :
                          msg_type == 8'd15    ? 8'd0  : 8'd0);
always @(posedge clk)
    msg_send_header_r <= msg_send_header;
always @(posedge clk)
    addr_subline_r <= msg_type == 8'd14 ? msg_addr[5:4] : 2'b0;
always @(posedge clk)
    hit_bram_r <= hit_bram;
always @(posedge clk)
    mem_process_next_val_r <= mem_process_next_val;
always @(posedge clk) begin
    buf_out_mem_r[8] <= buf_out_mem[8];
    buf_out_mem_r[7] <= buf_out_mem[7];
    buf_out_mem_r[6] <= buf_out_mem[6];
    buf_out_mem_r[5] <= buf_out_mem[5];
    buf_out_mem_r[4] <= buf_out_mem[4];
    buf_out_mem_r[3] <= buf_out_mem[3];
    buf_out_mem_r[2] <= buf_out_mem[2];
    buf_out_mem_r[1] <= buf_out_mem[1];
    buf_out_mem_r[0] <= buf_out_mem[0];
end
assign bram_r_val_hit = bram_r_val & hit_bram_r;
assign bram_w_val_hit = bram_w_val & hit_bram_r;
assign bram_ce      = bram_r_val_hit | bram_w_val_hit;
assign bram_rdwen   = bram_r_val_hit;
bram_sdp_wrapper #(
    .NAME           ("bram_boot"                    ),
    .DEPTH          (256         ),
    .ADDR_WIDTH     (8    ),
    .BITMASK_WIDTH  (512    ),
    .DATA_WIDTH     (512    )
) bram (
    .MEMCLK         (clk            ),
    .A              (bram_addr      ),
    .CE             (bram_ce        ),
    .RDWEN          (bram_rdwen     ),
    .BW             (bram_w_mask    ),
    .DIN            (bram_data_in   ),
    .DOUT           (bram_data_out  )
);
l2_encoder encoder(
    .msg_dst_chipid             (msg_src_chipid),
    .msg_dst_x                  (msg_src_x),
    .msg_dst_y                  (msg_src_y),
    .msg_dst_fbits              (msg_src_fbits),
    .msg_length                 (msg_send_length),
    .msg_type                   (msg_send_type),
    .msg_mshrid                 (msg_mshrid),
    .msg_data_size              ({3{1'b0}}),
    .msg_cache_type             ({1{1'b0}}),
    .msg_subline_vector         ({4{1'b0}}),
    .msg_mesi                   ({2{1'b0}}),
    .msg_l2_miss                (msg_addr[40-1]),
    .msg_subline_id             ({2{1'b0}}),
    .msg_last_subline           ({1{1'b1}}),
    .msg_addr                   (msg_addr),
    .msg_src_chipid             ({14{1'b0}}),
    .msg_src_x                  ({8{1'b0}}),
    .msg_src_y                  ({8{1'b0}}),
    .msg_src_fbits              ({4{1'b0}}),
    .msg_sdid                   ({10{1'b0}}),
    .msg_lsid                   ({6{1'b0}}),
    .msg_header                 (msg_send_header)
);
reg [8-1:0] buf_out_counter_f;
reg [8-1:0] buf_out_counter_next;
reg [3:0] buf_out_rd_ptr_f;
reg [3:0] buf_out_rd_ptr_next;
always @ *
begin
    noc_valid_out = (buf_out_counter_f != 0);
end
always @ *
begin
    mem_ready_in = (buf_out_counter_f == 0);
end
always @ *
begin
    if (noc_valid_out && noc_ready_out)
    begin
        buf_out_counter_next = buf_out_counter_f - 1;
    end
    else if (mem_valid_in && mem_ready_in)
    begin
        buf_out_counter_next = msg_send_length + 1;
    end
    else
    begin
        buf_out_counter_next = buf_out_counter_f;
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        buf_out_counter_f <= 0;
    end
    else
    begin
        buf_out_counter_f <= buf_out_counter_next;
    end
end
always @ *
begin
    if (mem_valid_in && mem_ready_in)
    begin
        buf_out_rd_ptr_next = 0;
    end
    else if (noc_valid_out && noc_ready_out)
    begin
        buf_out_rd_ptr_next = buf_out_rd_ptr_f + 1;
    end
    else
    begin
        buf_out_rd_ptr_next = buf_out_rd_ptr_f;
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        buf_out_rd_ptr_f <= 0;
    end
    else
    begin
        buf_out_rd_ptr_f <= buf_out_rd_ptr_next;
    end
end
always @ *
begin
    noc_valid_out = (buf_out_counter_f != 0);
end
always @ *
begin
    
    noc_data_out = 0;
    if (buf_out_rd_ptr_f < 9)
        noc_data_out = buf_out_mem[buf_out_rd_ptr_f];
end
function integer clogb2;
  input [31:0] value;
  begin
    value = value - 1;
    for (clogb2 = 0; value > 0; clogb2 = clogb2 + 1) begin
      value = value >> 1;
    end
  end
endfunction
endmodule
module net_int_sync (
input clk_emac,
input clk_ciop,
input rst_n,
input net_int,
(* ASYNC_REG = "TRUE" *) output reg sync_int);
(* ASYNC_REG = "TRUE" *) reg int_buffer_ff;
(* ASYNC_REG = "TRUE" *) reg ack_buffer_ff;
(* ASYNC_REG = "TRUE" *) reg sync_ack;
(* ASYNC_REG = "TRUE" *) reg store_int;
   
always @(posedge clk_emac or posedge net_int) begin
    if (~rst_n) begin
        store_int <= 1'b0;
    end
    
    else if (net_int) begin
        store_int <= 1'b1;
    end
    
    else if (sync_ack) begin
        store_int <= 1'b0;
    end
end
always @(posedge clk_ciop) begin
    if (~rst_n) begin
        int_buffer_ff <= 1'b0;
        sync_int <= 1'b0;
    end
    else begin
        int_buffer_ff <= store_int;
        sync_int <= int_buffer_ff;
    end
end
always @(posedge clk_emac) begin
    if (~rst_n) begin
        ack_buffer_ff <= 1'b0;
        sync_ack <= 1'b0;
    end
    else begin
        ack_buffer_ff <= sync_int;
        sync_ack <= ack_buffer_ff;
    end
end
endmodule
         
         
   
    
   
    
       
        
        
    
  
   
     
    
   
   
    
    
module uart_mux (
    input               axi_clk,
    input               axi_rst_n,
    input               uart_boot_en,
    input               uart_timeout_en,
    input               init_done,
    
    output              writer_start,
    input               writer_finish,
    output  reg [2:0]   writer_str_sel,
    output              reader_start,
    input               reader_stop,
    output              test_start,
    input               test_good_end,
    input               test_bad_end,
    
    input   [12:0]      init_axi_awaddr, 
    input               init_axi_awvalid,
    output              init_axi_awready,
    input   [31:0]      init_axi_wdata,  
    input   [3:0 ]      init_axi_wstrb,  
    input               init_axi_wvalid, 
    output              init_axi_wready, 
    output  [1:0]       init_axi_bresp,  
    output              init_axi_bvalid, 
    input               init_axi_bready,
    
    input   [12:0]      writer_axi_awaddr,
    input               writer_axi_awvalid,
    output              writer_axi_awready,
    input   [31:0]      writer_axi_wdata,
    input   [3:0]       writer_axi_wstrb,
    input               writer_axi_wvalid,
    output              writer_axi_wready,
    output  [1:0]       writer_axi_bresp,
    output              writer_axi_bvalid,
    input               writer_axi_bready,
    input   [31:0]      writer_axi_araddr,
    input               writer_axi_arvalid,
    output              writer_axi_arready,
    output  [31:0]      writer_axi_rdata,
    output  [1:0]       writer_axi_rresp,
    output              writer_axi_rvalid,
    input               writer_axi_rready,
    
    input   [12:0]      core_axi_awaddr,
    input               core_axi_awvalid,
    output              core_axi_awready,
    input   [31:0]      core_axi_wdata,
    input   [3:0]       core_axi_wstrb,
    input               core_axi_wvalid,
    output              core_axi_wready,
    output  [1:0]       core_axi_bresp,
    output              core_axi_bvalid,
    input               core_axi_bready,
    input   [31:0]      core_axi_araddr,
    input               core_axi_arvalid,
    output              core_axi_arready,
    output  [31:0]      core_axi_rdata,
    output  [1:0]       core_axi_rresp,
    output              core_axi_rvalid,
    input               core_axi_rready,
    
    input   [31:0]      reader_axi_araddr,
    input               reader_axi_arvalid,
    output              reader_axi_arready,
    output  [31:0]      reader_axi_rdata,
    output  [1:0]       reader_axi_rresp,
    output              reader_axi_rvalid,
    input               reader_axi_rready,
    
    output   reg    [12:0]  s_axi_awaddr,
    output   reg            s_axi_awvalid,
    input                   s_axi_awready,
    output   reg    [31:0]  s_axi_wdata,
    output   reg    [3:0 ]  s_axi_wstrb,
    output   reg            s_axi_wvalid,
    input                   s_axi_wready,
    input           [1:0]   s_axi_bresp,
    input                   s_axi_bvalid,
    output   reg            s_axi_bready,
    output   reg    [12:0]  s_axi_araddr,
    output   reg            s_axi_arvalid,
    input                   s_axi_arready,
    input           [31:0]  s_axi_rdata,
    input           [1:0]   s_axi_rresp,
    input                   s_axi_rvalid,
    output   reg            s_axi_rready
);
localparam INIT_SEL         = 0;
localparam WRITER_SEL       = 1;
localparam READER_SEL       = 2;
localparam TEST_SEL         = 3;
wire [2:0]  mux_sel_rst_state;
wire        asm_test_timeout;
wire                    pc_good_trap;
wire                    pc_bad_trap;
reg     [2:0]       mux_sel;
reg     [63:0]      asm_test_cycle_cnt;
reg                 uart_boot_en_ff;
reg                 uart_timeout_en_ff;
always @(posedge axi_clk) begin
    uart_boot_en_ff <= uart_boot_en;
    uart_timeout_en_ff <= uart_timeout_en;
end
assign mux_sel_rst_state  = uart_boot_en_ff ? INIT_SEL : TEST_SEL ;
always @(posedge axi_clk) begin
    if (~axi_rst_n) begin
        mux_sel <= mux_sel_rst_state;
        writer_str_sel <= 0;
    end
    else begin
        case (mux_sel)
        INIT_SEL: begin
            if (init_done) begin
                mux_sel <= WRITER_SEL;
                writer_str_sel <= 0;
            end
        end
        WRITER_SEL: begin
            if (writer_finish) begin
                mux_sel <= READER_SEL;
            end
        end
        READER_SEL: begin
            if (reader_stop)
                mux_sel <= TEST_SEL;
        end
        TEST_SEL: begin
            mux_sel <=  pc_good_trap | pc_bad_trap | asm_test_timeout ? WRITER_SEL   : mux_sel;
            writer_str_sel <=   pc_good_trap        ?   1  :
                                pc_bad_trap         ?   2  :
                                asm_test_timeout    ?   3 : writer_str_sel;         
        end
        default: begin
            mux_sel <= mux_sel;
        end
        endcase
    end
end
assign writer_start = mux_sel == WRITER_SEL;
assign reader_start = mux_sel == READER_SEL;
assign test_start   = mux_sel == TEST_SEL;
assign  core_axi_awready    = s_axi_awready;
assign  core_axi_wready     = s_axi_wready;
assign  core_axi_bresp      = s_axi_bresp;
assign  core_axi_bvalid     = s_axi_bvalid;
assign  core_axi_arready    = s_axi_arready;
assign  core_axi_rdata      = s_axi_rdata;
assign  core_axi_rresp      = s_axi_rresp;
assign  core_axi_rvalid     = s_axi_rvalid;
assign  init_axi_awready    = s_axi_awready;
assign  init_axi_wready     = s_axi_wready;
assign  init_axi_bresp      = s_axi_bresp;
assign  init_axi_bvalid     = s_axi_bvalid;
assign  writer_axi_awready  = s_axi_awready;
assign  writer_axi_wready   = s_axi_wready;
assign  writer_axi_bresp    = s_axi_bresp;
assign  writer_axi_bvalid   = s_axi_bvalid;
assign  writer_axi_arready  = s_axi_arready;
assign  writer_axi_rdata    = s_axi_rdata;
assign  writer_axi_rresp    = s_axi_rresp;
assign  writer_axi_rvalid   = s_axi_rvalid;
assign  reader_axi_arready  = s_axi_arready;
assign  reader_axi_rdata    = s_axi_rdata;
assign  reader_axi_rresp    = s_axi_rresp;
assign  reader_axi_rvalid   = s_axi_rvalid;
always @(*) begin
    
    s_axi_awaddr    = 13'b0;
    s_axi_awvalid   = 1'b0;
    s_axi_wdata     = 32'b0;
    s_axi_wstrb     = 4'b0;
    s_axi_wvalid    = 1'b0;
    s_axi_bready    = 1'b0;
    s_axi_araddr    = 13'b0;
    s_axi_arvalid   = 1'b0;
    s_axi_rready    = 1'b0;
    case(mux_sel)
        INIT_SEL: begin
            s_axi_awaddr    = init_axi_awaddr;
            s_axi_awvalid   = init_axi_awvalid;
            s_axi_wdata     = init_axi_wdata;
            s_axi_wstrb     = init_axi_wstrb;
            s_axi_wvalid    = init_axi_wvalid;
            s_axi_bready    = init_axi_bready;
        end
        WRITER_SEL: begin
            s_axi_awaddr    = writer_axi_awaddr;
            s_axi_awvalid   = writer_axi_awvalid;
            s_axi_wdata     = writer_axi_wdata;
            s_axi_wstrb     = writer_axi_wstrb;
            s_axi_wvalid    = writer_axi_wvalid;
            s_axi_bready    = writer_axi_bready;
            s_axi_araddr    = writer_axi_araddr;
            s_axi_arvalid   = writer_axi_arvalid;
            s_axi_rready    = writer_axi_rready;
        end
        READER_SEL: begin
            s_axi_araddr    = reader_axi_araddr;
            s_axi_arvalid   = reader_axi_arvalid;
            s_axi_rready    = reader_axi_rready;
        end
        TEST_SEL: begin
            s_axi_awaddr    = core_axi_awaddr;
            s_axi_awvalid   = core_axi_awvalid;
            s_axi_wdata     = core_axi_wdata;
            s_axi_wstrb     = core_axi_wstrb;
            s_axi_wvalid    = core_axi_wvalid;
            s_axi_bready    = core_axi_bready;
            s_axi_araddr    = core_axi_araddr;
            s_axi_arvalid   = core_axi_arvalid;
            s_axi_rready    = core_axi_rready;
        end
        default: ;
    endcase
end
always @(posedge axi_clk) begin
    if (~axi_rst_n)
        asm_test_cycle_cnt <= 64'b0;
    else
        asm_test_cycle_cnt <=   reader_start & reader_stop      ?   64'b0                   :
                                test_start & ~asm_test_timeout  ?   asm_test_cycle_cnt + 1  :
                                                                    asm_test_cycle_cnt      ;
end
   
    assign asm_test_timeout = 1'b0;
    assign pc_good_trap     = 1'b0;
    assign pc_bad_trap      = 1'b0;
  
endmodule
    
    
    
     
    
    
    
    
    
    
    
    
    
    
    
    
         
         
   
    
   
    
       
        
        
    
  
   
     
    
   
   
    
    
module uart_reader (
    input                                 axi_clk,      
    input                                 axi_rst_n,    
    input                                 start,        
    output  reg                           stop,       
    output  [31:0]                        m_axi_araddr,
    output                                m_axi_arvalid,
    input                                 m_axi_arready,
    input   [31:0]                        m_axi_rdata,
    input   [1:0]                         m_axi_rresp,
    input                                 m_axi_rvalid,
    output                                m_axi_rready,
    input   [14-1:0]       chip_id,
    input   [8-1:0]            x_id,
    input   [8-1:0]            y_id,
    output                                noc_valid,
    output  [64-1:0]         noc_data,
    input                                 noc_ready
);
localparam  RD_STOP             = 0;
localparam  TEST_RXRD           = 1;
localparam  WAIT_RXRD_RESP      = 2;
localparam  READ_DATA           = 3;
localparam  WAIT_DATA           = 4;
localparam  IDLE                = 0;
localparam  ADDR                = 1;
localparam  BLK_NUM             = 2;
localparam  BLK                 = 3;
localparam  NOC_INTF_IDLE       = 0;
localparam  NOC_INTF_HDR        = 1;
localparam  NOC_INTF_DATA       = 2;
localparam  NOC_HDR_LEN         = 3;
reg             start_r;
reg             active;
reg             finish;
reg     [2:0]   rd_state;
reg     [1:0]                     gr_state;
reg     [1:0]                     gr_state_r;
reg     [40-1   : 0]  gr_addr;
reg     [8-1   : 0]  gr_blk_num;
reg     [8*64-1    : 0]  gr_blk;
reg     [clogb2(255+1)-1: 0]  gr_blk_cnt;
reg     [clogb2(255+1)-1: 0]  pcblk_in_strgblk_cnt;
reg     [clogb2(255+1)-1: 0]  pcblk_in_strgblk_cnt_r;
reg     [clogb2(255+1)-1: 0]  strgblk_in_gr_cnt;
reg     [clogb2(255+1)-1: 0]  strgblk_in_gr_cnt_prev;
reg     [7:0]   flit_cnt; 
reg     [40-1   : 0]  start_window;
reg     [8*64-1  : 0]    gr_blk_r;
reg     [1:0]                     noc_intf_state;
reg     [2:0]                     noc_cnt;
wire            launch;
wire            rresp_rx_rdy;
wire            rresp_rx_not_rdy;
wire            r_sent;
wire            state_rd_stop;
wire            state_test_rxrd;
wire            state_read_data;
wire            state_wait_data;
wire            gr_state_idle;
wire            gr_state_addr;
wire            gr_state_blk_num;
wire            gr_state_blk;
wire            gr_end;
wire    [7:0]   rdata;
wire            end_detected;
wire            storage_msg_ready;
wire    [40-1:0]    blk_addr;
wire            noc_last_hdr_val;
wire            noc_last_data_val;
wire    [64-1:0]       noc_hdr1_data;
wire    [64-1:0]       noc_hdr2_data;
wire    [64-1:0]       noc_hdr3_data;
wire    [8*64-1:0]       data_to_storage;
wire    [64-1:0]       noc_data_to_send [8-1:0];
wire [14-1:0]       source_chip_id;
wire [14-1:0]       dest_chip_id;
wire [8-1:0]            dest_x_id;
wire [8-1:0]            dest_y_id;
genvar i;
assign source_chip_id = chip_id;
assign dest_chip_id = chip_id;
assign dest_x_id = x_id;
assign dest_y_id = y_id;
assign m_axi_rready = 1'b1;
assign launch = start & ~start_r;
assign rresp_rx_rdy     = m_axi_rvalid & m_axi_rdata[0];
assign rresp_rx_not_rdy = m_axi_rvalid & ~m_axi_rdata[0];
assign r_sent        = m_axi_arvalid & m_axi_arready;
assign state_rd_stop       = rd_state == IDLE;
assign state_test_rxrd  = rd_state == TEST_RXRD;
assign state_read_data  = rd_state == READ_DATA;
assign state_wait_data  = rd_state == WAIT_DATA;
assign rdata_val        = m_axi_rvalid & state_wait_data;
assign rdata            = m_axi_rdata[7:0];
assign gr_state_idle    = gr_state == IDLE;
assign gr_state_addr    = gr_state == ADDR;
assign gr_state_blk_num = gr_state == BLK_NUM;
assign gr_state_blk     = gr_state == BLK;
assign gr_end           = (gr_state_r == BLK) & (gr_state == ADDR);
assign end_detected     = gr_state_blk_num & 
                          (gr_addr == 40'hffffffffff) &
                          rdata_val & (rdata == 8'b0);
always @(posedge axi_clk) begin
  start_r <= start;
end
always @(posedge axi_clk) begin
    active <= launch  ? 1'b1  :
              stop    ? 1'b0  : active;   
end
always @(posedge axi_clk) begin
  if (~axi_rst_n) begin
    finish <= 1'b0;    
  end
  else begin
    finish <= launch                ? 1'b0  :
              active & end_detected ? 1'b1  : finish;
  end
end
always @(posedge axi_clk) begin
  if (~axi_rst_n) begin
    stop <= 1'b0;    
  end
  else begin
    stop <= launch | ~active         ? 1'b0  :
            active & state_rd_stop   ? 1'b1  : stop;
  end
end
always @(posedge axi_clk) begin
  if (~axi_rst_n) begin
    rd_state <= RD_STOP;        
  end
  else begin
  
     
    case(rd_state)
      RD_STOP: begin
        if (launch)
          rd_state <= WAIT_DATA;
      end
      WAIT_DATA: begin
        if (m_axi_rvalid)
          rd_state <= finish ? RD_STOP : WAIT_DATA;
      end
      default: begin
      end
    endcase
    
  end
end
assign m_axi_arvalid  = (active & state_test_rxrd) |
                        (active & state_read_data) ;
assign m_axi_araddr   = (active & state_test_rxrd) ? 32'h1014 : 32'h1000;
always @(posedge axi_clk) begin
    start_window <= rdata_val ? {start_window[40-9:0], rdata} : start_window;
end
always @(posedge axi_clk) begin
  if (~axi_rst_n) begin
    gr_state <= IDLE;    
  end
  else begin
    case (gr_state)
      IDLE: begin
        if (start_window == 40'haaaaaaaaaa)
          gr_state <= ADDR;
      end
      ADDR: begin
        if (flit_cnt == 40/8)
          gr_state <= BLK_NUM;
        else if (finish)
          gr_state <= IDLE;
      end
      BLK_NUM: begin
        if (flit_cnt == 1)
          gr_state <= BLK;
      end
      BLK: begin
        if (gr_blk_cnt == gr_blk_num)
          gr_state <= ADDR;
      end
      default: begin
         gr_state  <= gr_state;
      end
    endcase
  end
end
always @(posedge axi_clk) begin
  if (~axi_rst_n) begin
    flit_cnt <= 8'b0;    
  end
  else begin
    flit_cnt <= (gr_state_addr & (flit_cnt == 40/8))       |
                (gr_state_blk_num & (flit_cnt == 1)) |
                (gr_state_blk & (flit_cnt == 8*64/8))         ? 8'b0         :
                active & rdata_val & ~gr_state_idle                     ? flit_cnt + 1 : flit_cnt;
  end
end
always @(posedge axi_clk) begin
    gr_addr <= rdata_val & gr_state_addr  ? {gr_addr[40-9:0], rdata} :
                                             gr_addr;
end
always @(posedge axi_clk) begin
  if (~axi_rst_n)
    gr_blk_num <= {8{1'b0}};
  else
    gr_blk_num <= rdata_val & gr_state_blk_num ? rdata : gr_blk_num;
end
always @(posedge axi_clk) begin
    gr_blk <= rdata_val & gr_state_blk  ? {gr_blk[8*64-9:0], rdata} :
                                          gr_blk;
end
always @(posedge axi_clk) begin
  if (~axi_rst_n)
    gr_blk_cnt <= {clogb2(255+1){1'b0}};
  else
    gr_blk_cnt <= gr_state_blk & (flit_cnt == 8*64/8) ? gr_blk_cnt + 1            :
                  gr_blk_cnt == gr_blk_num                      ? {clogb2(255+1){1'b0}} :
                                                                  gr_blk_cnt;
end
always @(posedge axi_clk) begin
  if (~axi_rst_n) begin
    pcblk_in_strgblk_cnt <= {clogb2(255+1){1'b0}};    
  end
  else begin
    pcblk_in_strgblk_cnt <= gr_state_blk & (flit_cnt == 8*64/8) ? pcblk_in_strgblk_cnt + 1        :
                      (pcblk_in_strgblk_cnt == 1) | gr_end  ? {clogb2(255+1){1'b0}} :
                                                                      pcblk_in_strgblk_cnt;
  end
end
always @(posedge axi_clk) begin
    pcblk_in_strgblk_cnt_r <= pcblk_in_strgblk_cnt;
end
always @(posedge axi_clk) begin
  if (~axi_rst_n) begin
    strgblk_in_gr_cnt <= {clogb2(255+1){1'b0}};    
  end
  else begin
    strgblk_in_gr_cnt <= gr_state_blk & (pcblk_in_strgblk_cnt == 1)   ? strgblk_in_gr_cnt + 1         :
                     gr_end                                               ? {clogb2(255+1){1'b0}} :
                                                                            strgblk_in_gr_cnt;
  end
end
always @(posedge axi_clk) begin
  if (~axi_rst_n)
    strgblk_in_gr_cnt_prev <= {clogb2(255+1){1'b0}};
  else
    strgblk_in_gr_cnt_prev <= noc_last_hdr_val ? strgblk_in_gr_cnt : strgblk_in_gr_cnt_prev;
end
always @(posedge axi_clk) begin
    gr_state_r <= gr_state;
end
assign storage_msg_ready = active                                           & 
                          ((pcblk_in_strgblk_cnt_r == 1) | gr_end) &
                          (gr_addr != 40'hffffffffff);
always @(posedge axi_clk) begin
  gr_blk_r <= gr_state_blk & (flit_cnt == 8*64/8)   ? gr_blk : gr_blk_r;
end
assign data_to_storage = gr_blk_r;
assign blk_addr = gr_addr + (strgblk_in_gr_cnt_prev << 6);
always @(posedge axi_clk) begin
  if (~axi_rst_n) begin
    noc_intf_state <= NOC_INTF_IDLE;
  end
  else begin
    case (noc_intf_state)
      NOC_INTF_IDLE: begin
        if (storage_msg_ready)
          noc_intf_state <= NOC_INTF_HDR;
      end
      NOC_INTF_HDR: begin
        if (noc_last_hdr_val)
          noc_intf_state <= NOC_INTF_DATA;
      end
      NOC_INTF_DATA: begin
        if (noc_last_data_val)
          noc_intf_state <= NOC_INTF_IDLE;
      end
      default: begin
      end
    endcase
  end
end
always @(posedge axi_clk) begin
  if (~axi_rst_n) begin
    noc_cnt <= 3'b0;
  end
  else begin
    noc_cnt <=  noc_last_hdr_val | noc_last_data_val  ? 3'b0        :
                noc_valid & noc_ready                 ? noc_cnt + 1 : noc_cnt;  
  end
end
assign noc_valid = noc_intf_state != NOC_INTF_IDLE;
assign noc_hdr1_data      = {chip_id, 8'h0, 8'h0, 4'h0, 8'ha, 8'h14, 8'h0, 6'h0};
assign noc_hdr2_data      = {8'h0, blk_addr, 16'h0};
assign noc_hdr3_data      = {chip_id, x_id, y_id, 4'b0, 30'h0};
generate
  for (i = 0; i < 8; i = i + 1) begin: NOC_DATA
    assign noc_data_to_send[i] = data_to_storage[64*(i+1)-1:64*i];
  end
endgenerate
assign noc_data           = (noc_intf_state == NOC_INTF_HDR) & (noc_cnt == 0) ? noc_hdr1_data :
                            (noc_intf_state == NOC_INTF_HDR) & (noc_cnt == 1) ? noc_hdr2_data :
                            (noc_intf_state == NOC_INTF_HDR) & (noc_cnt == 2) ? noc_hdr3_data :
                                                                                noc_data_to_send[noc_cnt];
assign noc_last_hdr_val   = (noc_intf_state == NOC_INTF_HDR)  &
                            (noc_cnt == NOC_HDR_LEN-1)        &
                            noc_ready;
assign noc_last_data_val  = (noc_intf_state == NOC_INTF_DATA) &
                            (noc_cnt == 8-1)       &
                            noc_ready; 
function integer clogb2;
  input [31:0] value;
  begin
    value = value - 1;
    for (clogb2 = 0; value > 0; clogb2 = clogb2 + 1) begin
      value = value >> 1;
    end
  end
endfunction
endmodule
    
    
    
     
    
    
    
    
    
    
    
    
    
    
    
    
   
    
   
    
       
        
        
    
  
   
     
    
   
   
    
    
module uart_top (
    input                                   axi_clk,
    input                                   rst_n,
   
    output                                  uart_tx,
    input                                   uart_rx,
    output                  uart_interrupt,
    input                                   uart_lb_sw,
    input                                   uart_boot_en,
    input                                   uart_timeout_en,
    output                                  test_start,
    input                                   test_good_end,
    input                                   test_bad_end,
    output                                  uart_rst_out_n,
    input                                   init_calib_complete,
    input [14-1:0]          chip_id,
    input [8-1:0]                x_id,
    input [8-1:0]                y_id,
    
    input                                   xbar_uart_noc2_valid,
    input [64-1:0]             xbar_uart_noc2_data,     
    output                                  uart_xbar_noc2_ready,
    output                                  uart_xbar_noc3_valid,
    output [64-1:0]            uart_xbar_noc3_data,  
    input                                   xbar_uart_noc3_ready,
    
    
    output                                  uart_xbar_noc2_valid,
    output [64-1:0]            uart_xbar_noc2_data,  
    input                                   xbar_uart_noc2_ready,
    input                                   xbar_uart_noc3_valid,
    input [64-1:0]             xbar_uart_noc3_data,     
    output                                  uart_xbar_noc3_ready
);
wire  uart16550_tx;
wire  uart16550_rx;
wire  [12:0]      s_axi_awaddr;
wire              s_axi_awvalid;
wire              s_axi_awready;
wire  [31:0]      s_axi_wdata;
wire  [3:0 ]      s_axi_wstrb;
wire              s_axi_wvalid;
wire              s_axi_wready;
wire  [1:0]       s_axi_bresp;
wire              s_axi_bvalid;
wire              s_axi_bready;
wire  [12:0]      s_axi_araddr;
wire              s_axi_arvalid;
wire              s_axi_arready;
wire  [31:0]      s_axi_rdata;
wire  [1:0]       s_axi_rresp;
wire              s_axi_rvalid;
wire              s_axi_rready;
wire              init_done;
wire              atg_init_done;
wire              writer_start;
wire              writer_finish;
wire  [2:0]       writer_str_sel;
wire              reader_start;
wire              reader_stop;
wire [12:0]                        core_axi_awaddr;
wire                               core_axi_awvalid;
wire                               core_axi_awready;
wire [31:0]                        core_axi_wdata;
wire [3:0]                         core_axi_wstrb;
wire                               core_axi_wvalid;
wire                               core_axi_wready;
wire [1:0]                         core_axi_bresp;
wire                               core_axi_bvalid;
wire                               core_axi_bready;
wire [12:0]                        core_axi_araddr;
wire                               core_axi_arvalid;
wire                               core_axi_arready;
wire [31:0]                        core_axi_rdata;
wire [1:0]                         core_axi_rresp;
wire                               core_axi_rvalid;
wire                               core_axi_rready;
(* DONT_TOUCH = "yes" *)wire    [64-1:0]  core_axi_awaddr_unmasked;
(* DONT_TOUCH = "yes" *)wire    [64-1:0]  core_axi_araddr_unmasked;
assign core_axi_awaddr = (core_axi_awaddr_unmasked[12:0] << 2)  | 13'h1000;
assign core_axi_araddr = (core_axi_araddr_unmasked[12:0] << 2)  | 13'h1000;
assign uart_xbar_noc3_ready = 1'b1;
noc_axilite_bridge #(
    .SLAVE_RESP_BYTEWIDTH   (1)
) noc_axilite_bridge (
    .clk                    (axi_clk                ),
    .rst                    (~rst_n             ),  
           
    .splitter_bridge_val    (xbar_uart_noc2_valid   ),
    .splitter_bridge_data   (xbar_uart_noc2_data  ),
    .bridge_splitter_rdy    (uart_xbar_noc2_ready   ),
    .bridge_splitter_val    (uart_xbar_noc3_valid   ),
    .bridge_splitter_data   (uart_xbar_noc3_data  ),
    .splitter_bridge_rdy    (xbar_uart_noc3_ready   ),
       
    
    
    .m_axi_awaddr        (core_axi_awaddr_unmasked),
    .m_axi_awvalid       (core_axi_awvalid),
    .m_axi_awready       (core_axi_awready),
    
    .m_axi_wdata         (core_axi_wdata),
    .m_axi_wstrb         (core_axi_wstrb),
    .m_axi_wvalid        (core_axi_wvalid),
    .m_axi_wready        (core_axi_wready),
    
    .m_axi_araddr        (core_axi_araddr_unmasked),
    .m_axi_arvalid       (core_axi_arvalid),
    .m_axi_arready       (core_axi_arready),
    
    .m_axi_rdata         (core_axi_rdata),
    .m_axi_rresp         (core_axi_rresp),
    .m_axi_rvalid        (core_axi_rvalid),
    .m_axi_rready        (core_axi_rready),
    
    .m_axi_bresp         (core_axi_bresp),
    .m_axi_bvalid        (core_axi_bvalid),
    .m_axi_bready        (core_axi_bready)
    
);
assign uart_tx        = uart_lb_sw ? uart_rx  : uart16550_tx;
assign uart16550_rx   = uart_rx; 
   
  
    
       
      assign init_done = 1'b1;
      
    
  
  
     
    assign writer_finish      = 1'b1;
    
   
  assign reader_stop = 1'b1;
  
 
  assign uart_rst_out_n = 1'b1;
uart_mux   uart_mux (
  .axi_clk              (axi_clk            ),
  .axi_rst_n            (rst_n              ),
  .uart_boot_en         (uart_boot_en       ),
  .uart_timeout_en      (uart_timeout_en    ),
  .init_done            (init_done          ),
  .writer_start         (writer_start       ),
  .writer_finish        (writer_finish      ),
  .writer_str_sel       (writer_str_sel     ),
  .reader_start         (reader_start       ),
  .reader_stop          (reader_stop        ),
  .test_start           (test_start         ),
  .test_good_end        (test_good_end      ),
  .test_bad_end         (test_bad_end       ),
 
  .core_axi_awaddr      (core_axi_awaddr    ),
  .core_axi_awvalid     (core_axi_awvalid   ),
  .core_axi_awready     (core_axi_awready   ),
  .core_axi_wdata       (core_axi_wdata     ),
  .core_axi_wstrb       (core_axi_wstrb     ),
  .core_axi_wvalid      (core_axi_wvalid    ),
  .core_axi_wready      (core_axi_wready    ),
  .core_axi_bresp       (core_axi_bresp     ),
  .core_axi_bvalid      (core_axi_bvalid    ),
  .core_axi_bready      (core_axi_bready    ),
  .core_axi_araddr      (core_axi_araddr    ),
  .core_axi_arvalid     (core_axi_arvalid   ),
  .core_axi_arready     (core_axi_arready   ),
  .core_axi_rdata       (core_axi_rdata     ),
  .core_axi_rresp       (core_axi_rresp     ),
  .core_axi_rvalid      (core_axi_rvalid    ),
  .core_axi_rready      (core_axi_rready    ),
  .s_axi_awaddr         (s_axi_awaddr       ),
  .s_axi_awvalid        (s_axi_awvalid      ),
  .s_axi_awready        (s_axi_awready      ),
  .s_axi_wdata          (s_axi_wdata        ),
  .s_axi_wstrb          (s_axi_wstrb        ),
  .s_axi_wvalid         (s_axi_wvalid       ),
  .s_axi_wready         (s_axi_wready       ),
  .s_axi_bresp          (s_axi_bresp        ),
  .s_axi_bvalid         (s_axi_bvalid       ),
  .s_axi_bready         (s_axi_bready       ),
  .s_axi_araddr         (s_axi_araddr       ),
  .s_axi_arvalid        (s_axi_arvalid      ),
  .s_axi_arready        (s_axi_arready      ),
  .s_axi_rdata          (s_axi_rdata        ),
  .s_axi_rresp          (s_axi_rresp        ),
  .s_axi_rvalid         (s_axi_rvalid       ),
  .s_axi_rready         (s_axi_rready       )
);
   
  
    
    
      
    
  
endmodule
         
         
   
    
   
    
       
        
        
    
  
   
     
    
   
   
    
    
module  uart_writer (
  input                 axi_clk,
  input                 axi_rst_n,
  input                 start,
  output  reg           finish,
  input   [2:0]         str_sel,
  output  [12:0]        m_axi_awaddr,
  output                m_axi_awvalid,
  input                 m_axi_awready,
  output  [31:0]        m_axi_wdata,
  output  [3:0]         m_axi_wstrb,
  output                m_axi_wvalid,
  input                 m_axi_wready,
  input   [1:0]         m_axi_bresp,
  input                 m_axi_bvalid,
  output                m_axi_bready,
  output  [31:0]        m_axi_araddr,
  output                m_axi_arvalid,
  input                 m_axi_arready,
  input   [31:0]        m_axi_rdata,
  input   [1:0]         m_axi_rresp,
  input                 m_axi_rvalid,
  output                m_axi_rready
);
localparam LINE_CNTR_WIDTH = 9;
localparam LINE_NUMBER = 16;
localparam CHAR_WIDTH = 8;
localparam WAIT_TX    = 0;
localparam WAIT_RRESP = 1;
localparam SEND_DATA  = 2;
localparam LINE_0_LEN = 4;
localparam LINE_1_LEN = 6;
localparam LINE_2_LEN = 6;
localparam LINE_3_LEN = 7;
wire  [LINE_CNTR_WIDTH-1:0] str_len [LINE_NUMBER-1:0];
assign str_len[0] = LINE_0_LEN;
assign str_len[1] = LINE_1_LEN;
assign str_len[2] = LINE_1_LEN;
assign str_len[3] = LINE_3_LEN;
reg   [CHAR_WIDTH-1:0]  line_0 [LINE_0_LEN-1:0];  
reg   [CHAR_WIDTH-1:0]  line_1 [LINE_1_LEN-1:0];  
reg   [CHAR_WIDTH-1:0]  line_2 [LINE_2_LEN-1:0];  
reg   [CHAR_WIDTH-1:0]  line_3 [LINE_3_LEN-1:0];  
always @(posedge axi_clk) begin
  line_0[0] <= 8'h44;
  line_0[1] <= 8'h4f;
  line_0[2] <= 8'h4e;
  line_0[3] <= 8'h45;
end
always @(posedge axi_clk) begin
  line_1[0] <= 8'h50;
  line_1[1] <= 8'h41;
  line_1[2] <= 8'h53;
  line_1[3] <= 8'h53;
  line_1[4] <= 8'h45;
  line_1[5] <= 8'h44;
end
always @(posedge axi_clk) begin
  line_2[0] <= 8'h46;
  line_2[1] <= 8'h41;
  line_2[2] <= 8'h49;
  line_2[3] <= 8'h4c;
  line_2[4] <= 8'h45;
  line_2[5] <= 8'h44;
end
always @(posedge axi_clk) begin
  line_3[0] <= 8'h54;
  line_3[1] <= 8'h49;
  line_3[2] <= 8'h4d;
  line_3[3] <= 8'h45;
  line_3[4] <= 8'h4f;
  line_3[5] <= 8'h55;
  line_3[6] <= 8'h54;
end
assign m_axi_bready   = 1'b1;
assign m_axi_rready   = 1'b1;
reg [1:0]   state;
reg         start_r;
reg         writer_active;
reg [LINE_CNTR_WIDTH-1:0]   char_cnt;
wire          ar_sent;
wire          tx_sent;
wire          launch_writer;
wire  [7:0]   curr_char;
wire  [LINE_CNTR_WIDTH-1:0]   curr_line_len;
wire [CHAR_WIDTH-1:0]   char_0;
wire [CHAR_WIDTH-1:0]   char_1;
wire [CHAR_WIDTH-1:0]   char_2;
wire [CHAR_WIDTH-1:0]   char_3;
assign ar_sent         = m_axi_arvalid & m_axi_arready;
assign tx_sent        = m_axi_wvalid  & m_axi_wready;
assign state_wait_tx  = state == WAIT_TX;
assign state_send_d   = state == SEND_DATA;
always @(posedge axi_clk) begin
  start_r <= start;
end
assign launch_writer = start & ~start_r;
always @(posedge axi_clk) begin
  if (~axi_rst_n)
    writer_active <= 1'b0;
  else
    writer_active <= launch_writer    ? 1'b1  :
                     finish           ? 1'b0  : writer_active;
end
always @(posedge axi_clk) begin
  if (~axi_rst_n)
    finish <= 1'b0;
  else
    finish <= writer_active & (char_cnt == curr_line_len);
end
assign rresp_tx_emp     = m_axi_rvalid & m_axi_rdata[6];
assign rresp_tx_no_emp  = m_axi_rvalid & ~m_axi_rdata[6];
assign m_axi_arvalid    = writer_active & state_wait_tx;
assign m_axi_araddr     = 32'h1014;
assign m_axi_wvalid     = writer_active & state_send_d;
assign m_axi_wdata      = curr_char;
assign m_axi_awvalid    = writer_active & state_send_d;
assign m_axi_awaddr     = 32'h1000;
assign m_axi_wstrb      = 4'hf;
always @(posedge axi_clk) begin
  if (~axi_rst_n) begin
    state <= WAIT_TX;
  end
  else begin
  
  
    state <= SEND_DATA;
  
  end
end
always @(posedge axi_clk) begin
  if (~axi_rst_n)
    char_cnt <= {LINE_CNTR_WIDTH{1'b0}};
  else begin
    char_cnt <= launch_writer             ? {LINE_CNTR_WIDTH{1'b0}} :
                writer_active & tx_sent   ?  char_cnt + 1           : char_cnt;
  end
end
assign char_0 = line_0[char_cnt];
assign char_1 = line_1[char_cnt];
assign char_2 = line_2[char_cnt];
assign char_3 = line_3[char_cnt];
assign curr_char =  ({8{str_sel == 0}} & char_0) |
                    ({8{str_sel == 1}}   & char_1) |
                    ({8{str_sel == 2}}   & char_2) |
                    ({8{str_sel == 3}}  & char_3) ;
assign curr_line_len = str_len[str_sel];
endmodule
module io_xbar_space_avail_top (valid,
		    yummy,
		    spc_avail,
		    clk,
		    reset);
parameter BUFFER_SIZE = 4;
parameter BUFFER_BITS = 3;
   
 
input valid;			
input yummy;			
output spc_avail;		
input clk;
input reset;
reg yummy_f;
reg valid_f;
reg [BUFFER_BITS-1:0] count_f;
reg is_one_f;
reg is_two_or_more_f;
wire [BUFFER_BITS-1:0] count_plus_1;
wire [BUFFER_BITS-1:0] count_minus_1;
wire up;
wire down;
reg [BUFFER_BITS-1:0] count_temp;
assign count_plus_1 = count_f + 1'b1;
assign count_minus_1 = count_f - 1'b1;
assign spc_avail = (is_two_or_more_f | yummy_f | (is_one_f & ~valid_f));
assign up = yummy_f & ~valid_f;
assign down = ~yummy_f & valid_f;
always @ (count_f or count_plus_1 or count_minus_1 or up or down)
begin
	case (count_f)
	0:
		begin
			if(up)
			begin
				count_temp <= count_plus_1;
			end
			else
			begin
				count_temp <= count_f;
			end
		end
	BUFFER_SIZE:
		begin
			if(down)
			begin
				count_temp <= count_minus_1;
			end
			else
			begin
				count_temp <= count_f;
			end
		end
	default:
		begin
			case ({up, down})
				2'b10:	count_temp <= count_plus_1;
				2'b01:	count_temp <= count_minus_1;
				default:	count_temp <= count_f;
			endcase
		end
	endcase
end
wire top_bits_zero_temp = ~| count_temp[BUFFER_BITS-1:1];
always @ (posedge clk)
begin
	if(reset)
	begin
	   count_f <= BUFFER_SIZE;
	   yummy_f <= 1'b0;
	   valid_f <= 1'b0;
	   is_one_f <= (BUFFER_SIZE == 1);
	   is_two_or_more_f <= (BUFFER_SIZE >= 2);
	end
	else
	begin
	   count_f <= count_temp;
	   yummy_f <= yummy;
	   valid_f <= valid;
	   is_one_f         <= top_bits_zero_temp & count_temp[0];
   	   is_two_or_more_f <= ~top_bits_zero_temp;
	end
end
endmodule
      
  
          
      
    
         
module jtag(
    input clk,
    input rst_n,
    
    input wire jtag_clk,
    input wire jtag_rst_l,
    input wire jtag_modesel,
    input wire jtag_datain,
    output wire jtag_dataout,
    output wire jtag_dataout_en,
    
    output wire jtag_tiles_ucb_val,
    output wire [4-1:0] jtag_tiles_ucb_data,
    
    input wire tiles_jtag_ucb_val,
    input wire [4-1:0] tiles_jtag_ucb_data,
    output wire ctap_oram_req_val,
    output wire [4-1:0] ctap_oram_req_misc,
    input wire [64-1:0] oram_ctap_res_data,
    
    
    
    output wire [127:0] ctap_clk_en,
    output wire ctap_oram_clk_en
    );
wire sys_clk = clk;
wire jtag_ctap_reg_wr_en;
wire [4-1:0] jtag_ctap_reg_sel;
wire [128-1:0] jtag_ctap_data;
wire jtag_ctap_reg_wr_en_sync;
wire [4-1:0] jtag_ctap_reg_sel_sync;
wire [128-1:0] jtag_ctap_data_sync;
wire [128-1:0] ctap_jtag_data;
wire ctap_jtag_interrupt_bit;
wire [128-1:0] ctap_jtag_data_sync;
wire ctap_jtag_interrupt_bit_sync;
wire ctap_ucb_tx_val;
wire [128-1:0] ctap_ucb_tx_data;
wire [(128/4)-1:0] ctap_ucb_tx_data_vec;
wire ctap_ucb_rx_val;
wire [128-1:0] ctap_ucb_rx_data;
jtag_interface jtag_interface(
    .jtag_clk(jtag_clk),
    .jtag_rst_l(jtag_rst_l),
    .jtag_modesel(jtag_modesel),
    .jtag_datain(jtag_datain),
    .jtag_dataout(jtag_dataout),
    .jtag_dataout_en(jtag_dataout_en),
    .ctap_jtag_data(ctap_jtag_data_sync),
    .ctap_jtag_interrupt_bit(ctap_jtag_interrupt_bit_sync),
    .jtag_ctap_data(jtag_ctap_data),
    .jtag_ctap_reg_wr_en(jtag_ctap_reg_wr_en),
    .jtag_ctap_reg_sel(jtag_ctap_reg_sel)
    );
jtag_ctap ctap(
    .clk(clk),
    .rst_n(rst_n),
    
    .ctap_jtag_data(ctap_jtag_data),
    .ctap_jtag_interrupt_bit(ctap_jtag_interrupt_bit),
    .jtag_ctap_data(jtag_ctap_data_sync),
    .jtag_ctap_reg_wr_en(jtag_ctap_reg_wr_en_sync),
    .jtag_ctap_reg_sel(jtag_ctap_reg_sel_sync),
    .ctap_ucb_tx_val(ctap_ucb_tx_val),
    .ctap_ucb_tx_data(ctap_ucb_tx_data),
    .ctap_ucb_tx_data_vec(ctap_ucb_tx_data_vec),
    .ctap_ucb_rx_val(ctap_ucb_rx_val),
    .ctap_ucb_rx_data(ctap_ucb_rx_data),
    .ctap_oram_req_val(ctap_oram_req_val),
    .ctap_oram_req_misc(ctap_oram_req_misc),
    .oram_ctap_res_data(oram_ctap_res_data),
    
    
    
    .ctap_clk_en(ctap_clk_en),
    .ctap_oram_clk_en(ctap_oram_clk_en)
    );
synchronizer #(1) u_jtag_ctap_reg_wr_en_sync 
   ( .syncdata (jtag_ctap_reg_wr_en_sync),
     .presyncdata (jtag_ctap_reg_wr_en),
     .clk (sys_clk)
     );
assign jtag_ctap_reg_sel_sync = jtag_ctap_reg_sel;
assign jtag_ctap_data_sync = jtag_ctap_data;
assign ctap_jtag_data_sync = ctap_jtag_data;
synchronizer #(1) u_ctap_jtag_interrupt_bit_sync 
   ( .syncdata (ctap_jtag_interrupt_bit_sync),
     .presyncdata (ctap_jtag_interrupt_bit),
     .clk (jtag_clk)
     );
jtag_ucb_receiver ucb_rx(
    .clk(clk),
    .rst_n(rst_n),
    .ctap_ucb_rx_val(ctap_ucb_rx_val),
    .ctap_ucb_rx_data(ctap_ucb_rx_data),
    .tiles_jtag_ucb_val(tiles_jtag_ucb_val),
    .tiles_jtag_ucb_data(tiles_jtag_ucb_data)
    );
jtag_ucb_transmitter ucb_tx(
    .clk(clk),
    .rst_n(rst_n),
    .ctap_ucb_tx_val(ctap_ucb_tx_val),
    .ctap_ucb_tx_data(ctap_ucb_tx_data),
    .ctap_ucb_tx_data_vec(ctap_ucb_tx_data_vec),
    .jtag_tiles_ucb_val(jtag_tiles_ucb_val),
    .jtag_tiles_ucb_data(jtag_tiles_ucb_data)
    );
endmodule
  
          
      
    
         
module jtag_interface(
    
    input wire jtag_clk,
    input wire jtag_rst_l,
    input wire jtag_modesel,
    input wire jtag_datain,
    output wire jtag_dataout,
    output wire jtag_dataout_en,
    
    input wire [128-1:0] ctap_jtag_data,
    input wire ctap_jtag_interrupt_bit,
    output reg [128-1:0] jtag_ctap_data,
    output reg jtag_ctap_reg_wr_en,
    output reg [4-1:0] jtag_ctap_reg_sel
    );
wire jtag_clk_l = ~jtag_clk;
wire [18-1:0]   tap_instructions;
wire [18-1:0]   next_tap_instructions;
wire          tap_capture_dr_state;       
wire          tap_shift_dr_state;         
                                          
wire          tap_pause_dr_state;         
wire          tap_update_dr_state;        
wire          tap_shift_exit2_dr_state;   
wire          tap_update_ir_state;        
wire          tap_bypass_sel;
wire          instr_bypass;
wire          instr_idcode;
wire          instr_highz;
wire          instr_clamp;
reg [31:0]    idcode;
reg [31:0]    next_idcode;
reg [128-1:0] scratch_reg;
reg [128-1:0] scratch_reg_next;
wire          tap_scratch_sel;
wire          tap_so;
wire          instr_ctap_instruction_reg_sel;
wire          instr_ctap_data0_reg_sel;
wire          instr_ctap_address_reg_sel;
wire          instr_ctap_interrupt_bit_sel;
wire          next_instr_ctap_instruction_reg_sel;
wire          next_instr_ctap_data0_reg_sel;
wire          next_instr_ctap_address_reg_sel;
parameter TAP_CMD_LO    = 0,
    TAP_CMD_HI    = 6 - 1;
jtag_interface_tap u_tap_controller (
    
    .tck (jtag_clk),
    .tck_l (jtag_clk_l),
    .trst_n (jtag_rst_l),
    .tms (jtag_modesel),
    .tdi (jtag_datain),
    .so (tap_so),
    .bypass_sel (tap_bypass_sel), 
    .dft_pin_pscan(1'b0),
    
    .capture_dr_state (tap_capture_dr_state),
    .shift_dr_state (tap_shift_dr_state),
    .pause_dr_state (tap_pause_dr_state),
    .update_dr_state (tap_update_dr_state),
    .shift_exit2_dr_state (tap_shift_exit2_dr_state), 
    .update_ir_state (tap_update_ir_state),
    .clock_dr  (), 
    .tdo (jtag_dataout),
    .tdo_en (jtag_dataout_en),
    .instructions (tap_instructions), 
    .next_instructions (next_tap_instructions) 
    );
wire [6-1:0] tap_inst = tap_instructions[TAP_CMD_HI:TAP_CMD_LO];
wire [6-1:0] next_tap_inst = next_tap_instructions[TAP_CMD_HI:TAP_CMD_LO];
assign instr_bypass           = tap_inst == {6{1'b1}}
                                | (tap_instructions[TAP_CMD_HI:TAP_CMD_HI-3] == 4'b0001   
                                & (|tap_instructions[TAP_CMD_HI-4:TAP_CMD_LO]))
                                | (tap_instructions[TAP_CMD_HI:TAP_CMD_HI-3] == 4'b0100   
                                & (|tap_instructions[TAP_CMD_HI-4:TAP_CMD_LO]))
                                | tap_inst == 6'h19
                                | tap_inst == 6'h27
                                | tap_inst == 6'h2F
                                | tap_instructions[TAP_CMD_HI:TAP_CMD_HI-1] == 2'd3;
assign instr_idcode           = tap_inst == 6'h01;
assign instr_highz            = tap_inst == 6'h03;
assign instr_clamp            = tap_inst == 6'h04;
assign instr_ctap_instruction_reg_sel = tap_inst == 6'h08;
assign instr_ctap_data0_reg_sel = tap_inst == 6'h09;
assign instr_ctap_address_reg_sel = tap_inst == 6'h0a;
assign instr_ctap_interrupt_bit_sel = tap_inst == 6'h0b;
assign next_instr_ctap_instruction_reg_sel = next_tap_inst == 6'h08;
assign next_instr_ctap_data0_reg_sel = next_tap_inst == 6'h09;
assign next_instr_ctap_address_reg_sel = next_tap_inst == 6'h0a;
assign tap_scratch_sel = instr_ctap_instruction_reg_sel | instr_ctap_data0_reg_sel 
                        | instr_ctap_address_reg_sel;
assign tap_bypass_sel   = instr_highz  | instr_clamp | instr_bypass;
assign tap_so =   
       (idcode[0]                 & instr_idcode) 
       | (scratch_reg[128-1]   & tap_scratch_sel)
       | (ctap_jtag_interrupt_bit   & instr_ctap_interrupt_bit_sel)
       
       
       
       
       
       
       
       
       
       
       
       ;
wire [3:0] jtag_id = 4'b0;
always @ *
begin
    if (instr_idcode & tap_capture_dr_state)
        next_idcode = { jtag_id[3:0], 16'h1AAA, 11'h03E, 1'b1 };
    else begin
        if (instr_idcode & tap_shift_dr_state)
            
            next_idcode = { jtag_datain, idcode[31:1] }; 
        else
            next_idcode = idcode[31:0];
    end
end
always @ (posedge jtag_clk)
begin
    if (!jtag_rst_l)
    begin
        scratch_reg <= 128'b0;
        idcode <= 0;
    end
    else
    begin
        scratch_reg <= scratch_reg_next;
        idcode <= next_idcode;
    end
end
reg           scratch_reg_shift;
reg           scratch_reg_load;
always @ * 
begin
    scratch_reg_shift = tap_scratch_sel & tap_shift_dr_state;
    scratch_reg_load = tap_scratch_sel & tap_capture_dr_state;
    if (scratch_reg_shift)
        scratch_reg_next = {scratch_reg[128-2:0], jtag_datain};
    else if (scratch_reg_load)
        scratch_reg_next[128-1:0] = ctap_jtag_data[128-1:0];
    else
        scratch_reg_next = scratch_reg;
    
    jtag_ctap_data = scratch_reg;
    
    jtag_ctap_reg_wr_en = tap_update_dr_state && tap_scratch_sel;
end
reg [4-1:0] ctap_reg_sel;
reg [4-1:0] ctap_reg_sel_next;
always @ (posedge jtag_clk)
begin
    if (!jtag_rst_l)
    begin
        ctap_reg_sel <= 0;
    end
    else
        ctap_reg_sel <= ctap_reg_sel_next;
end
reg next_ctap_data0_sel;
always @ *
begin
    
    next_ctap_data0_sel = tap_update_ir_state & next_instr_ctap_data0_reg_sel;
    if (next_ctap_data0_sel)
        ctap_reg_sel_next = 4'd1;
    else if (next_instr_ctap_instruction_reg_sel)
        ctap_reg_sel_next = 4'd2;
    else if (next_instr_ctap_address_reg_sel)
        ctap_reg_sel_next = 4'd3;
    else
        ctap_reg_sel_next = ctap_reg_sel;
    
    jtag_ctap_reg_sel = ctap_reg_sel;
end
endmodule
  
    
    
    
    
    
    
    
        
        
        
        
        
        
        
        
        
        
        
 
        
        
        
        
  
          
      
    
         
module jtag_interface_tap(
instructions, next_instructions, capture_dr_state, shift_dr_state, 
pause_dr_state, update_dr_state, shift_exit2_dr_state, 
update_ir_state, clock_dr, tdo, tdo_en, 
tck, tck_l, trst_n, tms, tdi, so, bypass_sel, dft_pin_pscan
);
input  tck;
input  tck_l;
input  trst_n;
input  tms;
input  tdi;
input  so;
input  bypass_sel;
input  dft_pin_pscan;
output [18-1:0] instructions;
output [18-1:0] next_instructions;
output                capture_dr_state;
output                shift_dr_state;
output                pause_dr_state;
output                update_dr_state;
output                shift_exit2_dr_state;
output                update_ir_state;
output                clock_dr;
output                tdo;
output                tdo_en; 
                  
wire [18-1:0]   instructions;
reg [18-1:0]    next_instructions;
wire                  capture_dr_state;
wire                  shift_dr_state;
wire                  pause_dr_state;
wire                  update_dr_state;
wire                  shift_exit2_dr_state;
wire                  update_ir_state;
wire                  clock_dr;
wire                  tdo;
wire                  tdo_en; 
parameter TAP_RESET     = 16'h0001,
      TAP_TEST      = 16'h0002,
      TAP_SEL_DR    = 16'h0004,
      TAP_CAP_DR    = 16'h0008,
      TAP_SHIFT_DR  = 16'h0010,
      TAP_EXIT1_DR  = 16'h0020,
      TAP_PAUSE_DR  = 16'h0040,
      TAP_EXIT2_DR  = 16'h0080,
      TAP_UPDATE_DR = 16'h0100,
      TAP_SEL_IR    = 16'h0200,
      TAP_CAP_IR    = 16'h0400,
      TAP_SHIFT_IR  = 16'h0800,
      TAP_EXIT1_IR  = 16'h1000,
      TAP_PAUSE_IR  = 16'h2000,
      TAP_EXIT2_IR  = 16'h4000,
      TAP_UPDATE_IR = 16'h8000,
      TAP_STATE_WIDTH = 16;
parameter TAP_RESET_BIT     =  0,
      TAP_CAP_DR_BIT    =  3,
      TAP_SHIFT_DR_BIT  =  4,
      TAP_PAUSE_DR_BIT  =  6,
      TAP_EXIT2_DR_BIT  =  7,
      TAP_UPDATE_DR_BIT =  8,
      TAP_CAP_IR_BIT    = 10,
      TAP_SHIFT_IR_BIT  = 11,
      TAP_UPDATE_IR_BIT = 15;
wire [15:0] tap_state;
reg [15:0]  next_tap_state;
wire        tap_state_reset_negedge;
wire        capture_shift_dr;
wire        next_tap_state_reset_negedge;
wire        next_capture_shift_dr;
reg         next_tdo;
wire        next_tdo_en;
wire [18-1:0] new_instructions;
reg [18-1:0] next_new_instructions;
wire                reset_muxed;
wire                instructions_rst_l;
wire                tdi_ff;
wire                tdi_ff_en;
wire                tdi_ff_rst_l;
always @ ( tap_state or tms) begin
   case (tap_state)
      TAP_RESET: begin
     if (tms)
        next_tap_state = TAP_RESET;
     else
        next_tap_state = TAP_TEST;
      end
      TAP_TEST: begin
     if (tms)
        next_tap_state = TAP_SEL_DR;
     else
        next_tap_state = TAP_TEST;
      end
      TAP_SEL_DR: begin
     if (tms)
        next_tap_state = TAP_SEL_IR;
     else
        next_tap_state = TAP_CAP_DR;
      end
      TAP_CAP_DR: begin
     if (tms)
        next_tap_state = TAP_EXIT1_DR;
     else
        next_tap_state = TAP_SHIFT_DR;
      end
      TAP_SHIFT_DR: begin
     if (tms)
        next_tap_state = TAP_EXIT1_DR;
     else
        next_tap_state = TAP_SHIFT_DR;
      end
      TAP_EXIT1_DR: begin
     if (tms)
        next_tap_state = TAP_UPDATE_DR;
     else
        next_tap_state = TAP_PAUSE_DR;
      end
      TAP_PAUSE_DR: begin
     if (tms)
        next_tap_state = TAP_EXIT2_DR;
     else
        next_tap_state = TAP_PAUSE_DR;
      end
      TAP_EXIT2_DR: begin
     if (tms)
        next_tap_state = TAP_UPDATE_DR;
     else
        next_tap_state = TAP_SHIFT_DR;
      end
      TAP_UPDATE_DR: begin
     if (tms)
        next_tap_state = TAP_SEL_DR;
     else
        next_tap_state = TAP_TEST;
      end
      TAP_SEL_IR: begin
     if (tms)
        next_tap_state = TAP_RESET;
     else
        next_tap_state = TAP_CAP_IR;
      end
      TAP_CAP_IR: begin
     if (tms)
        next_tap_state = TAP_EXIT1_IR;
     else
        next_tap_state = TAP_SHIFT_IR;
      end
      TAP_SHIFT_IR:  begin
     if (tms)
        next_tap_state = TAP_EXIT1_IR;
     else
        next_tap_state = TAP_SHIFT_IR;
      end
      TAP_EXIT1_IR:  begin
     if (tms)
        next_tap_state = TAP_UPDATE_IR;
     else
        next_tap_state = TAP_PAUSE_IR;
      end
      TAP_PAUSE_IR:  begin
     if (tms)
        next_tap_state = TAP_EXIT2_IR;
     else
        next_tap_state = TAP_PAUSE_IR;
      end
      TAP_EXIT2_IR:  begin
     if (tms)
        next_tap_state = TAP_UPDATE_IR;
     else
        next_tap_state = TAP_SHIFT_IR;
      end
      TAP_UPDATE_IR: begin
     if (tms)
        next_tap_state = TAP_SEL_DR;
     else
        next_tap_state = TAP_TEST;
      end
      default: next_tap_state = {TAP_STATE_WIDTH{1'bx}};
   endcase
end
assign capture_dr_state     = tap_state[TAP_CAP_DR_BIT];
assign shift_dr_state       = tap_state[TAP_SHIFT_DR_BIT];
assign pause_dr_state       = tap_state[TAP_PAUSE_DR_BIT];
assign update_dr_state      = tap_state[TAP_UPDATE_DR_BIT];
assign update_ir_state      = tap_state[TAP_UPDATE_IR_BIT];
assign shift_exit2_dr_state = tap_state[TAP_SHIFT_DR_BIT] | tap_state[TAP_EXIT2_DR_BIT];
always @ ( new_instructions or tap_state or tdi) begin
   if (tap_state[TAP_CAP_IR_BIT])       
      next_new_instructions = { {18-1{1'b0}}, 1'b1 };
   else begin
      if (tap_state[TAP_SHIFT_IR_BIT])  
     next_new_instructions = { tdi, new_instructions[18-1:1] };
      else
     next_new_instructions = new_instructions;
   end
end
always @ ( instructions or new_instructions or tap_state) begin
   if (tap_state[TAP_UPDATE_IR_BIT])
      next_instructions = new_instructions;
   else
      next_instructions = instructions;
end
assign next_tap_state_reset_negedge = tap_state[TAP_RESET_BIT];
assign reset_muxed = dft_pin_pscan ? 1'b0 : tap_state_reset_negedge;
assign instructions_rst_l = ~reset_muxed & trst_n;
assign tdi_ff_en    = tap_state[TAP_SHIFT_DR_BIT];
assign tdi_ff_rst_l = ~(bypass_sel & tap_state[TAP_CAP_DR_BIT]);
assign next_tdo_en = tap_state[TAP_SHIFT_IR_BIT] | tap_state[TAP_SHIFT_DR_BIT];
always @ ( bypass_sel or new_instructions or so
      or tap_state or tdi_ff) begin
   if (tap_state[TAP_SHIFT_IR_BIT])
      next_tdo = new_instructions[0];
   else if (bypass_sel)
      next_tdo = tdi_ff;
   else
      next_tdo = so;
end
assign next_capture_shift_dr = tap_state[TAP_SHIFT_DR_BIT] | tap_state[TAP_CAP_DR_BIT];
assign clock_dr              = tck & capture_shift_dr;
dff_ns #(1) u_dffsl_tap_state_reset_negedge
   ( .din (next_tap_state_reset_negedge),
     .clk (tck_l),
     .q (tap_state_reset_negedge)
     );
dffsl_async_ns #(1) u_dffsl_tap_state0
   ( .din (next_tap_state[0]),
     .clk (tck),
     .set_l (trst_n),
     .q (tap_state[0])
     );
dffrl_async_ns #(TAP_STATE_WIDTH-1) u_dffrl_async_tap_state 
   ( .din (next_tap_state[TAP_STATE_WIDTH-1:1]),
     .clk (tck),
     .rst_l (trst_n),
     .q (tap_state[TAP_STATE_WIDTH-1:1])
     );
dffsl_async_ns #(1) u_dffsl_new_instructions0
   ( .din (next_new_instructions[0]),
     .clk (tck),
     .set_l (trst_n),
     .q (new_instructions[0])
     );
dffrl_async_ns #(18-1) u_dffrl_async_new_instructions 
   ( .din (next_new_instructions[18-1:1]),
     .clk (tck),
     .rst_l (trst_n),
     .q (new_instructions[18-1:1])
     );
dffsl_async_ns #(1) u_dffsl_instructions0
   ( .din (next_instructions[0]),
     .clk (tck_l),
     .set_l (instructions_rst_l),
     .q (instructions[0])
     );
dffrl_async_ns #(18-1) u_dffrl_async_instructions 
   ( .din (next_instructions[18-1:1]),
     .clk (tck_l),
     .rst_l (instructions_rst_l),
     .q (instructions[18-1:1])
     );
dffrl_async_ns #(1) u_dffrl_async_capture_shift_dr 
   ( .din (next_capture_shift_dr),
     .clk (tck_l),
     .rst_l (trst_n),
     .q (capture_shift_dr)
     );
dffrl_async_ns #(1) u_dffrl_async_tdo 
   ( .din (next_tdo),
     .clk (tck_l),
     .rst_l (trst_n),
     .q (tdo)
     );
dffrl_async_ns #(1) u_dffrl_async_tdo_en 
   ( .din (next_tdo_en),
     .clk (tck_l),
     .rst_l (trst_n),
     .q (tdo_en)
     );
dffrle_ns #(1) u_dffrle_tdi_ff
   ( .din (tdi),
     .clk (tck),
     .en (tdi_ff_en),
     .rst_l (tdi_ff_rst_l),
     .q (tdi_ff)
     );
endmodule
  
          
      
    
         
module jtag_ctap(
    input wire clk,
    input wire rst_n,
    
    input wire [128-1:0] jtag_ctap_data,
    input wire jtag_ctap_reg_wr_en,
    input wire [4-1:0] jtag_ctap_reg_sel,
    output reg [128-1:0] ctap_jtag_data,
    output reg ctap_jtag_interrupt_bit,
    
    output reg ctap_ucb_tx_val,
    output reg [128-1:0] ctap_ucb_tx_data,
    output reg [(128/4)-1:0] ctap_ucb_tx_data_vec,
    
    
    input wire ctap_ucb_rx_val,
    input wire [128-1:0] ctap_ucb_rx_data,
    output reg ctap_oram_req_val,
    output reg [4-1:0] ctap_oram_req_misc,
    input wire [64-1:0] oram_ctap_res_data,
    
    
    
    output reg [127:0] ctap_clk_en,
    output reg ctap_oram_clk_en
    );
reg [32-1:0] jtag_req;
reg [32-1:0] jtag_req_misc;
reg [32-1:0] jtag_req_next;
reg jtag_req_val;
reg jtag_req_val_next;
reg [128-1:0] data_reg;
reg [128-1:0] data_reg_next;
reg [32-1:0] jtag_address;
reg [32-1:0] jtag_address_next;
reg interrupt_bit;
reg interrupt_bit_next;
reg response_interrupt_en;
reg clear_interrupt_en;
reg capture_ucb_data_en;
reg [127:0] ctap_clk_en_reg;
reg [127:0] ctap_clk_en_reg_next;
reg ctap_oram_clk_en_reg;
reg ctap_oram_clk_en_reg_next;
reg [128-1:0] rtap_packet;
reg rtap_val;
reg capture_oram_response;
reg capture_oram_response_next;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        jtag_req <= 0;
        data_reg <= 0;
        jtag_address <= 0;
        interrupt_bit <= 0;
        jtag_req_val <= 0;
        capture_oram_response <= 0;
        ctap_clk_en_reg <= ~(128'b0);
        ctap_oram_clk_en_reg <= 1'b0; 
    end
    else
    begin
        jtag_req <= jtag_req_next;
        data_reg <= data_reg_next;
        jtag_address <= jtag_address_next;
        interrupt_bit <= interrupt_bit_next;
        jtag_req_val <= jtag_req_val_next;
        capture_oram_response <= capture_oram_response_next;
        ctap_clk_en_reg <= ctap_clk_en_reg_next;
        ctap_oram_clk_en_reg <= ctap_oram_clk_en_reg_next;
    end
end
reg data_reg_wr_en;
reg inst_wr_en;
reg addr_wr_en;
always @ *
begin
    data_reg_wr_en = 0;
    inst_wr_en = 0;
    addr_wr_en = 0;
    if (jtag_ctap_reg_wr_en)
    begin
        if (jtag_ctap_reg_sel == 4'd1)
            data_reg_wr_en = 1'b1;
        if (jtag_ctap_reg_sel == 4'd2)
            inst_wr_en = 1'b1;
        if (jtag_ctap_reg_sel == 4'd3)
            addr_wr_en = 1'b1;
    end
    
    if (data_reg_wr_en)
    begin
        data_reg_next = 0;
        data_reg_next[63:0] = jtag_ctap_data[63:0]; 
    end
    else if (capture_ucb_data_en)
        data_reg_next[128-1:0] = rtap_packet[128-1:0];
    
    
    else if (capture_oram_response)
        data_reg_next = oram_ctap_res_data;
    else
        data_reg_next = data_reg;
    
    if (inst_wr_en)
        jtag_req_next = jtag_ctap_data;
    else
        jtag_req_next = jtag_req;
    
    if (addr_wr_en)
        jtag_address_next = jtag_ctap_data;
    else
        jtag_address_next = jtag_address;
end
reg jtag_ctap_reg_wr_en_d1;
always @ (posedge clk)
begin
    if (!rst_n)
        jtag_ctap_reg_wr_en_d1 <= 1'b0;
    else
        jtag_ctap_reg_wr_en_d1 <= jtag_ctap_reg_wr_en;
end
always @ *
begin
    jtag_req_val_next = 0;
    if (jtag_req_val == 1'b1)
        jtag_req_val_next = 1'b0;
    else
    begin
        if (jtag_ctap_reg_wr_en_d1 == 1'b1 && jtag_ctap_reg_wr_en == 1'b0 && jtag_ctap_reg_sel == 4'd2)
            jtag_req_val_next = 1'b1;
    end
end
reg [128-1:0] ctap_packet;
reg [(128/4)-1:0] ctap_packet_vec;
reg ctap_packet_val;
reg [32-1:0] ctap_header;
reg [32-1:0] ctap_address;
reg [64-1:0] ctap_data;
always @ *
begin
    ctap_packet_vec = 0;
    ctap_packet_val = 0;
    ctap_packet = 0;
    jtag_req_misc = jtag_req[15:0];
    clear_interrupt_en = 1'b0;
    ctap_oram_req_val = 0;
    ctap_oram_req_misc = 0;
    capture_oram_response_next = 0;
    ctap_clk_en_reg_next = ctap_clk_en_reg;
    ctap_oram_clk_en_reg_next = ctap_oram_clk_en_reg;
    if (jtag_req_val)
    begin
        
        ctap_packet_val = 1'b1;
        case (jtag_req[31:24])
            8'd2:
            begin
                clear_interrupt_en = 1'b1;
                ctap_packet_val = 1'b0;
            end
            8'd9:
            begin
                ctap_oram_req_val = 1'b1;
                ctap_oram_req_misc = jtag_req_misc[4-1:0];
                capture_oram_response_next = 1'b1;
                ctap_packet_val = 1'b0;
            end
            8'd12:
            begin
                ctap_clk_en_reg_next = data_reg[127:0];
                ctap_packet_val = 1'b0;
            end
            8'd13:
            begin
                ctap_oram_clk_en_reg_next = data_reg[0];
                ctap_packet_val = 1'b0;
            end
        endcase
    end
    ctap_header[32-1:0] = jtag_req[32-1:0];
    ctap_address[32-1:0] = jtag_address[32-1:0];
    ctap_data = data_reg[64-1:0];
    ctap_packet[31:0] = ctap_header;
    ctap_packet[63:32] = ctap_address;
    ctap_packet[127:64] = ctap_data;
    ctap_packet_vec = 32'hffffffff;
    
end
reg ret_val;
always @ *
begin
    ret_val = rtap_val;
    capture_ucb_data_en = 1'b0;
    response_interrupt_en = 1'b0;
    if (ret_val)
    begin
        response_interrupt_en = 1'b1;
        capture_ucb_data_en = 1'b1;
    end
end
always @ *
begin
    interrupt_bit_next = interrupt_bit;
    if (response_interrupt_en)
        interrupt_bit_next = 1'b1;
    else if (clear_interrupt_en)
        interrupt_bit_next = 1'b0;
    
    ctap_jtag_interrupt_bit = interrupt_bit;
    ctap_clk_en = ctap_clk_en_reg;
    ctap_oram_clk_en = ctap_oram_clk_en_reg;
end
always @ *
begin
    ctap_jtag_data = data_reg;
end
always @ *
begin
    ctap_ucb_tx_val = ctap_packet_val;
    ctap_ucb_tx_data = ctap_packet;
    ctap_ucb_tx_data_vec = ctap_packet_vec;
end
always @ *
begin
    rtap_packet = ctap_ucb_rx_data;
    rtap_val = ctap_ucb_rx_val;
end
    
    
    
endmodule
  
          
      
    
         
module jtag_ucb_receiver(
    input wire clk,
    input wire rst_n,
    
    output reg ctap_ucb_rx_val,
    output reg [128-1:0] ctap_ucb_rx_data,
    
    
    input wire tiles_jtag_ucb_val,
    input wire [4-1:0] tiles_jtag_ucb_data
    
    );
wire tiles_val;
wire [128-1:0] tiles_data;
ucb_bus_in #(4, 128-64) ucb_in_tiles(
    .vld(tiles_jtag_ucb_val),
    .data(tiles_jtag_ucb_data),
    .stall(),
    .clk(clk),
    .rst_l(rst_n),
    .indata_buf_vld(tiles_val),
    .indata_buf(tiles_data),
    .stall_a1(1'b0)
    );
always @ *
begin
    ctap_ucb_rx_val = tiles_val;
    ctap_ucb_rx_data = 4'b0;
    if (tiles_val)
        ctap_ucb_rx_data = tiles_data;
end
endmodule
  
          
      
    
         
module jtag_ucb_transmitter(
    input wire clk,
    input wire rst_n,
    
    input wire ctap_ucb_tx_val,
    input wire [128-1:0] ctap_ucb_tx_data,
    input wire [(128/4)-1:0] ctap_ucb_tx_data_vec,
    
    output wire jtag_tiles_ucb_val,
    output wire [4-1:0] jtag_tiles_ucb_data
    );
ucb_bus_out #(4, 128-64) ucb_out(
    .vld(jtag_tiles_ucb_val),
    .data(jtag_tiles_ucb_data),
    .outdata_buf_busy(),
    .clk(clk),
    .rst_l(rst_n),
    .stall(1'b0),
    .outdata_buf_in(ctap_ucb_tx_data),
    .outdata_vec_in(ctap_ucb_tx_data_vec),
    .outdata_buf_wr(ctap_ucb_tx_val)
    );
endmodule
    
    
    
     
    
    
    
    
    
    
    
    
    
    
    
    
 
module mc_top (
    output                          mc_ui_clk_sync_rst,
    input                           core_ref_clk,
    input   [64-1:0]   mc_flit_in_data,
    input                           mc_flit_in_val,
    output                          mc_flit_in_rdy,
    output  [64-1:0]   mc_flit_out_data,
    output                          mc_flit_out_val,
    input                           mc_flit_out_rdy,
    input                           uart_boot_en,
    
 
    input                           sys_clk,
    output                          ddr_cas_n,
    output                          ddr_ras_n,
    output                          ddr_we_n,
 
    output [15-1:0]   ddr_addr,
    output [3-1:0]     ddr_ba,
    output [1-1:0]     ddr_ck_n,
    output [1-1:0]     ddr_ck_p,
    output [1-1:0]    ddr_cke,
    output                          ddr_reset_n,
    inout  [64-1:0]     ddr_dq,
    inout  [8-1:0]    ddr_dqs_n,
    inout  [8-1:0]    ddr_dqs_p,
    output [1-1:0]     ddr_cs_n,
 
 
 
    output [8-1:0]     ddr_dm,
 
    output [1-1:0]    ddr_odt,
    output                          init_calib_complete_out,
    input                           sys_rst_n
);
reg     [31:0]                      delay_cnt;
reg                                 ui_clk_syn_rst_delayed;
wire                                init_calib_complete;
wire                                afifo_rst_1;
wire                                afifo_rst_2;
 wire                               app_en;
 wire    [3-1 :0]  app_cmd;
 wire    [29-1:0]  app_addr;
 wire                               app_rdy;
 wire                               app_wdf_wren;
 wire    [512-1:0]  app_wdf_data;
 wire    [64-1:0]  app_wdf_mask;
 wire                               app_wdf_rdy;
 wire                               app_wdf_end;
 wire    [512-1:0]  app_rd_data;
 wire                               app_rd_data_end;
 wire                               app_rd_data_valid;
 wire                               core_app_en;
 wire    [3-1 :0]  core_app_cmd;
 wire    [29-1:0]  core_app_addr;
 wire                               core_app_rdy;
 wire                               core_app_wdf_wren;
 wire    [512-1:0]  core_app_wdf_data;
 wire    [64-1:0]  core_app_wdf_mask;
 wire                               core_app_wdf_rdy;
 wire                               core_app_wdf_end;
 wire    [512-1:0]  core_app_rd_data;
 wire                               core_app_rd_data_end;
 wire                               core_app_rd_data_valid;
wire                                noc_mig_bridge_rst;
wire                                noc_mig_bridge_init_done;
 
wire                                app_sr_req;
wire                                app_ref_req;
wire                                app_zq_req;
wire                                app_sr_active;
wire                                app_ref_ack;
wire                                app_zq_ack;
wire                                ui_clk;
wire                                ui_clk_sync_rst;
wire                                trans_fifo_val;
wire    [64-1:0]       trans_fifo_data;
wire                                trans_fifo_rdy;
wire                                fifo_trans_val;
wire    [64-1:0]       fifo_trans_data;
wire                                fifo_trans_rdy;
reg                                 afifo_ui_rst_r;
reg                                 afifo_ui_rst_r_r;
reg                                 ui_clk_sync_rst_r;
reg                                 ui_clk_sync_rst_r_r;
always @(posedge core_ref_clk) begin
    if (~sys_rst_n)
        delay_cnt <= 32'h1ff;
    else begin
        delay_cnt <= (delay_cnt != 0) & ~ui_clk_sync_rst_r_r ? delay_cnt - 1 : delay_cnt;
    end
end
always @(posedge core_ref_clk) begin
    if (ui_clk_sync_rst)
        ui_clk_syn_rst_delayed <= 1'b1;
    else begin
        ui_clk_syn_rst_delayed <= delay_cnt != 0;
    end
end
assign mc_ui_clk_sync_rst   = ui_clk_syn_rst_delayed;
assign afifo_rst_1 = ui_clk_syn_rst_delayed;
always @(posedge ui_clk) begin
    afifo_ui_rst_r <= afifo_rst_1;
    afifo_ui_rst_r_r <= afifo_ui_rst_r;
end
always @(posedge core_ref_clk) begin
    ui_clk_sync_rst_r   <= ui_clk_sync_rst;
    ui_clk_sync_rst_r_r <= ui_clk_sync_rst_r;
end
assign afifo_rst_2 = afifo_ui_rst_r_r | ui_clk_sync_rst;
assign app_ref_req = 1'b0;
assign app_sr_req = 1'b0;
assign app_zq_req = 1'b0;
assign app_en                   = core_app_en;
assign app_cmd                  = core_app_cmd;
assign app_addr                 = core_app_addr;
assign app_wdf_wren             = core_app_wdf_wren;
assign app_wdf_data             = core_app_wdf_data;
assign app_wdf_mask             = core_app_wdf_mask;
assign app_wdf_end              = core_app_wdf_end;
assign noc_mig_bridge_rst       = ui_clk_sync_rst;
assign noc_mig_bridge_init_done = init_calib_complete;
assign init_calib_complete_out  = init_calib_complete & ~ui_clk_syn_rst_delayed;
assign core_app_rdy             = app_rdy;
assign core_app_wdf_rdy         = app_wdf_rdy;
assign core_app_rd_data_valid   = app_rd_data_valid;
assign core_app_rd_data_end     = app_rd_data_end;
assign core_app_rd_data         = app_rd_data;
noc_bidir_afifo  mig_afifo  (
    .clk_1           (core_ref_clk      ),
    .rst_1           (afifo_rst_1       ),
    .clk_2           (ui_clk            ),
    .rst_2           (afifo_rst_2       ),
    
    .flit_in_val_1   (mc_flit_in_val    ),
    .flit_in_data_1  (mc_flit_in_data   ),
    .flit_in_rdy_1   (mc_flit_in_rdy    ),
    .flit_out_val_2  (fifo_trans_val    ),
    .flit_out_data_2 (fifo_trans_data   ),
    .flit_out_rdy_2  (fifo_trans_rdy    ),
    
    .flit_in_val_2   (trans_fifo_val    ),
    .flit_in_data_2  (trans_fifo_data   ),
    .flit_in_rdy_2   (trans_fifo_rdy    ),
    .flit_out_val_1  (mc_flit_out_val   ),
    .flit_out_data_1 (mc_flit_out_data  ),
    .flit_out_rdy_1  (mc_flit_out_rdy   )
);
assign app_en                   = core_app_en;
assign app_cmd                  = core_app_cmd;
assign app_addr                 = core_app_addr;
assign app_wdf_wren             = core_app_wdf_wren;
assign app_wdf_data             = core_app_wdf_data;
assign app_wdf_mask             = core_app_wdf_mask;
assign app_wdf_end              = core_app_wdf_end;
assign noc_mig_bridge_rst       = ui_clk_sync_rst;
assign noc_mig_bridge_init_done = init_calib_complete;
assign init_calib_complete_out  = init_calib_complete & ~ui_clk_syn_rst_delayed;
assign core_app_rdy             = app_rdy;
assign core_app_wdf_rdy         = app_wdf_rdy;
assign core_app_rd_data_valid   = app_rd_data_valid;
assign core_app_rd_data_end     = app_rd_data_end;
assign core_app_rd_data         = app_rd_data;
noc_mig_bridge    #  (
    .MIG_APP_ADDR_WIDTH (29        ),
    .MIG_APP_DATA_WIDTH (512        )
)   noc_mig_bridge   (
    .clk                (ui_clk                     ),  
    .rst                (noc_mig_bridge_rst         ),  
    .uart_boot_en       (uart_boot_en               ),
    .flit_in            (fifo_trans_data            ),
    .flit_in_val        (fifo_trans_val             ),
    .flit_in_rdy        (fifo_trans_rdy             ),
    .flit_out           (trans_fifo_data            ),
    .flit_out_val       (trans_fifo_val             ),
    .flit_out_rdy       (trans_fifo_rdy             ),
    .app_rdy            (core_app_rdy               ),
    .app_wdf_rdy        (core_app_wdf_rdy           ),
    .app_rd_data        (core_app_rd_data           ),
    .app_rd_data_end    (core_app_rd_data_end       ),
    .app_rd_data_valid  (core_app_rd_data_valid     ),
    .phy_init_done      (noc_mig_bridge_init_done   ),
    .app_wdf_wren_reg   (core_app_wdf_wren          ),
    .app_wdf_data_out   (core_app_wdf_data          ),
    .app_wdf_mask_out   (core_app_wdf_mask          ),
    .app_wdf_end_out    (core_app_wdf_end           ),
    .app_addr_out       (core_app_addr              ),
    .app_en_reg         (core_app_en                ),
    .app_cmd_reg        (core_app_cmd               )
);
 
                        
 
mig_7series_0   mig_7series_0 (
    
    .ddr3_addr                      (ddr_addr),
    .ddr3_ba                        (ddr_ba),
    .ddr3_cas_n                     (ddr_cas_n),
    .ddr3_ck_n                      (ddr_ck_n),
    .ddr3_ck_p                      (ddr_ck_p),
    .ddr3_cke                       (ddr_cke),
    .ddr3_ras_n                     (ddr_ras_n),
    .ddr3_reset_n                   (ddr_reset_n),
    .ddr3_we_n                      (ddr_we_n),
    .ddr3_dq                        (ddr_dq),
    .ddr3_dqs_n                     (ddr_dqs_n),
    .ddr3_dqs_p                     (ddr_dqs_p),
    .ddr3_cs_n                      (ddr_cs_n),
 
    .ddr3_dm                        (ddr_dm),
    .ddr3_odt                       (ddr_odt),
 
    .init_calib_complete            (init_calib_complete),
    
    .app_addr                       (app_addr),
    .app_cmd                        (app_cmd),
    .app_en                         (app_en),
    .app_wdf_data                   (app_wdf_data),
    .app_wdf_end                    (app_wdf_end),
    .app_wdf_wren                   (app_wdf_wren),
    .app_rd_data                    (app_rd_data),
    .app_rd_data_end                (app_rd_data_end),
    .app_rd_data_valid              (app_rd_data_valid),
    .app_rdy                        (app_rdy),
    .app_wdf_rdy                    (app_wdf_rdy),
    .app_sr_req                     (app_sr_req),
    .app_ref_req                    (app_ref_req),
    .app_zq_req                     (app_zq_req),
    .app_sr_active                  (app_sr_active),
    .app_ref_ack                    (app_ref_ack),
    .app_zq_ack                     (app_zq_ack),
    .ui_clk                         (ui_clk),
    .ui_clk_sync_rst                (ui_clk_sync_rst),
    .app_wdf_mask                   (app_wdf_mask),
    
    .sys_clk_i                      (sys_clk),
    .sys_rst                        (sys_rst_n)
);
 
 
 
 
                        
 
 
  
  
  
endmodule 
    
    
    
     
    
    
    
    
    
    
    
    
    
    
    
    
module memory_zeroer
#(
    parameter MIG_APP_ADDR_WIDTH          = 28,
    parameter MIG_APP_DATA_WIDTH          = 128, 
    parameter MIG_APP_MASK_WIDTH          = MIG_APP_DATA_WIDTH / 8
)
(
    input   clk,
    input   rst_n,
    input   init_calib_complete_in,
    output  init_calib_complete_out,
    
    input                           app_rdy_in,
    input                           app_wdf_rdy_in,
    input                           app_wdf_wren_in,
    input [MIG_APP_DATA_WIDTH-1:0]  app_wdf_data_in,
    input [MIG_APP_MASK_WIDTH-1:0]  app_wdf_mask_in,
    input                           app_wdf_end_in,
    input [MIG_APP_ADDR_WIDTH-1:0]  app_addr_in,
    input                           app_en_in,
    input [2:0]                     app_cmd_in,
    output                          app_wdf_wren_out,
    output [MIG_APP_DATA_WIDTH-1:0] app_wdf_data_out,
    output [MIG_APP_MASK_WIDTH-1:0] app_wdf_mask_out,
    output                          app_wdf_end_out,
    output [MIG_APP_ADDR_WIDTH-1:0] app_addr_out,
    output                          app_en_out,
    output [2:0]                    app_cmd_out
);
localparam reg [63:0] BOARD_MEM_SIZE_MB = 1024;
localparam reg [63:0] MAX_MEM_ADDR      = (BOARD_MEM_SIZE_MB * 2**20) / 8;
localparam reg [63:0] WORDS_PER_WR      = 8;
wire                          app_wdf_wren;
wire [MIG_APP_DATA_WIDTH-1:0] app_wdf_data;
wire [MIG_APP_MASK_WIDTH-1:0] app_wdf_mask;
wire                          app_wdf_end;
wire [MIG_APP_ADDR_WIDTH-1:0] app_addr;
wire                          app_en;
wire [2:0]                    app_cmd;
wire zeroing_done;
reg [MIG_APP_ADDR_WIDTH:0] address_f;
wire [MIG_APP_ADDR_WIDTH:0] address_next;
reg  [7:0] extra_time_f;
wire [7:0] extra_time_next;
wire extra_time_done;
assign address_next = (init_calib_complete_in & app_rdy_in & app_wdf_rdy_in & (address_f <= MAX_MEM_ADDR)) ? address_f + WORDS_PER_WR : address_f;
always @(posedge clk)
begin
    if (~rst_n)
    begin
        address_f <= {MIG_APP_ADDR_WIDTH+1{1'b0}};
        extra_time_f <= 8'b11111111;
    end
    else
    begin
        address_f <= address_next;
        extra_time_f <= extra_time_next;
    end
end
assign zeroing_done = (address_f >= MAX_MEM_ADDR);
assign extra_time_next = ((~zeroing_done) | (extra_time_f == 8'b0)) ? extra_time_f : (extra_time_f - 1'b1);
assign extra_time_done = zeroing_done & (extra_time_f == 8'b0);
assign init_calib_complete_out = init_calib_complete_in & extra_time_done;
assign app_wdf_wren = 1'b1 & app_rdy_in & app_wdf_rdy_in;
assign app_wdf_wren_out = zeroing_done ? app_wdf_wren_in : app_wdf_wren;
assign app_wdf_data = {MIG_APP_DATA_WIDTH{1'b0}};
assign app_wdf_data_out = zeroing_done ? app_wdf_data_in : app_wdf_data;
assign app_wdf_mask = {MIG_APP_MASK_WIDTH{1'b0}};
assign app_wdf_mask_out = zeroing_done ? app_wdf_mask_in : app_wdf_mask;
assign app_wdf_end = 1'b1;
assign app_wdf_end_out = zeroing_done ? app_wdf_end_in : app_wdf_end;
assign app_addr = address_f[MIG_APP_ADDR_WIDTH-1:0];
assign app_addr_out = zeroing_done ? app_addr_in : app_addr;
assign app_en = 1'b1 & app_rdy_in & app_wdf_rdy_in;
assign app_en_out = zeroing_done ? app_en_in : app_en;
assign app_cmd = 3'b000;
assign app_cmd_out = zeroing_done ? app_cmd_in : app_cmd;
endmodule
    
    
    
     
    
    
    
    
    
    
    
    
    
    
    
    
module noc_mig_bridge # (
  parameter MIG_APP_ADDR_WIDTH          = 28,
  parameter MIG_APP_DATA_WIDTH          = 128, 
  parameter MIG_APP_MASK_WIDTH          = MIG_APP_DATA_WIDTH / 8,
  parameter IN_FLIGHT_LIMIT             = 16, 
  parameter BUFFER_ADDR_SIZE            = 4 
)
(
  input                             clk,
  input                             rst,
   
   input                                uart_boot_en,
  
   input       [64-1:0]           flit_in,
   input                                 flit_in_val,
   output                                flit_in_rdy,
   output      [64-1:0]           flit_out,
   output                                flit_out_val,
   input                                 flit_out_rdy,
  
   input                                 app_rdy,
   input                                 app_wdf_rdy,
   input       [MIG_APP_DATA_WIDTH-1:0]  app_rd_data,
   input                                 app_rd_data_end,
   input                                 app_rd_data_valid,
   input                                 phy_init_done,
   output reg                            app_wdf_wren_reg,
   output      [MIG_APP_DATA_WIDTH-1:0]  app_wdf_data_out,
   output      [MIG_APP_MASK_WIDTH-1:0]  app_wdf_mask_out,
   output                                app_wdf_end_out,
   output      [MIG_APP_ADDR_WIDTH-1:0]  app_addr_out,
   output reg                            app_en_reg,
   output reg  [2:0]                     app_cmd_reg
);
localparam CL_ADDR_WIDTH = 40 - 6;
localparam APP_DATA_WIDTH              = 512; 
localparam APP_MASK_WIDTH              = APP_DATA_WIDTH / 8;   
localparam MAX_PKT_LEN                 = 11; 
localparam MAX_PKT_LEN_LOG             = clogb2(MAX_PKT_LEN);
localparam LOC_ADDR_HI                 = (16 + 40 - 1);
localparam LOC_ADDR_LO                 = 16 + 6;
localparam RATIO        = APP_DATA_WIDTH / MIG_APP_DATA_WIDTH;  
localparam RATIO_WIDTH  = clogb2(RATIO);
localparam WORD_SIZE_LOG = clogb2(8);
integer i;
reg [64-1:0]           pkt_w1        [IN_FLIGHT_LIMIT-1:0];
reg [64-1:0]           pkt_w2        [IN_FLIGHT_LIMIT-1:0];
reg [64-1:0]           pkt_w3        [IN_FLIGHT_LIMIT-1:0]; 
reg [APP_DATA_WIDTH-1:0]  pkt_data_buf  [IN_FLIGHT_LIMIT-1:0];
 reg [2:0]                     pkt_state_buf [IN_FLIGHT_LIMIT-1:0];
 reg [8-1:0]   pkt_cmd_buf   [IN_FLIGHT_LIMIT-1:0];
reg [64-1:0]           in_data_buf[MAX_PKT_LEN-4:0]; 
reg [BUFFER_ADDR_SIZE-1:0]    buf_current_in;  
reg [BUFFER_ADDR_SIZE-1:0]    buf_current_out; 
reg [MAX_PKT_LEN_LOG-1:0]     remaining_flits; 
reg [2:0]                     acc_state;
reg [BUFFER_ADDR_SIZE-1:0]    buf_current_cmd;  
reg                           r_app_en;         
reg [BUFFER_ADDR_SIZE-1:0]    buf_current_data_rcv;
reg [MAX_PKT_LEN_LOG-1:0]     remaining_flt_out;
reg [64-1:0]           flit_out_buffer[MAX_PKT_LEN-1:0];
reg [BUFFER_ADDR_SIZE-1:0]    buf_current_wdf; 
reg                           buf_wdf_data_half;  
reg                           r_app_wdf_wren;     
wire                        app_wdf_wren;
wire  [APP_DATA_WIDTH-1:0]  app_wdf_data;
wire  [APP_MASK_WIDTH-1:0]  app_wdf_mask;
wire                        app_wdf_end;
wire  [CL_ADDR_WIDTH-1:0]   cl_addr;
wire                        app_en;
wire  [2:0]                 app_cmd;
reg                        app_wdf_wren_r;
reg  [APP_DATA_WIDTH-1:0]  app_wdf_data_r;
reg  [APP_MASK_WIDTH-1:0]  app_wdf_mask_r;
reg                        app_wdf_end_r;
reg                        app_wdf_wren_r_r;
reg  [APP_DATA_WIDTH-1:0]  app_wdf_data_r_r;
reg  [APP_MASK_WIDTH-1:0]  app_wdf_mask_r_r;
reg                        app_wdf_end_r_r;
reg       [APP_DATA_WIDTH-1:0]  app_rd_data_reg;
reg                             app_rd_data_end_reg;
reg                             app_rd_data_valid_reg;
reg       [CL_ADDR_WIDTH-1:0]      cl_addr_reg;
reg      [APP_DATA_WIDTH-1:0]   app_wdf_data_reg;
reg      [APP_MASK_WIDTH-1:0]   app_wdf_mask_reg;
reg                             app_wdf_end_reg;
reg   [5:0]     cmd_part;
reg             cmd_pending;
reg             wdf_pending;
reg   [5:0]     wdf_part;
reg   [5:0]     rd_part;
wire            cmd_send_end;
wire  [5:0]     cmd_part_next;
wire            app_rdy_trans;
wire            wdf_send_end;
wire  [5:0]     wdf_part_next;
wire            app_wdf_rdy_trans;
wire            rd_last;
wire  [5:0]     rd_part_next;
wire  [MIG_APP_DATA_WIDTH-1:0]  wdf_data_part [RATIO-1:0];
wire  [MIG_APP_MASK_WIDTH-1:0]  wdf_mask_part [RATIO-1:0];
reg   [MIG_APP_DATA_WIDTH-1:0]  app_rd_data_part [RATIO-1:0];
wire  [APP_DATA_WIDTH-1:0]      app_rd_data_trans;
always @(posedge clk) begin
  app_rd_data_reg       <= app_rd_data_trans;
  app_rd_data_end_reg   <= rd_last;
  app_rd_data_valid_reg <= rd_last;
end
assign flit_in_rdy  = (acc_state != 4 && !rst && phy_init_done);
always @(posedge clk) begin
  if(rst) begin
    
    buf_current_in <= 0;
    remaining_flits <= 0;
    acc_state = 0;
    
    for(i=0; i < IN_FLIGHT_LIMIT; i=i+1) begin
      pkt_w1        [i] <= 0;
      pkt_w2        [i] <= 0;
      pkt_w3        [i] <= 0;
      
      pkt_cmd_buf   [i] <= 0;
      
    end
    for(i=0; i < MAX_PKT_LEN-3; i = i + 1) begin
      in_data_buf[i] <= 0;
    end
  end
  else begin
    if(flit_in_val) begin
      
      case (acc_state) 
      
      0: begin 
        
        pkt_w1        [buf_current_in] <= flit_in;
        pkt_cmd_buf   [buf_current_in] <= flit_in[21:14];
        remaining_flits <= flit_in[29:22]-1;    
        acc_state       <= 1;
      end
      
      1: begin
        pkt_w2        [buf_current_in] <= flit_in;  
        remaining_flits <= remaining_flits-1;
        acc_state <= 2;
      end
      
      2: begin
        pkt_w3        [buf_current_in] <= flit_in;
        
        if(remaining_flits == 0) begin 
            
            if(buf_current_in+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}} == buf_current_out) begin
                buf_current_in <= buf_current_in + 1;
                
                acc_state <= 4;
            end
            else begin
                buf_current_in <= buf_current_in + 1;
                
                acc_state <= 0;
            end
        end
        else begin 
            remaining_flits <= remaining_flits-1;
            acc_state <= 3;
        end
      end
      
      3: begin
        in_data_buf[remaining_flits] <= flit_in;
        remaining_flits <= remaining_flits - 1;
        
        if((remaining_flits == 0)) begin
            buf_current_in <= buf_current_in+1;
            if (buf_current_in+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}} != buf_current_out) begin	
                acc_state <= 0;
            end
            else begin
                acc_state <= 4;
            end
        end
      end
      
      4: begin 
        if(buf_current_in != buf_current_out) begin
            
            acc_state <= 0;
        end
      end
      default: begin
        
      end
      endcase
    end
  end
end
generate begin
  genvar ii;
  for (ii = 0; ii < IN_FLIGHT_LIMIT; ii = ii + 1) begin: IN_STATE
    always @(posedge clk) begin
      if(rst) begin
        pkt_data_buf[ii]  <= {APP_DATA_WIDTH{1'b0}};
        pkt_state_buf[ii] <= 5;
      end
      else begin
        pkt_data_buf[ii]  <= (ii == buf_current_in) & flit_in_val &
                             (acc_state == 3) & (remaining_flits == 0)   ?   { flit_in, 
                                                                                        in_data_buf[1], 
                                                                                        in_data_buf[2],
                                                                                        in_data_buf[3],
                                                                                        in_data_buf[4],
                                                                                        in_data_buf[5],
                                                                                        in_data_buf[6],
                                                                                        in_data_buf[7]}   :
                              (ii == buf_current_data_rcv) & app_rd_data_valid_reg  ?   app_rd_data_reg   : 
                                                                                        pkt_data_buf[ii]  ;
        pkt_state_buf[ii] <= (ii == buf_current_in)   & 
                             flit_in_val                              ? ((acc_state == 0)                ?   0          :
                                                                         (acc_state == 2)   & 
                                                                         (remaining_flits == 0)                   ?   2      :
                                                                         (acc_state == 3) &
                                                                         (remaining_flits == 0)                   ?   1      :
                                                                         (acc_state == 4)     &
                                                                         (buf_current_in != buf_current_out)      ?   0          :
                                                                                                                  pkt_state_buf[ii]
                                                                         )                  :
                              (ii == buf_current_out)             & 
                              ((pkt_state_buf[ii] == 4) |
                               (pkt_state_buf[ii] == 5))  &
                              (remaining_flt_out == 0)                ?   5         :
                              (ii == buf_current_data_rcv)        &
                              app_rd_data_valid_reg               & 
                              app_rd_data_end_reg                     ?   4            :
                              (ii == buf_current_cmd)             &
                              app_en & app_rdy_trans                        ? ((pkt_cmd_buf[ii] == 8'd15) |
                                                                         (pkt_cmd_buf[ii] == 8'd20) ?    4            :
                                                                                                                      3     
                                                                        )                   :
                              (ii == buf_current_wdf)             &
                              app_wdf_wren                        &
                              app_wdf_rdy_trans                         &
                              (buf_wdf_data_half == 0)          ?   2      :
                                                                          pkt_state_buf[ii] ;                                                            
      end
    end
  end
end
endgenerate
always @(posedge clk) begin
  app_wdf_wren_r <= app_wdf_rdy_trans ? app_wdf_wren  : app_wdf_wren_r;
  app_wdf_data_r <= app_wdf_rdy_trans ? app_wdf_data  : app_wdf_data_r;
  app_wdf_mask_r <= app_wdf_rdy_trans ? app_wdf_mask  : app_wdf_mask_r;
  app_wdf_end_r  <= app_wdf_rdy_trans ? app_wdf_end   : app_wdf_end_r;
end
always @(posedge clk) begin
  app_wdf_wren_r_r <= app_wdf_rdy_trans   ? app_wdf_wren_r  : app_wdf_wren_r_r;
  app_wdf_data_r_r <= app_wdf_rdy_trans   ? app_wdf_data_r  : app_wdf_data_r_r;
  app_wdf_mask_r_r <= app_wdf_rdy_trans   ? app_wdf_mask_r  : app_wdf_mask_r_r;
  app_wdf_end_r_r  <= app_wdf_rdy_trans   ? app_wdf_end_r   : app_wdf_end_r_r;
end
always @(posedge clk) begin
  if (rst) begin
    app_wdf_wren_reg  <= 1'b0;
    app_wdf_data_reg  <= {APP_DATA_WIDTH{1'b0}};
    app_wdf_mask_reg  <= {APP_MASK_WIDTH{1'b0}};
    app_wdf_end_reg   <= 1'b0;
    app_en_reg        <= 1'b0;
    cl_addr_reg       <= {CL_ADDR_WIDTH{1'b0}};
    app_cmd_reg       <= {3{1'b0}};
  end else begin
    app_wdf_wren_reg  <= app_wdf_rdy_trans      ? app_wdf_wren_r_r : app_wdf_wren_reg;
    app_wdf_data_reg  <= app_wdf_rdy_trans      ? app_wdf_data_r_r : app_wdf_data_reg;
    app_wdf_mask_reg  <= app_wdf_rdy_trans      ? app_wdf_mask_r_r : app_wdf_mask_reg;
    app_wdf_end_reg   <= app_wdf_rdy_trans      ? app_wdf_end_r_r  : app_wdf_end_reg;
    app_en_reg        <= app_rdy_trans    ? app_en       : app_en_reg;
    cl_addr_reg      <= app_rdy_trans    ? cl_addr     : cl_addr_reg;
    app_cmd_reg       <= app_rdy_trans    ? app_cmd      : app_cmd_reg;
  end
end
wire [RATIO_WIDTH-1:0]  last_addr_bits [RATIO-1:0];
wire [RATIO-1:0]        inv_cmp [RATIO_WIDTH-1:0];
wire [RATIO_WIDTH-1:0]  curr_last_bits;
generate begin
  if (RATIO_WIDTH > 0) begin
    assign curr_last_bits = cmd_part[RATIO_WIDTH-1:0];
  end
end
endgenerate
assign cmd_send_end       = app_en_reg & (cmd_part == (RATIO - 1)) & app_rdy;
assign cmd_part_next      = cmd_part == (RATIO - 1) ? 6'b0 : cmd_part + 1;  
assign app_rdy_trans      = (~cmd_pending | cmd_send_end) & ~(app_en_reg & ~cmd_send_end);
always @(posedge clk) begin
  if (rst)
    cmd_pending <= 1'b0;
  else
    cmd_pending <=  app_en_reg & ~cmd_send_end ? 1'b1  :
                    cmd_send_end               ? 1'b0  : cmd_pending;
end
always @(posedge clk) begin
  if (rst)
    cmd_part <= 5'b0;
  else
    cmd_part <= app_en_reg & app_rdy ? cmd_part_next : cmd_part;
end
assign wdf_send_end     = app_wdf_wren_reg & (wdf_part == (RATIO - 1)) & app_wdf_rdy;
assign wdf_part_next    = wdf_part == (RATIO - 1) ? 6'b0 : wdf_part + 1;
assign app_wdf_rdy_trans    = (~wdf_pending | wdf_send_end) & ~(app_wdf_wren_reg & ~wdf_send_end);
always @(posedge clk) begin
  if (rst)
    wdf_pending <= 1'b0;
  else
    wdf_pending <=  app_wdf_wren_reg & ~wdf_send_end  ? 1'b1 :
                    wdf_send_end                      ? 1'b0 : wdf_pending;
end
always @(posedge clk) begin
  if (rst)
    wdf_part  <= 5'b0;
  else
    wdf_part  <= app_wdf_wren_reg & app_wdf_rdy ? wdf_part_next : wdf_part; 
end
generate begin
  genvar ii;
  for (ii = 0; ii < RATIO; ii = ii + 1) begin: APP_WDF
    assign wdf_data_part[ii] = app_wdf_data_reg[(ii+1)*MIG_APP_DATA_WIDTH - 1 : ii*MIG_APP_DATA_WIDTH];
    assign wdf_mask_part[ii] = app_wdf_mask_reg[(ii+1)*MIG_APP_MASK_WIDTH - 1 : ii*MIG_APP_MASK_WIDTH];
  end
end
endgenerate
generate begin
  if (RATIO_WIDTH > 0)
    assign app_addr_out = {cl_addr_reg, curr_last_bits, 3'b0}; 
  else
    assign app_addr_out = {cl_addr_reg, 3'b0};
end
endgenerate
assign app_wdf_data_out = wdf_data_part[wdf_part];
assign app_wdf_mask_out = wdf_mask_part[wdf_part];
assign app_wdf_end_out  = app_wdf_wren_reg;   
assign rd_part_next = rd_part == (RATIO - 1) ? 6'b0 : rd_part + 1;
assign rd_last      = (rd_part == (RATIO-1)) & app_rd_data_valid; 
always @(posedge clk) begin
  if (rst)
    rd_part   <= 5'b0;
  else
    rd_part   <= app_rd_data_valid ? rd_part_next : rd_part;
end
generate begin
  genvar ii;
  for (ii = 0; ii < RATIO; ii = ii + 1) begin: APP_RD
    always @(posedge clk) begin
      app_rd_data_part[ii] <= rd_part == ii ? app_rd_data : app_rd_data_part[ii]; 
    end
    if (ii == (RATIO-1)) 
      assign app_rd_data_trans[(ii+1)*MIG_APP_DATA_WIDTH-1 : ii*MIG_APP_DATA_WIDTH] = app_rd_data;
    else
      assign app_rd_data_trans[(ii+1)*MIG_APP_DATA_WIDTH-1 : ii*MIG_APP_DATA_WIDTH] = app_rd_data_part[ii];
  end
end
endgenerate
assign app_wdf_wren  = (pkt_state_buf[buf_current_wdf] == 1) ? 1'b1 : 1'b0;
assign app_wdf_data  = pkt_data_buf[buf_current_wdf];
assign app_wdf_mask  = {APP_MASK_WIDTH{1'b0}};
assign app_wdf_end   = (buf_wdf_data_half == 0);
assign app_en        = r_app_en;
  
  
wire  [CL_ADDR_WIDTH-1:0]   cl_addr_uart_boot;
wire  [48-1:0]   app_addr_virt;
wire  [29-1:0] storage_addr_out;   
assign app_addr_virt = pkt_w2[buf_current_cmd][((16 + 40 - 1)):(16)];
  storage_addr_trans #(
    .STORAGE_ADDR_WIDTH(29)
  ) cpu_mig_addr_translator (
    .va_byte_addr       (app_addr_virt        ),
    .storage_addr_out   (storage_addr_out     )
  );
  
  
  assign cl_addr_uart_boot   = {storage_addr_out, {WORD_SIZE_LOG{1'b0}}} >> 6;
  assign cl_addr      = uart_boot_en ? cl_addr_uart_boot : 
                                      pkt_w2[buf_current_cmd][LOC_ADDR_HI: LOC_ADDR_LO];  
assign app_cmd       = (pkt_cmd_buf[buf_current_cmd] == 8'd15 ||
                        pkt_cmd_buf[buf_current_cmd] == 8'd20) ? 3'b000 : 3'b001;
always@(posedge clk) begin
  if(rst) begin
    buf_current_wdf <= 0;
    buf_wdf_data_half <= 0;
    r_app_wdf_wren <= 0;
  end
  else begin
    if( (pkt_cmd_buf[buf_current_wdf] == 8'd14 || 
         pkt_cmd_buf[buf_current_wdf] == 8'd19) && 
        (pkt_state_buf[buf_current_wdf] != 5) ) 
    begin  
      buf_current_wdf <= buf_current_wdf + 1;
    end
    r_app_wdf_wren <= (pkt_state_buf[buf_current_wdf] == 1) ? 1 : 0;
    if(app_wdf_wren_r_r && app_wdf_rdy_trans) begin
      buf_current_wdf <= buf_current_wdf + 1;
    end
  end
end
always @(posedge clk) begin
  if(rst) begin
    buf_current_cmd <= 0;
    r_app_en <= 0;
  end
  else begin
    if(pkt_state_buf[buf_current_cmd] == 2) begin
      r_app_en <= 1;
    end
    if (app_en && app_rdy_trans) begin
      r_app_en <= 0;
      buf_current_cmd <= buf_current_cmd+1;
    end
    
  end
end
always @(posedge clk) begin
  if(rst) begin
    buf_current_data_rcv <= 0;
  end
	else begin
		if( (pkt_cmd_buf[buf_current_data_rcv] == 8'd15 || 
             pkt_cmd_buf[buf_current_data_rcv] == 8'd20) && 
            (pkt_state_buf[buf_current_data_rcv][2:0] != 5)) 
    begin 
      buf_current_data_rcv <= buf_current_data_rcv+1;
    end
    if(app_rd_data_valid_reg) begin 
      if (app_rd_data_end_reg) begin
        buf_current_data_rcv <= buf_current_data_rcv+1;
      end
    end
  end
end
assign flit_out = flit_out_buffer[remaining_flt_out-1];
assign flit_out_val = (pkt_state_buf[buf_current_out] == 4) & (remaining_flt_out > 0); 
always @(posedge clk) begin
  if(rst) begin
    buf_current_out <= IN_FLIGHT_LIMIT-1; 
    remaining_flt_out <= 0;
    for(i=0; i < MAX_PKT_LEN; i=i+1) begin
        flit_out_buffer[i] <= 64'h0;
    end
  end
  else begin
    if(pkt_state_buf[buf_current_out] == 4 ||
       pkt_state_buf[buf_current_out] == 5 ) begin
      if (remaining_flt_out == 0) begin
        
        if(pkt_state_buf[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}] == 4 ) begin
            buf_current_out <= buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}};
            
            if( pkt_cmd_buf[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}] == 8'd14 || 
                pkt_cmd_buf[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}] == 8'd19
                ) begin 
                remaining_flt_out <= 9;   
                
                flit_out_buffer[8][63:50  ]     <= pkt_w3[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}][63:50 ];
                flit_out_buffer[8][49:42       ]     <= pkt_w3[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}][49:42      ];
                flit_out_buffer[8][41:34       ]     <= pkt_w3[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}][41:34      ];
                flit_out_buffer[8][33:30   ]     <= pkt_w3[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}][33:30  ];
                flit_out_buffer[8][13:6      ]     <= pkt_w1[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}][13:6      ];
                flit_out_buffer[8][29:22] <= MAX_PKT_LEN-3;    
                
                if(pkt_cmd_buf[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}] == 8'd14) begin
                  flit_out_buffer[8][21:14] <=  8'd26; 
                end
                if(pkt_cmd_buf[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}] == 8'd19) begin
                  flit_out_buffer[8][21:14] <=  8'd24; 
                end 
        
                
                flit_out_buffer[8][5:0] <= {6{1'b0}};
                
                
                
                flit_out_buffer[0]  <= pkt_data_buf[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}][((8)*64)-1:(7)*64];
                flit_out_buffer[1]  <= pkt_data_buf[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}][((7)*64)-1:(6)*64];
                flit_out_buffer[2]  <= pkt_data_buf[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}][((6)*64)-1:(5)*64];
                flit_out_buffer[3]  <= pkt_data_buf[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}][((5)*64)-1:(4)*64];
                flit_out_buffer[4]  <= pkt_data_buf[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}][((4)*64)-1:(3)*64];
                flit_out_buffer[5]  <= pkt_data_buf[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}][((3)*64)-1:(2)*64];
                flit_out_buffer[6]  <= pkt_data_buf[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}][((2)*64)-1:(1)*64];
                flit_out_buffer[7]  <= pkt_data_buf[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}][((1)*64)-1:(0)*64];
            end
            else begin 
                flit_out_buffer[0][29:22] <= 0; 
                remaining_flt_out <= 1;
                flit_out_buffer[0][63:50  ] <= pkt_w3[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}][63:50 ];
                flit_out_buffer[0][49:42       ] <= pkt_w3[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}][49:42      ];
                flit_out_buffer[0][41:34       ] <= pkt_w3[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}][41:34      ];
                flit_out_buffer[0][33:30   ] <= pkt_w3[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}][33:30  ];
                flit_out_buffer[0][13:6      ] <= pkt_w1[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}][13:6      ];
                if(pkt_cmd_buf[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}] == 8'd15) begin
                  flit_out_buffer[0][21:14] <=  8'd27; 
                end
                if(pkt_cmd_buf[buf_current_out+{{BUFFER_ADDR_SIZE-1{1'b0}}, {1'b1}}] == 8'd20) begin
                  flit_out_buffer[0][21:14] <=  8'd25; 
                end
                
                flit_out_buffer[0][5:0] <= {6{1'b0}};
            end
         end
      end
      else begin
        if(flit_out_rdy && flit_out_val) begin
          remaining_flt_out <= remaining_flt_out-1;
        end
      end
    end
  end
end
function integer clogb2;
    input [31:0] value;
    begin
        value = value - 1;
        for (clogb2 = 0; value > 0; clogb2 = clogb2 + 1) begin
            value = value >> 1;
        end
    end
endfunction
endmodule
    
    
    
     
    
    
    
    
    
    
    
    
    
    
    
    
 
module f1_mc_top (
    input                           sys_clk,       
    input                           sys_rst_n,     
    input                           mc_clk,
    input   [64-1:0]   mc_flit_in_data,
    input                           mc_flit_in_val,
    output                          mc_flit_in_rdy,
    output  [64-1:0]   mc_flit_out_data,
    output                          mc_flit_out_val,
    input                           mc_flit_out_rdy,
    input                           uart_boot_en,
    output                          init_calib_complete_out,
    output                          mc_ui_clk_sync_rst,
    
    output wire [6     -1:0]    m_axi_awid,
    output wire [64   -1:0]    m_axi_awaddr,
    output wire [8    -1:0]    m_axi_awlen,
    output wire [3   -1:0]    m_axi_awsize,
    output wire [2  -1:0]    m_axi_awburst,
    output wire                                  m_axi_awlock,
    output wire [4  -1:0]    m_axi_awcache,
    output wire [3   -1:0]    m_axi_awprot,
    output wire [4    -1:0]    m_axi_awqos,
    output wire [4 -1:0]    m_axi_awregion,
    output wire [11   -1:0]    m_axi_awuser,
    output wire                                  m_axi_awvalid,
    input  wire                                  m_axi_awready,
    
    output wire  [6     -1:0]    m_axi_wid,
    output wire  [512   -1:0]    m_axi_wdata,
    output wire  [64   -1:0]    m_axi_wstrb,
    output wire                                   m_axi_wlast,
    output wire  [11   -1:0]    m_axi_wuser,
    output wire                                   m_axi_wvalid,
    input  wire                                   m_axi_wready,
    
    output wire  [6     -1:0]    m_axi_arid,
    output wire  [64   -1:0]    m_axi_araddr,
    output wire  [8    -1:0]    m_axi_arlen,
    output wire  [3   -1:0]    m_axi_arsize,
    output wire  [2  -1:0]    m_axi_arburst,
    output wire                                   m_axi_arlock,
    output wire  [4  -1:0]    m_axi_arcache,
    output wire  [3   -1:0]    m_axi_arprot,
    output wire  [4    -1:0]    m_axi_arqos,
    output wire  [4 -1:0]    m_axi_arregion,
    output wire  [11   -1:0]    m_axi_aruser,
    output wire                                   m_axi_arvalid,
    input  wire                                   m_axi_arready,
    
    input  wire  [6     -1:0]    m_axi_rid,
    input  wire  [512   -1:0]    m_axi_rdata,
    input  wire  [2   -1:0]    m_axi_rresp,
    input  wire                                   m_axi_rlast,
    input  wire  [11   -1:0]    m_axi_ruser,
    input  wire                                   m_axi_rvalid,
    output wire                                   m_axi_rready,
    
    input  wire  [6     -1:0]    m_axi_bid,
    input  wire  [2   -1:0]    m_axi_bresp,
    input  wire  [11   -1:0]    m_axi_buser,
    input  wire                                   m_axi_bvalid,
    output wire                                   m_axi_bready, 
    input wire                                    ddr_ready
);
reg pre_mc_rst_n;
reg mc_rst_n;
always @(negedge sys_rst_n or posedge mc_clk) begin 
    if(!sys_rst_n) begin
        pre_mc_rst_n <= 0;
        mc_rst_n <= 0;
    end else begin
        pre_mc_rst_n <= 1;
        mc_rst_n <= pre_mc_rst_n;
    end
end
wire                                trans_fifo_val;
wire    [64-1:0]       trans_fifo_data;
wire                                trans_fifo_rdy;
wire                                fifo_trans_val;
wire    [64-1:0]       fifo_trans_data;
wire                                fifo_trans_rdy;
wire [6     -1:0]     core_axi_awid;
wire [64   -1:0]     core_axi_awaddr;
wire [8    -1:0]     core_axi_awlen;
wire [3   -1:0]     core_axi_awsize;
wire [2  -1:0]     core_axi_awburst;
wire                               core_axi_awlock;
wire [4  -1:0]     core_axi_awcache;
wire [3   -1:0]     core_axi_awprot;
wire [4    -1:0]     core_axi_awqos;
wire [4 -1:0]     core_axi_awregion;
wire [11   -1:0]     core_axi_awuser;
wire                               core_axi_awvalid;
wire                               core_axi_awready;
wire  [6     -1:0]    core_axi_wid;
wire  [512   -1:0]    core_axi_wdata;
wire  [64   -1:0]    core_axi_wstrb;
wire                               core_axi_wlast;
wire  [11   -1:0]    core_axi_wuser;
wire                               core_axi_wvalid;
wire                               core_axi_wready;
wire  [6     -1:0]    core_axi_arid;
wire  [64   -1:0]    core_axi_araddr;
wire  [8    -1:0]    core_axi_arlen;
wire  [3   -1:0]    core_axi_arsize;
wire  [2  -1:0]    core_axi_arburst;
wire                               core_axi_arlock;
wire  [4  -1:0]    core_axi_arcache;
wire  [3   -1:0]    core_axi_arprot;
wire  [4    -1:0]    core_axi_arqos;
wire  [4 -1:0]    core_axi_arregion;
wire  [11   -1:0]    core_axi_aruser;
wire                               core_axi_arvalid;
wire                               core_axi_arready;
wire  [6     -1:0]    core_axi_rid;
wire  [512   -1:0]    core_axi_rdata;
wire  [2   -1:0]    core_axi_rresp;
wire                               core_axi_rlast;
wire  [11   -1:0]    core_axi_ruser;
wire                               core_axi_rvalid;
wire                               core_axi_rready;
wire  [6     -1:0]    core_axi_bid;
wire  [2   -1:0]    core_axi_bresp;
wire  [11   -1:0]    core_axi_buser;
wire                               core_axi_bvalid;
wire                               core_axi_bready;
wire                               init_calib_complete;
wire                               noc_axi4_bridge_rst;
wire                               noc_axi4_bridge_init_done;
noc_bidir_afifo  f1_mig_afifo  (
    .clk_1           (sys_clk      ),
    .rst_1           (~sys_rst_n   ),
    .clk_2           (mc_clk            ),
    .rst_2           (~mc_rst_n         ),
    
    .flit_in_val_1   (mc_flit_in_val    ),
    .flit_in_data_1  (mc_flit_in_data   ),
    .flit_in_rdy_1   (mc_flit_in_rdy    ),
    .flit_out_val_2  (fifo_trans_val    ),
    .flit_out_data_2 (fifo_trans_data   ),
    .flit_out_rdy_2  (fifo_trans_rdy    ),
    
    .flit_in_val_2   (trans_fifo_val    ),
    .flit_in_data_2  (trans_fifo_data   ),
    .flit_in_rdy_2   (trans_fifo_rdy    ),
    .flit_out_val_1  (mc_flit_out_val   ),
    .flit_out_data_1 (mc_flit_out_data  ),
    .flit_out_rdy_1  (mc_flit_out_rdy   )
);
assign m_axi_awid = core_axi_awid;
assign m_axi_awaddr = core_axi_awaddr;
assign m_axi_awlen = core_axi_awlen;
assign m_axi_awsize = core_axi_awsize;
assign m_axi_awburst = core_axi_awburst;
assign m_axi_awlock = core_axi_awlock;
assign m_axi_awcache = core_axi_awcache;
assign m_axi_awprot = core_axi_awprot;
assign m_axi_awqos = core_axi_awqos;
assign m_axi_awregion = core_axi_awregion;
assign m_axi_awuser = core_axi_awuser;
assign m_axi_awvalid = core_axi_awvalid;
assign core_axi_awready = m_axi_awready;
assign m_axi_wid = core_axi_wid;
assign m_axi_wdata = core_axi_wdata;
assign m_axi_wstrb = core_axi_wstrb;
assign m_axi_wlast = core_axi_wlast;
assign m_axi_wuser = core_axi_wuser;
assign m_axi_wvalid = core_axi_wvalid;
assign core_axi_wready = m_axi_wready;
assign m_axi_arid = core_axi_arid;
assign m_axi_araddr = core_axi_araddr;
assign m_axi_arlen = core_axi_arlen;
assign m_axi_arsize = core_axi_arsize;
assign m_axi_arburst = core_axi_arburst;
assign m_axi_arlock = core_axi_arlock;
assign m_axi_arcache = core_axi_arcache;
assign m_axi_arprot = core_axi_arprot;
assign m_axi_arqos = core_axi_arqos;
assign m_axi_arregion = core_axi_arregion;
assign m_axi_aruser = core_axi_aruser;
assign m_axi_arvalid = core_axi_arvalid;
assign core_axi_arready = m_axi_arready;
assign core_axi_rid = m_axi_rid;
assign core_axi_rdata = m_axi_rdata;
assign core_axi_rresp = m_axi_rresp;
assign core_axi_rlast = m_axi_rlast;
assign core_axi_ruser = m_axi_ruser;
assign core_axi_rvalid = m_axi_rvalid;
assign m_axi_rready = core_axi_rready;
assign core_axi_bid = m_axi_bid;
assign core_axi_bresp = m_axi_bresp;
assign core_axi_buser = m_axi_buser;
assign core_axi_bvalid = m_axi_bvalid;
assign m_axi_bready = core_axi_bready;
assign noc_axi4_bridge_rst       = ~mc_rst_n;
assign noc_axi4_bridge_init_done = init_calib_complete;
assign init_calib_complete_out  = init_calib_complete;
noc_axi4_bridge noc_axi4_bridge  (
    .clk                (mc_clk                    ),  
    .rst_n              (~noc_axi4_bridge_rst      ), 
    .uart_boot_en       (uart_boot_en              ),
    .phy_init_done      (noc_axi4_bridge_init_done ),
    .src_bridge_vr_noc2_val(fifo_trans_val),
    .src_bridge_vr_noc2_dat(fifo_trans_data),
    .src_bridge_vr_noc2_rdy(fifo_trans_rdy),
    .bridge_dst_vr_noc3_val(trans_fifo_val),
    .bridge_dst_vr_noc3_dat(trans_fifo_data),
    .bridge_dst_vr_noc3_rdy(trans_fifo_rdy),
    .m_axi_awid(core_axi_awid),
    .m_axi_awaddr(core_axi_awaddr),
    .m_axi_awlen(core_axi_awlen),
    .m_axi_awsize(core_axi_awsize),
    .m_axi_awburst(core_axi_awburst),
    .m_axi_awlock(core_axi_awlock),
    .m_axi_awcache(core_axi_awcache),
    .m_axi_awprot(core_axi_awprot),
    .m_axi_awqos(core_axi_awqos),
    .m_axi_awregion(core_axi_awregion),
    .m_axi_awuser(core_axi_awuser),
    .m_axi_awvalid(core_axi_awvalid),
    .m_axi_awready(core_axi_awready),
    .m_axi_wid(core_axi_wid),
    .m_axi_wdata(core_axi_wdata),
    .m_axi_wstrb(core_axi_wstrb),
    .m_axi_wlast(core_axi_wlast),
    .m_axi_wuser(core_axi_wuser),
    .m_axi_wvalid(core_axi_wvalid),
    .m_axi_wready(core_axi_wready),
    .m_axi_bid(core_axi_bid),
    .m_axi_bresp(core_axi_bresp),
    .m_axi_buser(core_axi_buser),
    .m_axi_bvalid(core_axi_bvalid),
    .m_axi_bready(core_axi_bready),
    .m_axi_arid(core_axi_arid),
    .m_axi_araddr(core_axi_araddr),
    .m_axi_arlen(core_axi_arlen),
    .m_axi_arsize(core_axi_arsize),
    .m_axi_arburst(core_axi_arburst),
    .m_axi_arlock(core_axi_arlock),
    .m_axi_arcache(core_axi_arcache),
    .m_axi_arprot(core_axi_arprot),
    .m_axi_arqos(core_axi_arqos),
    .m_axi_arregion(core_axi_arregion),
    .m_axi_aruser(core_axi_aruser),
    .m_axi_arvalid(core_axi_arvalid),
    .m_axi_arready(core_axi_arready),
    .m_axi_rid(core_axi_rid),
    .m_axi_rdata(core_axi_rdata),
    .m_axi_rresp(core_axi_rresp),
    .m_axi_rlast(core_axi_rlast),
    .m_axi_ruser(core_axi_ruser),
    .m_axi_rvalid(core_axi_rvalid),
    .m_axi_rready(core_axi_rready)
);
 
assign init_calib_complete = ddr_ready;
assign mc_ui_clk_sync_rst = ~mc_rst_n;
 
endmodule 
    
    
    
     
    
    
    
    
    
    
    
    
    
    
    
    
 
module noc_axi4_bridge (
    
    input  wire                                   clk,
    input  wire                                   rst_n,
    input  wire                                   uart_boot_en,
    input  wire                                   phy_init_done, 
    
    input  wire                                   src_bridge_vr_noc2_val,
    input  wire [64-1:0]             src_bridge_vr_noc2_dat,
    output wire                                   src_bridge_vr_noc2_rdy,
    output wire                                   bridge_dst_vr_noc3_val,
    output wire [64-1:0]             bridge_dst_vr_noc3_dat,
    input  wire                                   bridge_dst_vr_noc3_rdy,
    
    output wire [6     -1:0]    m_axi_awid,
    output wire [64   -1:0]    m_axi_awaddr,
    output wire [8    -1:0]    m_axi_awlen,
    output wire [3   -1:0]    m_axi_awsize,
    output wire [2  -1:0]    m_axi_awburst,
    output wire                              m_axi_awlock,
    output wire [4  -1:0]    m_axi_awcache,
    output wire [3   -1:0]    m_axi_awprot,
    output wire [4    -1:0]    m_axi_awqos,
    output wire [4 -1:0]    m_axi_awregion,
    output wire [11   -1:0]    m_axi_awuser,
    output wire                              m_axi_awvalid,
    input  wire                              m_axi_awready,
    output wire  [6     -1:0]    m_axi_wid,
    output wire  [512   -1:0]    m_axi_wdata,
    output wire  [64   -1:0]    m_axi_wstrb,
    output wire                               m_axi_wlast,
    output wire  [11   -1:0]    m_axi_wuser,
    output wire                               m_axi_wvalid,
    input  wire                               m_axi_wready,
    output wire  [6     -1:0]    m_axi_arid,
    output wire  [64   -1:0]    m_axi_araddr,
    output wire  [8    -1:0]    m_axi_arlen,
    output wire  [3   -1:0]    m_axi_arsize,
    output wire  [2  -1:0]    m_axi_arburst,
    output wire                               m_axi_arlock,
    output wire  [4  -1:0]    m_axi_arcache,
    output wire  [3   -1:0]    m_axi_arprot,
    output wire  [4    -1:0]    m_axi_arqos,
    output wire  [4 -1:0]    m_axi_arregion,
    output wire  [11   -1:0]    m_axi_aruser,
    output wire                               m_axi_arvalid,
    input  wire                               m_axi_arready,
    input  wire  [6     -1:0]    m_axi_rid,
    input  wire  [512   -1:0]    m_axi_rdata,
    input  wire  [2   -1:0]    m_axi_rresp,
    input  wire                               m_axi_rlast,
    input  wire  [11   -1:0]    m_axi_ruser,
    input  wire                               m_axi_rvalid,
    output wire                               m_axi_rready,
    input  wire  [6     -1:0]    m_axi_bid,
    input  wire  [2   -1:0]    m_axi_bresp,
    input  wire  [11   -1:0]    m_axi_buser,
    input  wire                               m_axi_bvalid,
    output wire                               m_axi_bready
);
wire [192-1:0] deser_header;
wire [512-1:0] deser_data;
wire deser_val;
wire deser_rdy;
wire [192-1:0] read_req_header;
wire [1-1:0] read_req_id;
wire read_req_val;
wire read_req_rdy;
wire [512-1:0] read_resp_data;
wire [1-1:0] read_resp_id;
wire read_resp_val;
wire read_resp_rdy;
wire write_req_val;
wire [192-1:0] write_req_header;
wire [1-1:0] write_req_id;
wire [512-1:0] write_req_data;
wire write_req_rdy;
wire [1-1:0] write_resp_id;
wire write_resp_val;
wire write_resp_rdy;
wire [192-1:0] ser_header;
wire [512-1:0] ser_data;
wire ser_val;
wire ser_rdy;
noc_axi4_bridge_buffer noc_axi4_bridge_buffer(
    .clk(clk),
    .rst_n(rst_n), 
    .deser_header(deser_header),
    .deser_data(deser_data),
    .deser_val(deser_val),
    .deser_rdy(deser_rdy),
    .read_req_header(read_req_header),
    .read_req_id(read_req_id),
    .read_req_val(read_req_val),
    .read_req_rdy(read_req_rdy),
    .read_resp_data(read_resp_data),
    .read_resp_id(read_resp_id),
    .read_resp_val(read_resp_val),
    .read_resp_rdy(read_resp_rdy),
    .write_req_header(write_req_header),
    .write_req_id(write_req_id),
    .write_req_data(write_req_data),
    .write_req_val(write_req_val), 
    .write_req_rdy(write_req_rdy),
    .write_resp_id(write_resp_id), 
    .write_resp_val(write_resp_val), 
    .write_resp_rdy(write_resp_rdy), 
    .ser_header(ser_header), 
    .ser_data(ser_data), 
    .ser_val(ser_val), 
    .ser_rdy(ser_rdy)
);
noc_axi4_bridge_deser noc_axi4_bridge_deser(
    .clk(clk), 
    .rst_n(rst_n), 
    .flit_in(src_bridge_vr_noc2_dat), 
    .flit_in_val(src_bridge_vr_noc2_val), 
    .flit_in_rdy(src_bridge_vr_noc2_rdy), 
    .phy_init_done(phy_init_done),
    .header_out(deser_header), 
    .data_out(deser_data), 
    .out_val(deser_val), 
    .out_rdy(deser_rdy)
);
noc_axi4_bridge_read noc_axi4_bridge_read (
    .clk(clk), 
    .rst_n(rst_n), 
    .uart_boot_en(uart_boot_en), 
    
    .req_val(read_req_val),
    .req_header(read_req_header),
    .req_id(read_req_id),
    .req_rdy(read_req_rdy),
    .resp_val(read_resp_val),
    .resp_id(read_resp_id),
    .resp_data(read_resp_data),
    .resp_rdy(read_resp_rdy),
    
    .m_axi_arid(m_axi_arid),
    .m_axi_araddr(m_axi_araddr),
    .m_axi_arlen(m_axi_arlen),
    .m_axi_arsize(m_axi_arsize),
    .m_axi_arburst(m_axi_arburst),
    .m_axi_arlock(m_axi_arlock),
    .m_axi_arcache(m_axi_arcache),
    .m_axi_arprot(m_axi_arprot), 
    .m_axi_arqos(m_axi_arqos),
    .m_axi_arregion(m_axi_arregion),
    .m_axi_aruser(m_axi_aruser),
    .m_axi_arvalid(m_axi_arvalid),
    .m_axi_arready(m_axi_arready),
    .m_axi_rid(m_axi_rid),
    .m_axi_rdata(m_axi_rdata),
    .m_axi_rresp(m_axi_rresp),
    .m_axi_rlast(m_axi_rlast), 
    .m_axi_ruser(m_axi_ruser),
    .m_axi_rvalid(m_axi_rvalid),
    .m_axi_rready(m_axi_rready)
);
noc_axi4_bridge_write noc_axi4_bridge_write (
    
    .clk(clk),
    .rst_n(rst_n),
    .uart_boot_en(uart_boot_en), 
    
    .req_val(write_req_val),
    .req_header(write_req_header),
    .req_id(write_req_id),
    .req_data(write_req_data),
    .req_rdy(write_req_rdy),
    .resp_val(write_resp_val),
    .resp_id(write_resp_id),
    .resp_rdy(write_resp_rdy),
    
    .m_axi_awid(m_axi_awid),
    .m_axi_awaddr(m_axi_awaddr),
    .m_axi_awlen(m_axi_awlen),
    .m_axi_awsize(m_axi_awsize),
    .m_axi_awburst(m_axi_awburst),
    .m_axi_awlock(m_axi_awlock),
    .m_axi_awcache(m_axi_awcache),
    .m_axi_awprot(m_axi_awprot),
    .m_axi_awqos(m_axi_awqos),
    .m_axi_awregion(m_axi_awregion),
    .m_axi_awuser(m_axi_awuser),
    .m_axi_awvalid(m_axi_awvalid),
    .m_axi_awready(m_axi_awready),
    .m_axi_wid(m_axi_wid),
    .m_axi_wdata(m_axi_wdata),
    .m_axi_wstrb(m_axi_wstrb),
    .m_axi_wlast(m_axi_wlast),
    .m_axi_wuser(m_axi_wuser),
    .m_axi_wvalid(m_axi_wvalid),
    .m_axi_wready(m_axi_wready),
    .m_axi_bid(m_axi_bid),
    .m_axi_bresp(m_axi_bresp),
    .m_axi_buser(m_axi_buser),
    .m_axi_bvalid(m_axi_bvalid),
    .m_axi_bready(m_axi_bready)
);
noc_axi4_bridge_ser noc_axi4_bridge_ser(
    .clk(clk), 
    .rst_n(rst_n), 
    .header_in(ser_header), 
    .data_in(ser_data), 
    .in_val(ser_val), 
    .in_rdy(ser_rdy), 
    .flit_out(bridge_dst_vr_noc3_dat), 
    .flit_out_val(bridge_dst_vr_noc3_val), 
    .flit_out_rdy(bridge_dst_vr_noc3_rdy)
);
endmodule
    
    
    
     
    
    
    
    
    
    
    
    
    
    
    
    
 
module noc_axi4_bridge_buffer (
  input clk, 
  input rst_n, 
  
  input [192-1:0] deser_header, 
  input [512-1:0] deser_data, 
  input deser_val, 
  output  deser_rdy,
  
  output [192-1:0] read_req_header, 
  output [1-1:0] read_req_id,
  output read_req_val, 
  input  read_req_rdy,
  
  input [512-1:0] read_resp_data, 
  input [1-1:0] read_resp_id,
  input read_resp_val, 
  output  read_resp_rdy,
  
  output [192-1:0] write_req_header, 
  output [1-1:0] write_req_id,
  output [512-1:0] write_req_data, 
  output write_req_val, 
  input  write_req_rdy,
  
  input [1-1:0] write_resp_id,
  input write_resp_val, 
  output  write_resp_rdy,
  
  output [192-1:0] ser_header, 
  output [512-1:0] ser_data, 
  output ser_val, 
  input  ser_rdy
);
localparam INVALID = 1'd0;
localparam WAITING = 1'd1;
localparam READ  = 1'd0;
localparam WRITE = 1'd1;
reg [2-1:0]                          pkt_state_buf ;
reg [192-1:0]   pkt_header[2-1:0];
reg [2-1:0]                          pkt_command;
reg [1-1:0]    fifo_in;
reg [1-1:0]    fifo_out;
reg preser_arb;
reg [2-1:0] bram_rdy;
reg [512-1:0] ser_data_f;
wire [192-1:0] ser_header_f;
reg ser_val_f;
reg [512-1:0] ser_data_ff;
reg [192-1:0] ser_header_ff;
reg ser_val_ff;
wire deser_go = (deser_rdy & deser_val);
wire read_req_go = (read_req_val & read_req_rdy);
wire read_resp_go = (read_resp_val & read_resp_rdy);
wire write_req_go = (write_req_val & write_req_rdy);
wire write_resp_go = (write_resp_val & write_resp_rdy);
wire req_go = read_req_go || write_req_go;
wire preser_rdy = ~ser_val_ff || ser_rdy;
wire ser_go = ser_val & ser_rdy;
always @(posedge clk) begin
    if(~rst_n) begin
        fifo_in <= {1{1'b0}};
        fifo_out <= {1{1'b0}};
    end 
    else begin
        fifo_in <= deser_go ? fifo_in + 1 : fifo_in;
        fifo_out <= req_go ? fifo_out + 1 : fifo_out;
    end
end
genvar i;
generate 
    for (i = 0; i < 2; i = i + 1) begin
        always @(posedge clk) begin
            if(~rst_n) begin
                pkt_state_buf[i] <= INVALID;
                pkt_header[i] <= 192'b0;
                pkt_command[i] <= 1'b0;
            end 
            else begin
                if ((i == fifo_in) & deser_go) begin
                    pkt_state_buf[i] <= WAITING;
                    pkt_header[i] <= deser_header;
                    pkt_command[i] <= (deser_header[21:14] == 8'd20) 
                                   || (deser_header[21:14] == 8'd15);
                end
                else if ((i == fifo_out) & req_go) begin
                      pkt_state_buf[i] <= INVALID;
                      pkt_header[i] <= 192'b0;
                      pkt_command[i] <= 1'b0;
                end
                else begin
                    pkt_state_buf[i] <= pkt_state_buf[i];
                    pkt_header[i] <= pkt_header[i];
                    pkt_command[i] <= pkt_command[i];
                end
            end
        end
    end
endgenerate
noc_axi4_bridge_sram_data noc_axi4_bridge_sram_data
(
    .MEMCLK(clk), 
    .RESET_N(rst_n),
    .CEA(1),
    .AA(write_req_id),
    .RDWENA(1'b1),
    .CEB(deser_go),
    .AB(fifo_in),
    .RDWENB(1'b0),
    .DOUTA(write_req_data),
    .BWB({512{1'b1}}),
    .DINB(deser_data)
);
assign read_req_val = (pkt_state_buf[fifo_out] == WAITING) && (pkt_command[fifo_out] == READ) && bram_rdy[fifo_out];
assign read_req_header = pkt_header[fifo_out];
assign read_req_id = fifo_out;
assign write_req_val = (pkt_state_buf[fifo_out] == WAITING) && (pkt_command[fifo_out] == WRITE) && bram_rdy[fifo_out];
assign write_req_header = pkt_header[fifo_out];
assign write_req_id = fifo_out;
assign deser_rdy = (pkt_state_buf[fifo_in] == INVALID);
always @(posedge clk) begin
    if(~rst_n) begin
        preser_arb <= 1'b0;
    end 
    else begin
        preser_arb <= preser_arb + 1'b1;
    end
end
noc_axi4_bridge_sram_req noc_axi4_bridge_sram_req
(
    .MEMCLK(clk), 
    .RESET_N(rst_n),
    .CEA(1),
    .AA(preser_arb ? write_resp_id : read_resp_id),
    .RDWENA(1'b1),
    .CEB(req_go),
    .AB(fifo_out),
    .RDWENB(1'b0),
    .DOUTA(ser_header_f),
    .BWB({192{1'b1}}),
    .DINB(pkt_header[fifo_out])
);
generate 
    for (i = 0; i < 2; i = i + 1) begin
        always @(posedge clk) begin
            if(~rst_n) begin
                bram_rdy[i] <= 1;
            end 
            else begin
                bram_rdy[i] <= (req_go & (i == fifo_out))               ? 0 
                             : (write_resp_go & (i == write_resp_id)) ? 1
                             : (read_resp_go & (i == read_resp_id))   ? 1
                             :                                          bram_rdy[i];
            end
        end
    end
endgenerate
assign read_resp_rdy = ~preser_arb & preser_rdy;
assign write_resp_rdy = preser_arb & preser_rdy;
always @(posedge clk) begin
    if(~rst_n) begin
        ser_data_f <= 0;
        ser_val_f <= 0;
        ser_header_ff <= 0;
        ser_val_ff <= 0;
        ser_data_ff <= 0;
    end 
    else begin
        if (preser_rdy) begin
            if (preser_arb) begin
                ser_val_f <= write_resp_val;
                ser_data_f <= 0;
            end
            else begin
                ser_val_f <= read_resp_val;
                ser_data_f <= read_resp_data;
            end
            ser_val_ff <= ser_val_f;
            ser_data_ff <= ser_data_f;
            ser_header_ff <= ser_header_f;
        end
        else begin
            ser_val_f <= ser_val_f;
            ser_data_f <= ser_data_f;
            ser_val_ff <= ser_val_ff;
            ser_data_ff <= ser_data_ff;
            ser_header_ff <= ser_header_ff;
        end
    end
end
assign ser_data = ser_data_ff;
assign ser_val = ser_val_ff;
assign ser_header = ser_header_ff;
endmodule
    
    
    
     
    
    
    
    
    
    
    
    
    
    
    
    
 
module noc_axi4_bridge_ser(
  input clk, 
  input rst_n, 
  input [192-1:0] header_in, 
  input [512-1:0] data_in, 
  input in_val, 
  output in_rdy, 
  output reg [64-1:0] flit_out, 
  output  flit_out_val, 
  input flit_out_rdy 
);
localparam ACCEPT = 2'd0;
localparam SEND_HEADER = 2'd1;
localparam SEND_DATA = 2'd2;
reg [512-1:0] data_in_f;
wire in_go = in_val & in_rdy;
wire flit_out_go = flit_out_val & flit_out_rdy;
always @(posedge clk) begin 
  if(~rst_n) begin
    data_in_f <= {512{1'b0}};
  end 
  else if (in_go) begin
    data_in_f <= data_in;
  end
  else begin
    data_in_f <= data_in_f;
  end
end
reg [1:0] state;
reg [8-1:0] remaining_flits;
assign flit_out_val = (state == SEND_HEADER) || (state == SEND_DATA);
assign in_rdy = (state == ACCEPT);
always @(posedge clk) begin
  if(~rst_n) begin
    state <= ACCEPT;
    remaining_flits <= 8'b0;
  end 
  else begin
    case (state)
      ACCEPT: begin
        state <= in_val ? SEND_HEADER : ACCEPT;
        remaining_flits <= 8'b0;
      end
      SEND_HEADER: begin
        if (flit_out_rdy) begin
          if (resp_header[29:22] == 0) begin
            state <= ACCEPT;
            remaining_flits <= 0;
          end
          else begin
            state <= SEND_DATA;
            remaining_flits <= resp_header[29:22];
          end
        end
        else begin
          state <= state;
          remaining_flits <= remaining_flits;
        end
      end
      SEND_DATA: begin
        if (remaining_flits == 8'b1) begin
          state <= flit_out_rdy ? ACCEPT : SEND_DATA;
          remaining_flits <= 0;
        end
        else begin
          state <= SEND_DATA;
          remaining_flits <= flit_out_rdy ? remaining_flits - 8'b1 : remaining_flits;
        end
      end
      default: begin
        
        state <= ACCEPT;
        remaining_flits <= 8'b0;
      end
    endcase 
  end
end
reg [64-1:0] resp_header;
always @(posedge clk) begin
  if (~rst_n) begin
    resp_header <= 64'b0;
  end
  else begin
    case (state)
      ACCEPT: begin
        if (in_go) begin
          resp_header[63:50  ]     <= header_in[191:178];
          resp_header[49:42       ]     <= header_in[177:170     ];
          resp_header[41:34       ]     <= header_in[169:162     ];
          resp_header[33:30   ]     <= header_in[161:158 ];
          resp_header[13:6      ]     <= header_in[13:6    ];
          resp_header[5:0   ]     <= {6{1'b0}};
          case (header_in[21:14])
            8'd19: begin
              resp_header[21:14    ]     <= 8'd24;
              resp_header[29:22  ]     <= 8; 
            end
            8'd20: begin
              resp_header[21:14    ]     <= 8'd25;
              resp_header[29:22  ]     <= 0;
            end
            8'd14: begin
              resp_header[21:14    ]     <= 8'd26;
              resp_header[29:22  ]     <= 8; 
            end
            8'd15: begin
              resp_header[21:14    ]     <= 8'd27;
              resp_header[29:22  ]     <= 0;
            end
            default: begin
              
              resp_header[21:14    ]     <= 8'b0;
              resp_header[29:22  ]     <= 0;
            end
          endcase 
        end
        else begin
          resp_header <= resp_header;
        end
      end
      SEND_HEADER: begin
        if (flit_out_go) begin
          resp_header <= 64'b0;
        end
        else begin
          resp_header <= resp_header;
        end
      end
      SEND_DATA: begin
        resp_header <= resp_header;
      end
      default: begin
        
        resp_header <= 64'b0;
      end
    endcase 
  end
end
always @(*) begin
  case (state)
    ACCEPT: begin
      flit_out = 64'b0;
    end
    SEND_HEADER: begin
      flit_out = resp_header;
    end
    SEND_DATA: begin
      flit_out = data_in_f >> (64 * (8 - remaining_flits));
    end
    default: begin
      flit_out = 64'b0;
    end
  endcase 
end
endmodule
    
    
    
     
    
    
    
    
    
    
    
    
    
    
    
    
 
module noc_axi4_bridge_deser (
  input clk, 
  input rst_n, 
  input [64-1:0] flit_in, 
  input  flit_in_val, 
  output flit_in_rdy, 
  input phy_init_done,
  output [192-1:0] header_out, 
  output [512-1:0] data_out, 
  output out_val, 
  input  out_rdy
);
localparam ACCEPT_W1   = 3'd0;
localparam ACCEPT_W2   = 3'd1;
localparam ACCEPT_W3   = 3'd2;
localparam ACCEPT_DATA = 3'd3;
localparam SEND        = 3'd4;
reg [64-1:0]           pkt_w1;
reg [64-1:0]           pkt_w2;
reg [64-1:0]           pkt_w3; 
reg [64-1:0]           in_data_buf[8-1:0]; 
reg [8-1:0]         remaining_flits; 
reg [2:0]                           state;
assign flit_in_rdy = (state != SEND) & phy_init_done;
wire flit_in_go = flit_in_val & flit_in_rdy;
assign out_val = (state == SEND);
always @(posedge clk) begin
  if(~rst_n) begin
    state <= ACCEPT_W1;
    remaining_flits <= 0;
    pkt_w1 <= 0;
    pkt_w2 <= 0;
    pkt_w3 <= 0;
  end 
  else begin
    case (state)
      ACCEPT_W1: begin
        if (flit_in_go) begin
          state <= ACCEPT_W2;
          remaining_flits <= flit_in[29:22]-1;
          pkt_w1 <= flit_in;  
        end
        else begin
          state <= state;
          remaining_flits <= remaining_flits;
          pkt_w1 <= pkt_w1;
        end
        pkt_w2 <= pkt_w2;
        pkt_w3 <= pkt_w3;  
      end
      ACCEPT_W2: begin
        if (flit_in_go) begin
          state <= ACCEPT_W3;
          remaining_flits <= remaining_flits - 1;
          pkt_w2 <= flit_in;
        end
        else begin
          state <= state;
          remaining_flits <= remaining_flits;
          pkt_w2 <= pkt_w2;
        end
        pkt_w1 <= pkt_w1;
        pkt_w3 <= pkt_w3;  
      end
      ACCEPT_W3: begin
        if (flit_in_go) begin
          if (remaining_flits == 0) begin
            state <= SEND;
            remaining_flits <= 0;
          end
          else begin
            state <= ACCEPT_DATA;
            remaining_flits <= remaining_flits - 1;
          end
          pkt_w3 <= flit_in;  
        end
        else begin
          state <= state;
          remaining_flits <= remaining_flits;
          pkt_w3 <= pkt_w3;  
        end
        pkt_w1 <= pkt_w1;
        pkt_w2 <= pkt_w2;
      end
      ACCEPT_DATA: begin
        if (flit_in_go) begin
          if (remaining_flits == 0) begin
            state <= SEND;
            remaining_flits <= 0;
          end
          else begin
            state <= ACCEPT_DATA;
            remaining_flits <= remaining_flits - 1;
          end
        end
        else begin
          state <= state;
          remaining_flits <= remaining_flits;
        end
        pkt_w1 <= pkt_w1;
        pkt_w2 <= pkt_w2;
        pkt_w3 <= pkt_w3;  
      end
      SEND: begin
        if (out_rdy) begin
          state <= ACCEPT_W1;
          remaining_flits <= 0;
          pkt_w1 <= 0;
          pkt_w2 <= 0;
          pkt_w3 <= 0;
        end
        else begin
          state <= state;
          remaining_flits <= remaining_flits;
          pkt_w1 <= pkt_w1;
          pkt_w2 <= pkt_w2;
          pkt_w3 <= pkt_w3;  
        end
      end
    endcase 
  end
end
genvar i;
generate
  for (i = 0; i < 8; i = i + 1) begin
    always @(posedge clk) begin
      if(~rst_n) begin
        in_data_buf[i] <= 0;
      end 
      else begin
        in_data_buf[i] <= (i == remaining_flits) & flit_in_val & (state == ACCEPT_DATA) ? flit_in 
                        : (state == SEND) & out_rdy                                     ? 0
                        :                                                                 in_data_buf[i];
      end
    end
  end
endgenerate
assign header_out = {pkt_w3, pkt_w2, pkt_w1};
assign data_out = {in_data_buf[0], in_data_buf[1], in_data_buf[2], in_data_buf[3], in_data_buf[4], in_data_buf[5], in_data_buf[6], in_data_buf[7]};
endmodule
    
    
    
     
    
    
    
    
    
    
    
    
    
    
    
    
 
module noc_axi4_bridge_read (
    
    input  wire                                          clk,
    input  wire                                          rst_n,
    input  wire                                          uart_boot_en, 
    
    input  wire                                          req_val,
    input  wire [192-1:0]                  req_header,
    input  wire [1-1:0]  req_id,
    output wire                                          req_rdy,
    output wire                                          resp_val,
    output wire [1-1:0]  resp_id,
    output  reg [512-1:0]                   resp_data,
    input  wire                                          resp_rdy,
    
    output wire  [6     -1:0]    m_axi_arid,
    output wire  [64   -1:0]    m_axi_araddr,
    output wire  [8    -1:0]    m_axi_arlen,
    output wire  [3   -1:0]    m_axi_arsize,
    output wire  [2  -1:0]    m_axi_arburst,
    output wire                               m_axi_arlock,
    output wire  [4  -1:0]    m_axi_arcache,
    output wire  [3   -1:0]    m_axi_arprot,
    output wire  [4    -1:0]    m_axi_arqos,
    output wire  [4 -1:0]    m_axi_arregion,
    output wire  [11   -1:0]    m_axi_aruser,
    output wire                               m_axi_arvalid,
    input  wire                               m_axi_arready,
    input  wire  [6     -1:0]    m_axi_rid,
    input  wire  [512   -1:0]    m_axi_rdata,
    input  wire  [2   -1:0]    m_axi_rresp,
    input  wire                               m_axi_rlast,
    input  wire  [11   -1:0]    m_axi_ruser,
    input  wire                               m_axi_rvalid,
    output wire                               m_axi_rready
);
localparam IDLE = 2'd0;
localparam GOT_REQ = 2'd1;
localparam GOT_RESP = 2'd2;
localparam SEND_RESP = 2'd3;
wire [64-1:0]addr_paddings = 64'b0;
    assign m_axi_arlen    = 8'b0; 
    assign m_axi_arsize   = 3'b110; 
    assign m_axi_arburst  = 2'b01; 
    assign m_axi_arlock   = 1'b0; 
    assign m_axi_arcache  = 4'b11; 
    assign m_axi_arprot   = 3'b0; 
    assign m_axi_arqos    = 4'b0; 
    assign m_axi_arregion = 4'b0; 
    assign m_axi_aruser   = 11'b0; 
wire m_axi_argo = m_axi_arvalid & m_axi_arready;
wire req_go = req_val & req_rdy;
reg req_state;
reg [192-1:0] req_header_f;
reg [1-1:0] req_id_f;
assign req_rdy = (req_state == IDLE);
assign m_axi_arvalid = (req_state == GOT_REQ);
always  @(posedge clk) begin
    if(~rst_n) begin
        req_header_f <= 0;
        req_id_f <= 0;
        req_state <= IDLE;
    end else begin
        case (req_state)
            IDLE: begin
                req_state <= req_go ? GOT_REQ : req_state;
                req_header_f <= req_go ? req_header : req_header_f;
                req_id_f <= req_go ? req_id : req_id_f;
            end
            GOT_REQ: begin
                req_state <= m_axi_argo ? IDLE : req_state;
                req_header_f <= m_axi_argo ? 0 : req_header_f;
                req_id_f <= m_axi_argo ? 0 : req_id_f;
            end
            default : begin
                
                req_header_f <= 0;
                req_id_f <= 0;
                req_state <= IDLE;
            end
        endcase
    end
end
assign m_axi_arid = {{6-1{1'b0}}, req_id_f};
wire [40-1:0] virt_addr = req_header_f[119:80];
wire [64-1:0] phys_addr;
storage_addr_trans #(
.STORAGE_ADDR_WIDTH(64)
) cpu_mig_waddr_translator (
    .va_byte_addr       (virt_addr  ),
    .storage_addr_out   (phys_addr  )
);
reg [6:0] size[2-1:0];
reg [5:0] offset[2-1:0];
reg [1-1:0] resp_id_f;
wire resp_go;
wire uncacheable = (virt_addr[40-1]) 
                || (req_header_f[21:14] == 8'd14);
generate begin
    genvar i;
    for (i = 0; i < 2; i = i + 1) begin
        always @(posedge clk) begin
            if(~rst_n) begin
                size[i] <= 7'b0;
                offset[i] <= 6'b0;
            end 
            else begin
                if ((i == req_id_f) && m_axi_argo) begin
                    if (uncacheable) begin
                        offset[i] <= virt_addr[5:0];
                        case (req_header_f[74:72])
                            3'b000: begin
                                size[i] <= 7'd0;
                            end
                            3'b001: begin
                                size[i] <= 7'd1;
                            end
                            3'b010: begin
                                size[i] <= 7'd2;
                            end
                            3'b011: begin
                                size[i] <= 7'd4;
                            end
                            3'b100: begin
                                size[i] <= 7'd8;
                            end
                            3'b101: begin
                                size[i] <= 7'd16;
                            end
                            3'b110: begin
                                size[i] <= 7'd32;
                            end
                            3'b111: begin
                                size[i] <= 7'd64;
                            end
                            default: begin
                                
                                size[i] <= 7'b0;
                            end
                        endcase
                    end
                    else begin
                        offset[i] <= 6'b0;
                        size[i] <= 7'd64;
                    end
                end
                else if ((i == resp_id_f) & resp_go) begin
                    size[i] <= 7'b0;
                    offset[i] <= 7'b0;
                end
                else begin
                    size[i] <= size[i];
                    offset[i] <= offset[i];
                end
            end
        end
    end
end
endgenerate
wire [64-1:0] addr = uart_boot_en ? {phys_addr[64-4:0], 3'b0} : virt_addr;
assign m_axi_araddr = {addr[64-1:6], 6'b0};
wire m_axi_rgo = m_axi_rvalid & m_axi_rready;
assign resp_go = resp_val & resp_rdy;
reg [1:0] resp_state;
assign resp_val = (resp_state == SEND_RESP);
assign m_axi_rready = (resp_state == IDLE);
always  @(posedge clk) begin
    if(~rst_n) begin
        resp_id_f <= 0;
        resp_state <= IDLE;
    end else begin
        case (resp_state)
            IDLE: begin
                resp_state <= m_axi_rgo ? GOT_RESP : resp_state;
                resp_id_f <= m_axi_rgo ? m_axi_rid : resp_id_f;
            end
            GOT_RESP: begin
                resp_state <= SEND_RESP;
                resp_id_f <= resp_id_f;
            end
            SEND_RESP: begin
                resp_state <= resp_go ? IDLE : resp_state;
                resp_id_f <= resp_go ? 0 : resp_id_f;
            end
            default : begin
                
                resp_id_f <= 0;
                resp_state <= IDLE;
            end
        endcase
    end
end
assign resp_id = resp_id_f;
reg [512-1:0] data_offseted;
always @(posedge clk) begin
    if(~rst_n) begin
        data_offseted <= 0;
    end 
    else begin
        data_offseted <= m_axi_rgo ? (m_axi_rdata >> (8*offset[m_axi_rid])) : 0;
    end
end
always @(posedge clk) begin
    if (~rst_n) begin
        resp_data <= {512{1'b0}};
    end 
    else begin
        case (resp_state)
            GOT_RESP: begin
                case (size[resp_id_f]) 
                    7'd0: begin 
                        resp_data <= {512{1'b0}};
                    end
                    7'd1: begin
                        resp_data <= {512/8{data_offseted[7:0]}};
                    end
                    7'd2: begin
                        resp_data <= {512/16{data_offseted[15:0]}};
                    end
                    7'd4: begin
                        resp_data <= {512/32{data_offseted[31:0]}};
                    end
                    7'd8: begin
                        resp_data <= {512/64{data_offseted[63:0]}};
                    end
                    7'd16: begin
                        resp_data <= {512/128{data_offseted[127:0]}};
                    end
                    7'd32: begin
                        resp_data <= {512/256{data_offseted[255:0]}};
                    end
                    default: begin
                        resp_data <= {512/512{data_offseted[511:0]}};
                    end
                endcase
            end
            SEND_RESP: begin
                resp_data <= resp_go ? {512{1'b0}} : resp_data;
            end
            default: begin
                resp_data <= {512{1'b0}};
            end
        endcase 
    end 
end
endmodule
    
    
    
     
    
    
    
    
    
    
    
    
    
    
    
    
 
module noc_axi4_bridge_write (
    
    input  wire                                                    clk,
    input  wire                                                    rst_n,
    input  wire                                                    uart_boot_en, 
    
    input  wire                                          req_val,
    input  wire [192-1:0]                  req_header,
    input  wire [1-1:0]  req_id,
    input  wire [512-1:0]                   req_data,
    output wire                                          req_rdy,
    output wire                                          resp_val,
    output wire [1-1:0]  resp_id,
    input  wire                                          resp_rdy,
    
    output wire [6     -1:0]     m_axi_awid,
    output wire [64   -1:0]     m_axi_awaddr,
    output wire [8    -1:0]     m_axi_awlen,
    output wire [3   -1:0]     m_axi_awsize,
    output wire [2  -1:0]     m_axi_awburst,
    output wire                               m_axi_awlock,
    output wire [4  -1:0]     m_axi_awcache,
    output wire [3   -1:0]     m_axi_awprot,
    output wire [4    -1:0]     m_axi_awqos,
    output wire [4 -1:0]     m_axi_awregion,
    output wire [11   -1:0]     m_axi_awuser,
    output wire                               m_axi_awvalid,
    input  wire                               m_axi_awready,
    output wire  [6     -1:0]    m_axi_wid,
    output wire  [512   -1:0]    m_axi_wdata,
    output wire  [64   -1:0]    m_axi_wstrb,
    output wire                               m_axi_wlast,
    output wire  [11   -1:0]    m_axi_wuser,
    output wire                               m_axi_wvalid,
    input  wire                               m_axi_wready,
    input  wire  [6     -1:0]    m_axi_bid,
    input  wire  [2   -1:0]    m_axi_bresp,
    input  wire  [11   -1:0]    m_axi_buser,
    input  wire                               m_axi_bvalid,
    output wire                               m_axi_bready
);
localparam IDLE = 3'd0;
localparam GOT_REQ = 3'd1;
localparam PREP_REQ = 3'd2;
localparam SENT_AW = 3'd3;
localparam SENT_W = 3'd4;
localparam GOT_RESP = 3'd1;
    assign m_axi_awlen    = 8'b0; 
    assign m_axi_awsize   = 3'b110; 
    assign m_axi_awburst  = 2'b01; 
    assign m_axi_awlock   = 1'b0; 
    assign m_axi_awcache  = 4'b11; 
    assign m_axi_awprot   = 3'b0; 
    assign m_axi_awqos    = 4'b0; 
    assign m_axi_awregion = 4'b0; 
    assign m_axi_awuser   = 11'b0; 
    assign m_axi_wuser    = 11'b0; 
wire [64-1:0] addr_paddings = 64'b0;
wire m_axi_awgo = m_axi_awvalid & m_axi_awready;
wire m_axi_wgo = m_axi_wvalid & m_axi_wready;
wire req_go = req_val & req_rdy;
assign m_axi_wlast = m_axi_wvalid;
reg [2:0] req_state;
reg [192-1:0] req_header_f;
reg [1-1:0] req_id_f;
reg [512-1:0] req_data_f;
assign req_rdy = (req_state == IDLE);
assign m_axi_awvalid = (req_state == PREP_REQ) || (req_state == SENT_W);
assign m_axi_wvalid = (req_state == PREP_REQ) || (req_state == SENT_AW);
always  @(posedge clk) begin
    if(~rst_n) begin
        req_header_f <= 0;
        req_id_f <= 0;
        req_state <= IDLE;
        req_data_f <= 0;
    end else begin
        case (req_state)
            IDLE: begin
                req_state <= req_go ? GOT_REQ : req_state;
                req_header_f <= req_go ? req_header : req_header_f;
                req_id_f <= req_go ? req_id : req_id_f;
                req_data_f <= req_data_f;
            end
            GOT_REQ: begin
                req_state <= PREP_REQ;
                req_header_f <= req_header_f;
                req_id_f <= req_id_f;
                req_data_f <= req_data; 
            end
            PREP_REQ: begin
                req_state <= (m_axi_awgo & m_axi_wgo) ? IDLE : m_axi_awgo ? SENT_AW : m_axi_wgo ? SENT_W : req_state;
                req_header_f <= (m_axi_awgo & m_axi_wgo) ? 0 : req_header_f;
                req_id_f <= (m_axi_awgo & m_axi_wgo) ? 0 : req_id_f;
                req_data_f <= (m_axi_awgo & m_axi_wgo) ? 0 : req_data_f;
            end
            SENT_AW: begin
                req_state <= m_axi_wgo ? IDLE : req_state;
                req_header_f <= m_axi_wgo ? 0 : req_header_f;
                req_id_f <= m_axi_wgo ? 0 : req_id_f;
                req_data_f <= m_axi_wgo ? 0 : req_data_f;
            end
            SENT_W: begin
                req_state <= m_axi_awgo ? IDLE : req_state;
                req_header_f <= m_axi_awgo ? 0 : req_header_f;
                req_id_f <= m_axi_awgo ? 0 : req_id_f;
                req_data_f <= m_axi_awgo ? 0 : req_data_f;
            end
            default : begin
                req_header_f <= 0;
                req_id_f <= 0;
                req_state <= IDLE;
                req_data_f <= 0;
            end
        endcase
    end
end
assign m_axi_awid = {{6-1{1'b0}}, req_id_f};
assign m_axi_wid = {{6-1{1'b0}}, req_id_f};
wire [40-1:0] virt_addr = req_header_f[119:80];
wire [64-1:0] phys_addr;
wire uncacheable = (virt_addr[40-1])
                || (req_header_f[21:14] == 8'd15);
storage_addr_trans #(
.STORAGE_ADDR_WIDTH(64)
) cpu_mig_raddr_translator (
    .va_byte_addr       (virt_addr  ),
    .storage_addr_out   (phys_addr  )
);
reg [64-1:0] strb_before_offset;
reg [5:0] offset;
reg [64-1:0] addr;
always @(posedge clk) begin
    if (~rst_n) begin
        offset <= 6'b0;
        strb_before_offset <= 64'b0;
        addr <= 64'b0;
    end
    else begin
        if (uncacheable) begin
            case (req_header_f[74:72])
                3'b000: begin
                    strb_before_offset <= 64'b0;
                end
                3'b001: begin
                    strb_before_offset <= 64'b1;
                end
                3'b010: begin
                    strb_before_offset <= 64'b11;
                end
                3'b011: begin
                    strb_before_offset <= 64'hf;
                end
                3'b100: begin
                    strb_before_offset <= 64'hff;
                end
                3'b101: begin
                    strb_before_offset <= 64'hffff;
                end
                3'b110: begin
                    strb_before_offset <= 64'hffffffff;
                end
                3'b111: begin
                    strb_before_offset <= 64'hffffffffffffffff;
                end
                default: begin
                    
                    strb_before_offset <= 64'b0;
                end
            endcase
        end
        else begin
            strb_before_offset <= 64'hffffffffffffffff;
        end
        offset <= uncacheable ? virt_addr[5:0] : 6'b0;
        addr <= uart_boot_en ? {phys_addr[64-4:0], 3'b0} : virt_addr;
    end
end
assign m_axi_awaddr = {addr[64-1:6], 6'b0};
assign m_axi_wstrb = strb_before_offset << offset;
assign m_axi_wdata = req_data_f << (8*offset);
wire m_axi_bgo = m_axi_bvalid & m_axi_bready;
wire resp_go = resp_val & resp_rdy;
reg [2:0] resp_state;
reg [1-1:0]resp_id_f;
assign resp_val = (resp_state == GOT_RESP);
assign m_axi_bready = (resp_state == IDLE);
always  @(posedge clk) begin
    if(~rst_n) begin
        resp_id_f <= 0;
        resp_state <= IDLE;
    end else begin
        case (resp_state)
            IDLE: begin
                resp_state <= m_axi_bgo ? GOT_RESP : resp_state;
                resp_id_f <= m_axi_bgo ? m_axi_bid : resp_id_f;
            end
            GOT_RESP: begin
                resp_state <= resp_go ? IDLE : resp_state;
                resp_id_f <= resp_go ? 0 : resp_id_f;
            end
            default : begin
                resp_state <= IDLE;
                resp_id_f <= 0;
            end
        endcase
    end
end
assign resp_id = resp_id_f;
endmodule
    
    
    
     
    
    
    
    
    
    
    
    
    
    
    
    
 
module axi4_zeroer (
    input   clk,
    input   rst_n,
    input   init_calib_complete_in,
    output  init_calib_complete_out,
    
    input wire  [6     -1:0]     s_axi_awid,
    input wire  [64   -1:0]     s_axi_awaddr,
    input wire  [8    -1:0]     s_axi_awlen,
    input wire  [3   -1:0]     s_axi_awsize,
    input wire  [2  -1:0]     s_axi_awburst,
    input wire                                s_axi_awlock,
    input wire  [4  -1:0]     s_axi_awcache,
    input wire  [3   -1:0]     s_axi_awprot,
    input wire  [4    -1:0]     s_axi_awqos,
    input wire  [4 -1:0]     s_axi_awregion,
    input wire  [11   -1:0]     s_axi_awuser,
    input wire                                s_axi_awvalid,
    output reg                                s_axi_awready,
    input wire   [6     -1:0]    s_axi_wid,
    input wire   [512   -1:0]    s_axi_wdata,
    input wire   [64   -1:0]    s_axi_wstrb,
    input wire                                s_axi_wlast,
    input wire   [11   -1:0]    s_axi_wuser,
    input wire                                s_axi_wvalid,
    output reg                                s_axi_wready,
    input wire   [6     -1:0]    s_axi_arid,
    input wire   [64   -1:0]    s_axi_araddr,
    input wire   [8    -1:0]    s_axi_arlen,
    input wire   [3   -1:0]    s_axi_arsize,
    input wire   [2  -1:0]    s_axi_arburst,
    input wire                                s_axi_arlock,
    input wire   [4  -1:0]    s_axi_arcache,
    input wire   [3   -1:0]    s_axi_arprot,
    input wire   [4    -1:0]    s_axi_arqos,
    input wire   [4 -1:0]    s_axi_arregion,
    input wire   [11   -1:0]    s_axi_aruser,
    input wire                                s_axi_arvalid,
    output reg                                s_axi_arready,
    output reg  [6     -1:0]     s_axi_rid,
    output reg  [512   -1:0]     s_axi_rdata,
    output reg  [2   -1:0]     s_axi_rresp,
    output reg                                s_axi_rlast,
    output reg  [11   -1:0]     s_axi_ruser,
    output reg                                s_axi_rvalid,
    input wire                                s_axi_rready,
    output reg  [6     -1:0]     s_axi_bid,
    output reg  [2   -1:0]     s_axi_bresp,
    output reg  [11   -1:0]     s_axi_buser,
    output reg                                s_axi_bvalid,
    input wire                                s_axi_bready,    
    
    output reg  [6     -1:0]     m_axi_awid,
    output reg  [64   -1:0]     m_axi_awaddr,
    output reg  [8    -1:0]     m_axi_awlen,
    output reg  [3   -1:0]     m_axi_awsize,
    output reg  [2  -1:0]     m_axi_awburst,
    output reg                                m_axi_awlock,
    output reg  [4  -1:0]     m_axi_awcache,
    output reg  [3   -1:0]     m_axi_awprot,
    output reg  [4    -1:0]     m_axi_awqos,
    output reg  [4 -1:0]     m_axi_awregion,
    output reg  [11   -1:0]     m_axi_awuser,
    output reg                                m_axi_awvalid,
    input  wire                               m_axi_awready,
    output reg   [6     -1:0]    m_axi_wid,
    output reg   [512   -1:0]    m_axi_wdata,
    output reg   [64   -1:0]    m_axi_wstrb,
    output reg                                m_axi_wlast,
    output reg   [11   -1:0]    m_axi_wuser,
    output reg                                m_axi_wvalid,
    input  wire                               m_axi_wready,
    output reg   [6     -1:0]    m_axi_arid,
    output reg   [64   -1:0]    m_axi_araddr,
    output reg   [8    -1:0]    m_axi_arlen,
    output reg   [3   -1:0]    m_axi_arsize,
    output reg   [2  -1:0]    m_axi_arburst,
    output reg                                m_axi_arlock,
    output reg   [4  -1:0]    m_axi_arcache,
    output reg   [3   -1:0]    m_axi_arprot,
    output reg   [4    -1:0]    m_axi_arqos,
    output reg   [4 -1:0]    m_axi_arregion,
    output reg   [11   -1:0]    m_axi_aruser,
    output reg                                m_axi_arvalid,
    input  wire                               m_axi_arready,
    input  wire  [6     -1:0]    m_axi_rid,
    input  wire  [512   -1:0]    m_axi_rdata,
    input  wire  [2   -1:0]    m_axi_rresp,
    input  wire                               m_axi_rlast,
    input  wire  [11   -1:0]    m_axi_ruser,
    input  wire                               m_axi_rvalid,
    output reg                                m_axi_rready,
    input  wire  [6     -1:0]    m_axi_bid,
    input  wire  [2   -1:0]    m_axi_bresp,
    input  wire  [11   -1:0]    m_axi_buser,
    input  wire                               m_axi_bvalid,
    output reg                                m_axi_bready
);
localparam reg [63:0] BOARD_MEM_SIZE_MB = 1024;
localparam reg [64-1:0] MAX_MEM_ADDR      = (BOARD_MEM_SIZE_MB * 2**20);
localparam REQUESTS_NEEDED  = MAX_MEM_ADDR / 64; 
localparam MAX_OUTSTANDING = 16;
wire zeroer_req_val;
wire zeroer_resp_rdy;
wire req_go;
wire resp_go;
reg [64-1:0] req_sent;
reg [64-1:0] resp_got;
reg [3:0] outstanding;
wire [64-1:0] zeroer_addr;
wire zeroer_wlast;
assign zeroer_req_val = init_calib_complete_in 
                      & (req_sent < REQUESTS_NEEDED) 
                      & (outstanding != MAX_OUTSTANDING-1) 
                      & m_axi_awready
                      & m_axi_wready
                      & rst_n;
assign zeroer_resp_rdy = init_calib_complete_in 
                       & (resp_got < REQUESTS_NEEDED) 
                       & rst_n;
assign req_go = zeroer_req_val;
assign resp_go = zeroer_resp_rdy & m_axi_bvalid;
always @(posedge clk) begin
    if(~rst_n) begin
        req_sent <= 0;
        resp_got <= 0;
        outstanding <= 0;
    end 
    else begin
        req_sent <= req_sent + req_go;
        resp_got <= resp_got + resp_go;
        outstanding <= req_go & resp_go ? outstanding 
                     : req_go           ? outstanding + 1 
                     : resp_go          ? outstanding - 1 
                     :                    outstanding;
    end
end
assign init_calib_complete_out = (req_sent == REQUESTS_NEEDED) & 
                                 (resp_got == REQUESTS_NEEDED);
assign zeroer_addr = req_sent * 64;
assign zeroer_wlast = zeroer_req_val;
always @(*) begin
    if (~init_calib_complete_out) begin
        m_axi_awid = 6'b0;
        m_axi_awaddr = zeroer_addr;
        m_axi_awlen = 8'b0;
        m_axi_awsize = 3'b110;
        m_axi_awburst = 2'b01;
        m_axi_awlock = 1'b0;
        m_axi_awcache = 4'b11;
        m_axi_awprot = 3'b10;
        m_axi_awqos = 4'b0;
        m_axi_awregion = 4'b0;
        m_axi_awuser = 11'b0;
        m_axi_awvalid = zeroer_req_val;
        m_axi_wid = 6'b0;
        m_axi_wdata = {512{1'b0}};
        m_axi_wstrb = {64{1'b1}};
        m_axi_wlast = zeroer_wlast;
        m_axi_wuser = 11'b0;
        m_axi_wvalid = zeroer_req_val;
        m_axi_arid = 6'b0;
        m_axi_araddr = 64'b0;
        m_axi_arlen = 8'b0;
        m_axi_arsize = 3'b110;
        m_axi_arburst = 2'b01;
        m_axi_arlock = 1'b0;
        m_axi_arcache = 4'b11;
        m_axi_arprot = 3'b10;
        m_axi_arqos = 4'b0;
        m_axi_arregion = 4'b0;
        m_axi_aruser = 11'b0;
        m_axi_arvalid = 1'b0;
        m_axi_rready = 1'b0;
        m_axi_bready = zeroer_resp_rdy;
        s_axi_awready = 1'b0;
        s_axi_wready = 1'b0;
        s_axi_arready = 1'b0;
        s_axi_rid = 6'b0;
        s_axi_rdata = 512'b0;
        s_axi_rresp = 2'b0;
        s_axi_rlast = 1'b0;
        s_axi_ruser = 11'b0;
        s_axi_rvalid = 1'b0;
        s_axi_bid = 6'b0;
        s_axi_bresp = 2'b0;
        s_axi_buser = 11'b0;
        s_axi_bvalid = 1'b0;
    end
    else begin
        m_axi_awid = s_axi_awid;
        m_axi_awaddr = s_axi_awaddr;
        m_axi_awlen = s_axi_awlen;
        m_axi_awsize = s_axi_awsize;
        m_axi_awburst = s_axi_awburst;
        m_axi_awlock = s_axi_awlock;
        m_axi_awcache = s_axi_awcache;
        m_axi_awprot = s_axi_awprot;
        m_axi_awqos = s_axi_awqos;
        m_axi_awregion = s_axi_awregion;
        m_axi_awuser = s_axi_awuser;
        m_axi_awvalid = s_axi_awvalid;
        s_axi_awready = m_axi_awready;
        m_axi_wid = s_axi_wid;
        m_axi_wdata = s_axi_wdata;
        m_axi_wstrb = s_axi_wstrb;
        m_axi_wlast = s_axi_wlast;
        m_axi_wuser = s_axi_wuser;
        m_axi_wvalid = s_axi_wvalid;
        s_axi_wready = m_axi_wready;
        m_axi_arid = s_axi_arid;
        m_axi_araddr = s_axi_araddr;
        m_axi_arlen = s_axi_arlen;
        m_axi_arsize = s_axi_arsize;
        m_axi_arburst = s_axi_arburst;
        m_axi_arlock = s_axi_arlock;
        m_axi_arcache = s_axi_arcache;
        m_axi_arprot = s_axi_arprot;
        m_axi_arqos = s_axi_arqos;
        m_axi_arregion = s_axi_arregion;
        m_axi_aruser = s_axi_aruser;
        m_axi_arvalid = s_axi_arvalid;
        s_axi_arready = m_axi_arready;
        s_axi_rid = m_axi_rid;
        s_axi_rdata = m_axi_rdata;
        s_axi_rresp = m_axi_rresp;
        s_axi_rlast = m_axi_rlast;
        s_axi_ruser = m_axi_ruser;
        s_axi_rvalid = m_axi_rvalid;
        m_axi_rready = s_axi_rready;
        s_axi_bid = m_axi_bid;
        s_axi_bresp = m_axi_bresp;
        s_axi_buser = m_axi_buser;
        s_axi_bvalid = m_axi_bvalid;
        m_axi_bready = s_axi_bready;
    end
end
endmodule
 
module noc_axi4_bridge_sram_data
(
input wire MEMCLK,
input wire RESET_N,
input wire CEA,
input wire [1-1:0] AA,
input wire RDWENA,
input wire CEB,
input wire [1-1:0] AB,
input wire RDWENB,
input wire [512-1:0] BWA,
input wire [512-1:0] DINA,
output wire [512-1:0] DOUTA,
input wire [512-1:0] BWB,
input wire [512-1:0] DINB,
output wire [512-1:0] DOUTB,
input wire [4-1:0] BIST_COMMAND,
input wire [4-1:0] BIST_DIN,
output reg [4-1:0] BIST_DOUT,
input wire [8-1:0] SRAMID
);
  
wire [512-1:0] DOUTA_bram;
wire [512-1:0] DOUTB_bram;
assign DOUTA = DOUTA_bram;
assign DOUTB = DOUTB_bram;
bram_1r1w_wrapper #(
   .NAME          (""             ),
   .DEPTH         (2),
   .ADDR_WIDTH    (1),
   .BITMASK_WIDTH (512),
   .DATA_WIDTH    (512)
)   noc_axi4_bridge_sram_data (
   .MEMCLK        (MEMCLK     ),
   .RESET_N        (RESET_N     ),
   .CEA        (CEA     ),
   .AA        (AA     ),
   .AB        (AB     ),
   .RDWENA        (RDWENA     ),
   .CEB        (CEB     ),
   .RDWENB        (RDWENB     ),
   .BWA        (BWA     ),
   .DINA        (DINA     ),
   .DOUTA        (DOUTA_bram     ),
   .BWB        (BWB     ),
   .DINB        (DINB     ),
   .DOUTB        (DOUTB_bram     )
);
      
  
 
 endmodule
 
module noc_axi4_bridge_sram_req
(
input wire MEMCLK,
input wire RESET_N,
input wire CEA,
input wire [1-1:0] AA,
input wire RDWENA,
input wire CEB,
input wire [1-1:0] AB,
input wire RDWENB,
input wire [192-1:0] BWA,
input wire [192-1:0] DINA,
output wire [192-1:0] DOUTA,
input wire [192-1:0] BWB,
input wire [192-1:0] DINB,
output wire [192-1:0] DOUTB,
input wire [4-1:0] BIST_COMMAND,
input wire [4-1:0] BIST_DIN,
output reg [4-1:0] BIST_DOUT,
input wire [8-1:0] SRAMID
);
  
wire [192-1:0] DOUTA_bram;
wire [192-1:0] DOUTB_bram;
assign DOUTA = DOUTA_bram;
assign DOUTB = DOUTB_bram;
bram_1r1w_wrapper #(
   .NAME          (""             ),
   .DEPTH         (2),
   .ADDR_WIDTH    (1),
   .BITMASK_WIDTH (192),
   .DATA_WIDTH    (192)
)   noc_axi4_bridge_sram_req (
   .MEMCLK        (MEMCLK     ),
   .RESET_N        (RESET_N     ),
   .CEA        (CEA     ),
   .AA        (AA     ),
   .AB        (AB     ),
   .RDWENA        (RDWENA     ),
   .CEB        (CEB     ),
   .RDWENB        (RDWENB     ),
   .BWA        (BWA     ),
   .DINA        (DINA     ),
   .DOUTA        (DOUTA_bram     ),
   .BWB        (BWB     ),
   .DINB        (DINB     ),
   .DOUTB        (DOUTB_bram     )
);
      
  
 
 endmodule
module async_fifo 
#(
	parameter DSIZE = 64,
	parameter ASIZE = 5,
	parameter MEMSIZE = 16 
)
(
	rdata, 
	rempty,
	rclk,
	ren,
	wdata,
	wfull,
	wclk,
	wval,
	wreset,
	rreset
	);
output  [DSIZE-1:0] 	rdata;
output			rempty;
output 			wfull;
input	[DSIZE-1:0]	wdata;
input			wval;
input			ren;
input			rclk;
input			wclk;
input 			wreset;
input			rreset;
reg	[ASIZE-1:0]	g_wptr;
reg	[ASIZE-1:0]	g_rptr;
reg	[ASIZE-1:0]	g_rsync1, g_rsync2;
reg	[ASIZE-1:0]	g_wsync1, g_wsync2;
reg	[DSIZE-1:0] 	fifo[MEMSIZE-1:0];
wire [ASIZE-1:0] b_wptr;
wire [ASIZE-1:0] b_wptr_next;
wire [ASIZE-1:0] g_wptr_next;
wire [ASIZE-1:0] b_rptr;
wire [ASIZE-1:0] b_rptr_next;
wire [ASIZE-1:0] g_rptr_next;
assign b_wptr[ASIZE-1:0] = ({1'b0, b_wptr[ASIZE-1:1]} ^ g_wptr[ASIZE-1:0]);
assign b_rptr[ASIZE-1:0] = ({1'b0, b_rptr[ASIZE-1:1]} ^ g_rptr[ASIZE-1:0]);
assign b_wptr_next = b_wptr + 1;
assign b_rptr_next = b_rptr + 1;
assign g_wptr_next[ASIZE-1:0] = {1'b0, b_wptr_next[ASIZE-1:1]} ^ b_wptr_next[ASIZE-1:0];
assign g_rptr_next[ASIZE-1:0] = {1'b0, b_rptr_next[ASIZE-1:1]} ^ b_rptr_next[ASIZE-1:0];
assign wfull =  (g_wptr[ASIZE-1]   != g_rsync2[ASIZE-1]  ) && 
		(g_wptr[ASIZE-2]   != g_rsync2[ASIZE-2]  ) &&
		(g_wptr[ASIZE-3:0] == g_rsync2[ASIZE-3:0]) ||
		(wreset || rreset);
assign rempty =  (g_wsync2[ASIZE-1:0] == g_rptr[ASIZE-1:0]) ||
	         (wreset || rreset);
assign rdata = fifo[b_rptr[ASIZE-2:0]];
always @(posedge rclk) begin
	if (rreset) begin
		g_rptr <= 0;
	end
	else if (ren && !rempty) begin
		g_rptr <= g_rptr_next;
	end
	g_wsync1 <= g_wptr;
	g_wsync2 <= g_wsync1;
end
always @(posedge wclk) begin
	if (wreset) begin
		g_wptr <= 0;
	end
	else if (wval && !wfull) begin
		fifo[b_wptr[ASIZE-2:0]] <= wdata;
		g_wptr <= g_wptr_next;
	end
	g_rsync1 <= g_rptr;
	g_rsync2 <= g_rsync1;
	
end
endmodule
module bram_1r1w_wrapper 
#(parameter NAME="", DEPTH=1, ADDR_WIDTH=1, BITMASK_WIDTH=1, DATA_WIDTH=1)
(
  input wire MEMCLK,
  input wire RESET_N,
  input wire CEA,
  input wire [ADDR_WIDTH-1:0] AA,
  input wire [ADDR_WIDTH-1:0] AB,
  input wire RDWENA,
  input wire CEB,
  input wire RDWENB,
  input wire [DATA_WIDTH-1:0] BWA,
  input wire [DATA_WIDTH-1:0] DINA,
  output reg [DATA_WIDTH-1:0] DOUTA,
  input wire [DATA_WIDTH-1:0] BWB,
  input wire [DATA_WIDTH-1:0] DINB,
  output wire [DATA_WIDTH-1:0] DOUTB
  
  
  
  
);
wire                            write_enable_in;
wire                            read_enable_in;
reg                             write_enable_in_reg;
reg   [ADDR_WIDTH-1:0    ]      WRITE_ADDRESS_REG;
reg   [ADDR_WIDTH-1:0    ]      WRITE_ADDRESS_REG_muxed;
reg   [BITMASK_WIDTH-1:0 ]      WRITE_BIT_MASK_REG;
reg   [DATA_WIDTH-1:0    ]      DIN_r;
reg                             read_enable_in_reg;
reg   [DATA_WIDTH-1:0    ]      bram_data_in_r;
wire                            bram_write_en;
reg                            bram_write_en_muxed;
wire                            bram_read_en;
wire                            bram_write_read_en;
reg  [DATA_WIDTH-1:0    ]      bram_data_write_read_out_reg;
reg  [DATA_WIDTH-1:0    ]      bram_data_read_out_reg;
reg  [DATA_WIDTH-1:0    ]      bram_data_in;
reg  [DATA_WIDTH-1:0    ]      bram_data_in_muxed;
wire  [DATA_WIDTH-1:0    ]      last_wrote_data;
wire                            rw_conflict;
reg                             rw_conflict_r;
wire                            ww_conflict;
reg                             ww_conflict_r;
assign read_enable_in    = CEA & (RDWENA == 1'b1);
assign write_enable_in   = CEB & (RDWENB == 1'b0);
wire [ADDR_WIDTH-1:0    ] READ_ADDRESS = AA;
wire [ADDR_WIDTH-1:0    ] WRITE_ADDRESS = AB;
wire [BITMASK_WIDTH-1:0    ] WRITE_BIT_MASK = BWB;
always @(posedge MEMCLK) begin
  write_enable_in_reg <= write_enable_in;
  WRITE_ADDRESS_REG   <= WRITE_ADDRESS;
  WRITE_BIT_MASK_REG  <= WRITE_BIT_MASK;
  DIN_r <= DINB;
  read_enable_in_reg  <= read_enable_in;
  bram_data_in_r <= bram_data_in;
  rw_conflict_r  <= rw_conflict;
  ww_conflict_r  <= ww_conflict;
  
end
assign rw_conflict      = write_enable_in_reg & read_enable_in & (WRITE_ADDRESS_REG == READ_ADDRESS);
assign ww_conflict      = write_enable_in_reg & write_enable_in & (WRITE_ADDRESS_REG == WRITE_ADDRESS);
assign DOUTB = {DATA_WIDTH{1'bx}}; 
always @ * begin
  bram_data_in = (DIN_r & WRITE_BIT_MASK_REG);
  if (ww_conflict_r)
    bram_data_in = bram_data_in | (bram_data_in_r & ~WRITE_BIT_MASK_REG);
  else
    bram_data_in = bram_data_in | (bram_data_write_read_out_reg & ~WRITE_BIT_MASK_REG);
  
  
  
  if (read_enable_in_reg) begin
    DOUTA = bram_data_read_out_reg; 
    if (rw_conflict_r) begin
      DOUTA = bram_data_in_r;
    end
  end
end
assign bram_write_en      = write_enable_in_reg;
assign bram_read_en         = (read_enable_in) & ~rw_conflict;             
assign bram_write_read_en         = (write_enable_in) & ~ww_conflict;             
reg [DATA_WIDTH-1:0] ram [DEPTH-1:0];
always @(posedge MEMCLK) begin
  if (bram_write_en_muxed) begin
    ram[WRITE_ADDRESS_REG_muxed] <= bram_data_in_muxed;
  end
  if (bram_read_en) begin
    bram_data_read_out_reg <= ram[READ_ADDRESS];
  end
  if (bram_write_read_en) begin
    bram_data_write_read_out_reg <= ram[WRITE_ADDRESS];
  end
end
localparam INIT_STATE = 1'd0;
localparam DONE_STATE  = 1'd1;
reg [ADDR_WIDTH-1:0] bist_index;
reg [ADDR_WIDTH-1:0] bist_index_next;
reg init_done;
reg init_done_next;
always @ (posedge MEMCLK)
begin
   if (!RESET_N)
   begin
      bist_index <= 0;
      init_done <= 0;
   end
   else
   begin
      bist_index <= bist_index_next;
      init_done <= init_done_next;
   end
end
always @ *
begin
   bist_index_next = init_done ? bist_index : bist_index + 1;
   init_done_next = ((|(~bist_index)) == 0) | init_done;
end
always @ *
begin
   if (!init_done)
   begin
      WRITE_ADDRESS_REG_muxed = bist_index;
      bram_write_en_muxed = 1'b1;
      bram_data_in_muxed = {DATA_WIDTH{1'b0}};
   end
   else
   begin
      WRITE_ADDRESS_REG_muxed = WRITE_ADDRESS_REG;
      bram_write_en_muxed = bram_write_en;
      bram_data_in_muxed = bram_data_in;
   end
end
endmodule
module bram_1rw_wrapper 
#(parameter NAME="", DEPTH=1, ADDR_WIDTH=1, BITMASK_WIDTH=1, DATA_WIDTH=1)
(
    input                         MEMCLK,
    input wire RESET_N,
    input                         CE,
    input   [ADDR_WIDTH-1:0]      A,
    input                         RDWEN,
    input   [BITMASK_WIDTH-1:0]   BW,
    input   [DATA_WIDTH-1:0]      DIN,
    output  [DATA_WIDTH-1:0]      DOUT
);
wire                            write_en;
wire                            read_en;
reg                             wen_r;
reg   [ADDR_WIDTH-1:0    ]      A_r;
reg   [BITMASK_WIDTH-1:0 ]      BW_r;
reg   [DATA_WIDTH-1:0    ]      DIN_r;
reg   [DATA_WIDTH-1:0    ]      DOUT_r;
reg                             ren_r;
reg   [DATA_WIDTH-1:0    ]      bram_data_in_r;
wire                            bram_wen;
wire                            bram_ren;
reg  [DATA_WIDTH-1:0    ]      bram_data_out;
wire  [DATA_WIDTH-1:0    ]      bram_data_in;
wire  [DATA_WIDTH-1:0    ]      up_to_date_data;
wire                            rw_conflict;
reg                             rw_conflict_r;
reg   [ADDR_WIDTH-1:0    ]      WRITE_ADDRESS_REG_muxed;
reg                            bram_write_en_muxed;
reg  [DATA_WIDTH-1:0    ]      bram_data_in_muxed;
assign write_en   = CE & (RDWEN == 1'b0);
assign read_en    = CE & (RDWEN == 1'b1);
always @(posedge MEMCLK) begin
   wen_r <= write_en;
   A_r   <= A;
   BW_r  <= BW;
   DIN_r <= DIN;
end
always @(posedge MEMCLK) begin
  ren_r  <= read_en;
end
always @(posedge MEMCLK)
   bram_data_in_r <= bram_data_in;
always @(posedge MEMCLK)
   rw_conflict_r  <= rw_conflict;
always @(posedge MEMCLK)
  DOUT_r  <= DOUT;
assign bram_data_in = (up_to_date_data & ~BW_r) | (DIN_r & BW_r);
assign rw_conflict      = wen_r & CE & (A_r == A);                         
assign up_to_date_data  = rw_conflict_r ? bram_data_in_r : bram_data_out;  
assign bram_ren         = (read_en | write_en) & ~rw_conflict;             
                                                                        
assign bram_wen      = wen_r;
assign DOUT          = ren_r ? up_to_date_data : DOUT_r;
reg [DATA_WIDTH-1:0] ram [DEPTH-1:0];
always @(posedge MEMCLK) begin
  if (bram_write_en_muxed) begin
      ram[WRITE_ADDRESS_REG_muxed] <= bram_data_in_muxed;
  end
  if (bram_ren) begin
    bram_data_out <= ram[A];
  end
end
 
localparam INIT_STATE = 1'd0;
localparam DONE_STATE  = 1'd1;
reg [ADDR_WIDTH-1:0] bist_index;
reg [ADDR_WIDTH-1:0] bist_index_next;
reg init_done;
reg init_done_next;
always @ (posedge MEMCLK)
begin
   if (!RESET_N)
   begin
      bist_index <= 0;
      init_done <= 0;
   end
   else
   begin
      bist_index <= bist_index_next;
      init_done <= init_done_next;
   end
end
always @ *
begin
   bist_index_next = init_done ? bist_index : bist_index + 1;
   init_done_next = ((|(~bist_index)) == 0) | init_done;
end
always @ *
begin
   if (!init_done)
   begin
      WRITE_ADDRESS_REG_muxed = bist_index;
      bram_write_en_muxed = 1'b1;
      bram_data_in_muxed = {DATA_WIDTH{1'b0}};
   end
   else
   begin
      WRITE_ADDRESS_REG_muxed = A_r;
      bram_write_en_muxed = bram_wen;
      bram_data_in_muxed = bram_data_in;
   end
end
endmodule
module synchronizer (
    clk,
    presyncdata,
    syncdata
    );
parameter SIZE = 1;
input wire clk;
input wire [SIZE-1:0] presyncdata;
output reg [SIZE-1:0] syncdata;
  reg [SIZE-1:0] presyncdata_tmp = {{SIZE}{1'b0}};
    
    
    
    
    
    
    
    
    
    
    
    
    
    
always @ (posedge clk)
begin
    presyncdata_tmp <= presyncdata;
    syncdata        <= presyncdata_tmp;
end
endmodule
 
module bw_r_rf16x160(
   
   dout, so_w, so_r,
   
   din, rd_adr, wr_adr, read_en, wr_en, rst_tri_en, word_wen,
   byte_wen, rd_clk, wr_clk, se, si_r, si_w, reset_l, sehold
   );
   input [159:0]  din; 
   input [3:0]    rd_adr;   
   input [3:0]    wr_adr;  
   input          read_en;
   input    wr_en;  
        
   input    rst_tri_en ; 
   input [3:0]    word_wen; 
          
   input [19:0]   byte_wen; 
                            
   input          rd_clk;
   input          wr_clk;
   input          se, si_r, si_w ;
   input    reset_l;
   input    sehold; 
   output [159:0] dout;
   output         so_w;
   output         so_r;
   
   wire _unused_ok = &{1'b0,
                      se,
                      si_r,
                      si_w,
                      1'b0};
   wire _unused_output = 1'b0;
   assign so_w = _unused_output;
   assign so_r = _unused_output;
   wire [159:0] bit_en; 
   
   reg [3:0] rd_adr_d1;
   reg [3:0] rd_adr_d2;
   reg [3:0] wr_adr_d1;
   reg wr_en_d1;
   reg [3:0] word_wen_d1;
   reg [19:0] byte_wen_d1;
   reg read_en_d1;
   reg read_en_d2;
   
   reg [159:0] inq_ary [15:0];
   
   assign dout = inq_ary[rd_adr_d1];
   
   always @ (posedge wr_clk)
   begin
      if (!reset_l)
      begin
         
         inq_ary[00] <= 160'b0;
         inq_ary[01] <= 160'b0;
         inq_ary[02] <= 160'b0;
         inq_ary[03] <= 160'b0;
         inq_ary[04] <= 160'b0;
         inq_ary[05] <= 160'b0;
         inq_ary[06] <= 160'b0;
         inq_ary[07] <= 160'b0;
         inq_ary[08] <= 160'b0;
         inq_ary[09] <= 160'b0;
         inq_ary[10] <= 160'b0;
         inq_ary[11] <= 160'b0;
         inq_ary[12] <= 160'b0;
         inq_ary[13] <= 160'b0;
         inq_ary[14] <= 160'b0;
         inq_ary[15] <= 160'b0;
      end
      else
      begin
         if (wr_en)
         begin
            inq_ary[wr_adr] <= (din & bit_en) | (inq_ary[wr_adr] & ~bit_en);
         end
      end
   end
   
   always @ (posedge rd_clk)
   begin
      
      rd_adr_d1 <= rd_adr;
      rd_adr_d2 <= rd_adr_d1;
      wr_adr_d1 <= wr_adr;
      wr_en_d1 <= wr_en;
      word_wen_d1 <= word_wen;
      byte_wen_d1 <= byte_wen;
      read_en_d1 <= read_en;
      read_en_d2 <= read_en_d1;
   end
   assign bit_en[0]  = word_wen[0] & byte_wen[0] & ~rst_tri_en;
   assign bit_en[1]  = word_wen[1] & byte_wen[0] & ~rst_tri_en;
   assign bit_en[2]  = word_wen[2] & byte_wen[0] & ~rst_tri_en;
   assign bit_en[3]  = word_wen[3] & byte_wen[0] & ~rst_tri_en;
   assign bit_en[4]  = word_wen[0] & byte_wen[0] & ~rst_tri_en;
   assign bit_en[5]  = word_wen[1] & byte_wen[0] & ~rst_tri_en;
   assign bit_en[6]  = word_wen[2] & byte_wen[0] & ~rst_tri_en;
   assign bit_en[7]  = word_wen[3] & byte_wen[0] & ~rst_tri_en;
   assign bit_en[8]  = word_wen[0] & byte_wen[1] & ~rst_tri_en;
   assign bit_en[9]  = word_wen[1] & byte_wen[1] & ~rst_tri_en;
   assign bit_en[10] = word_wen[2] & byte_wen[1] & ~rst_tri_en;
   assign bit_en[11] = word_wen[3] & byte_wen[1] & ~rst_tri_en;
   assign bit_en[12] = word_wen[0] & byte_wen[1] & ~rst_tri_en;
   assign bit_en[13] = word_wen[1] & byte_wen[1] & ~rst_tri_en;
   assign bit_en[14] = word_wen[2] & byte_wen[1] & ~rst_tri_en;
   assign bit_en[15] = word_wen[3] & byte_wen[1] & ~rst_tri_en;
   assign bit_en[16] = word_wen[0] & byte_wen[2] & ~rst_tri_en;
   assign bit_en[17] = word_wen[1] & byte_wen[2] & ~rst_tri_en;
   assign bit_en[18] = word_wen[2] & byte_wen[2] & ~rst_tri_en;
   assign bit_en[19] = word_wen[3] & byte_wen[2] & ~rst_tri_en;
   assign bit_en[20] = word_wen[0] & byte_wen[2] & ~rst_tri_en;
   assign bit_en[21] = word_wen[1] & byte_wen[2] & ~rst_tri_en;
   assign bit_en[22] = word_wen[2] & byte_wen[2] & ~rst_tri_en;
   assign bit_en[23] = word_wen[3] & byte_wen[2] & ~rst_tri_en;
   assign bit_en[24] = word_wen[0] & byte_wen[3] & ~rst_tri_en;
   assign bit_en[25] = word_wen[1] & byte_wen[3] & ~rst_tri_en;
   assign bit_en[26] = word_wen[2] & byte_wen[3] & ~rst_tri_en;
   assign bit_en[27] = word_wen[3] & byte_wen[3] & ~rst_tri_en;
   assign bit_en[28] = word_wen[0] & byte_wen[3] & ~rst_tri_en;
   assign bit_en[29] = word_wen[1] & byte_wen[3] & ~rst_tri_en;
   assign bit_en[30] = word_wen[2] & byte_wen[3] & ~rst_tri_en;
   assign bit_en[31] = word_wen[3] & byte_wen[3] & ~rst_tri_en;
   assign bit_en[32] = word_wen[0] & byte_wen[4] & ~rst_tri_en;
   assign bit_en[33] = word_wen[1] & byte_wen[4] & ~rst_tri_en;
   assign bit_en[34] = word_wen[2] & byte_wen[4] & ~rst_tri_en;
   assign bit_en[35] = word_wen[3] & byte_wen[4] & ~rst_tri_en;
   assign bit_en[36] = word_wen[0] & byte_wen[4] & ~rst_tri_en;
   assign bit_en[37] = word_wen[1] & byte_wen[4] & ~rst_tri_en;
   assign bit_en[38] = word_wen[2] & byte_wen[4] & ~rst_tri_en;
   assign bit_en[39] = word_wen[3] & byte_wen[4] & ~rst_tri_en;
   assign bit_en[40] = word_wen[0] & byte_wen[5] & ~rst_tri_en;
   assign bit_en[41] = word_wen[1] & byte_wen[5] & ~rst_tri_en;
   assign bit_en[42] = word_wen[2] & byte_wen[5] & ~rst_tri_en;
   assign bit_en[43] = word_wen[3] & byte_wen[5] & ~rst_tri_en;
   assign bit_en[44] = word_wen[0] & byte_wen[5] & ~rst_tri_en;
   assign bit_en[45] = word_wen[1] & byte_wen[5] & ~rst_tri_en;
   assign bit_en[46] = word_wen[2] & byte_wen[5] & ~rst_tri_en;
   assign bit_en[47] = word_wen[3] & byte_wen[5] & ~rst_tri_en;
   assign bit_en[48] = word_wen[0] & byte_wen[6] & ~rst_tri_en;
   assign bit_en[49] = word_wen[1] & byte_wen[6] & ~rst_tri_en;
   assign bit_en[50] = word_wen[2] & byte_wen[6] & ~rst_tri_en;
   assign bit_en[51] = word_wen[3] & byte_wen[6] & ~rst_tri_en;
   assign bit_en[52] = word_wen[0] & byte_wen[6] & ~rst_tri_en;
   assign bit_en[53] = word_wen[1] & byte_wen[6] & ~rst_tri_en;
   assign bit_en[54] = word_wen[2] & byte_wen[6] & ~rst_tri_en;
   assign bit_en[55] = word_wen[3] & byte_wen[6] & ~rst_tri_en;
   assign bit_en[56] = word_wen[0] & byte_wen[7] & ~rst_tri_en;
   assign bit_en[57] = word_wen[1] & byte_wen[7] & ~rst_tri_en;
   assign bit_en[58] = word_wen[2] & byte_wen[7] & ~rst_tri_en;
   assign bit_en[59] = word_wen[3] & byte_wen[7] & ~rst_tri_en;
   assign bit_en[60] = word_wen[0] & byte_wen[7] & ~rst_tri_en;
   assign bit_en[61] = word_wen[1] & byte_wen[7] & ~rst_tri_en;
   assign bit_en[62] = word_wen[2] & byte_wen[7] & ~rst_tri_en;
   assign bit_en[63] = word_wen[3] & byte_wen[7] & ~rst_tri_en;
   assign bit_en[64] = word_wen[0] & byte_wen[8] & ~rst_tri_en;
   assign bit_en[65] = word_wen[1] & byte_wen[8] & ~rst_tri_en;
   assign bit_en[66] = word_wen[2] & byte_wen[8] & ~rst_tri_en;
   assign bit_en[67] = word_wen[3] & byte_wen[8] & ~rst_tri_en;
   assign bit_en[68] = word_wen[0] & byte_wen[8] & ~rst_tri_en;
   assign bit_en[69] = word_wen[1] & byte_wen[8] & ~rst_tri_en;
   assign bit_en[70] = word_wen[2] & byte_wen[8] & ~rst_tri_en;
   assign bit_en[71] = word_wen[3] & byte_wen[8] & ~rst_tri_en;
   assign bit_en[72] = word_wen[0] & byte_wen[9] & ~rst_tri_en;
   assign bit_en[73] = word_wen[1] & byte_wen[9] & ~rst_tri_en;
   assign bit_en[74] = word_wen[2] & byte_wen[9] & ~rst_tri_en;
   assign bit_en[75] = word_wen[3] & byte_wen[9] & ~rst_tri_en;
   assign bit_en[76] = word_wen[0] & byte_wen[9] & ~rst_tri_en;
   assign bit_en[77] = word_wen[1] & byte_wen[9] & ~rst_tri_en;
   assign bit_en[78] = word_wen[2] & byte_wen[9] & ~rst_tri_en;
   assign bit_en[79] = word_wen[3] & byte_wen[9] & ~rst_tri_en;
   assign bit_en[80] = word_wen[0] & byte_wen[10] & ~rst_tri_en;
   assign bit_en[81] = word_wen[1] & byte_wen[10] & ~rst_tri_en;
   assign bit_en[82] = word_wen[2] & byte_wen[10] & ~rst_tri_en;
   assign bit_en[83] = word_wen[3] & byte_wen[10] & ~rst_tri_en;
   assign bit_en[84] = word_wen[0] & byte_wen[10] & ~rst_tri_en;
   assign bit_en[85] = word_wen[1] & byte_wen[10] & ~rst_tri_en;
   assign bit_en[86] = word_wen[2] & byte_wen[10] & ~rst_tri_en;
   assign bit_en[87] = word_wen[3] & byte_wen[10] & ~rst_tri_en;
   assign bit_en[88] = word_wen[0] & byte_wen[11] & ~rst_tri_en;
   assign bit_en[89] = word_wen[1] & byte_wen[11] & ~rst_tri_en;
   assign bit_en[90] = word_wen[2] & byte_wen[11] & ~rst_tri_en;
   assign bit_en[91] = word_wen[3] & byte_wen[11] & ~rst_tri_en;
   assign bit_en[92] = word_wen[0] & byte_wen[11] & ~rst_tri_en;
   assign bit_en[93] = word_wen[1] & byte_wen[11] & ~rst_tri_en;
   assign bit_en[94] = word_wen[2] & byte_wen[11] & ~rst_tri_en;
   assign bit_en[95] = word_wen[3] & byte_wen[11] & ~rst_tri_en;
   assign bit_en[96] = word_wen[0] & byte_wen[12] & ~rst_tri_en;
   assign bit_en[97] = word_wen[1] & byte_wen[12] & ~rst_tri_en;
   assign bit_en[98] = word_wen[2] & byte_wen[12] & ~rst_tri_en;
   assign bit_en[99] = word_wen[3] & byte_wen[12] & ~rst_tri_en;
   assign bit_en[100] = word_wen[0] & byte_wen[12] & ~rst_tri_en;
   assign bit_en[101] = word_wen[1] & byte_wen[12] & ~rst_tri_en;
   assign bit_en[102] = word_wen[2] & byte_wen[12] & ~rst_tri_en;
   assign bit_en[103] = word_wen[3] & byte_wen[12] & ~rst_tri_en;
   assign bit_en[104] = word_wen[0] & byte_wen[13] & ~rst_tri_en;
   assign bit_en[105] = word_wen[1] & byte_wen[13] & ~rst_tri_en;
   assign bit_en[106] = word_wen[2] & byte_wen[13] & ~rst_tri_en;
   assign bit_en[107] = word_wen[3] & byte_wen[13] & ~rst_tri_en;
   assign bit_en[108] = word_wen[0] & byte_wen[13] & ~rst_tri_en;
   assign bit_en[109] = word_wen[1] & byte_wen[13] & ~rst_tri_en;
   assign bit_en[110] = word_wen[2] & byte_wen[13] & ~rst_tri_en;
   assign bit_en[111] = word_wen[3] & byte_wen[13] & ~rst_tri_en;
   assign bit_en[112] = word_wen[0] & byte_wen[14] & ~rst_tri_en;
   assign bit_en[113] = word_wen[1] & byte_wen[14] & ~rst_tri_en;
   assign bit_en[114] = word_wen[2] & byte_wen[14] & ~rst_tri_en;
   assign bit_en[115] = word_wen[3] & byte_wen[14] & ~rst_tri_en;
   assign bit_en[116] = word_wen[0] & byte_wen[14] & ~rst_tri_en;
   assign bit_en[117] = word_wen[1] & byte_wen[14] & ~rst_tri_en;
   assign bit_en[118] = word_wen[2] & byte_wen[14] & ~rst_tri_en;
   assign bit_en[119] = word_wen[3] & byte_wen[14] & ~rst_tri_en;
   assign bit_en[120] = word_wen[0] & byte_wen[15] & ~rst_tri_en;
   assign bit_en[121] = word_wen[1] & byte_wen[15] & ~rst_tri_en;
   assign bit_en[122] = word_wen[2] & byte_wen[15] & ~rst_tri_en;
   assign bit_en[123] = word_wen[3] & byte_wen[15] & ~rst_tri_en;
   assign bit_en[124] = word_wen[0] & byte_wen[15] & ~rst_tri_en;
   assign bit_en[125] = word_wen[1] & byte_wen[15] & ~rst_tri_en;
   assign bit_en[126] = word_wen[2] & byte_wen[15] & ~rst_tri_en;
   assign bit_en[127] = word_wen[3] & byte_wen[15] & ~rst_tri_en;
   assign bit_en[128] = word_wen[0] & byte_wen[16] & ~rst_tri_en;
   assign bit_en[129] = word_wen[1] & byte_wen[16] & ~rst_tri_en;
   assign bit_en[130] = word_wen[2] & byte_wen[16] & ~rst_tri_en;
   assign bit_en[131] = word_wen[3] & byte_wen[16] & ~rst_tri_en;
   assign bit_en[132] = word_wen[0] & byte_wen[16] & ~rst_tri_en;
   assign bit_en[133] = word_wen[1] & byte_wen[16] & ~rst_tri_en;
   assign bit_en[134] = word_wen[2] & byte_wen[16] & ~rst_tri_en;
   assign bit_en[135] = word_wen[3] & byte_wen[16] & ~rst_tri_en;
   assign bit_en[136] = word_wen[0] & byte_wen[17] & ~rst_tri_en;
   assign bit_en[137] = word_wen[1] & byte_wen[17] & ~rst_tri_en;
   assign bit_en[138] = word_wen[2] & byte_wen[17] & ~rst_tri_en;
   assign bit_en[139] = word_wen[3] & byte_wen[17] & ~rst_tri_en;
   assign bit_en[140] = word_wen[0] & byte_wen[17] & ~rst_tri_en;
   assign bit_en[141] = word_wen[1] & byte_wen[17] & ~rst_tri_en;
   assign bit_en[142] = word_wen[2] & byte_wen[17] & ~rst_tri_en;
   assign bit_en[143] = word_wen[3] & byte_wen[17] & ~rst_tri_en;
   assign bit_en[144] = word_wen[0] & byte_wen[18] & ~rst_tri_en;
   assign bit_en[145] = word_wen[1] & byte_wen[18] & ~rst_tri_en;
   assign bit_en[146] = word_wen[2] & byte_wen[18] & ~rst_tri_en;
   assign bit_en[147] = word_wen[3] & byte_wen[18] & ~rst_tri_en;
   assign bit_en[148] = word_wen[0] & byte_wen[18] & ~rst_tri_en;
   assign bit_en[149] = word_wen[1] & byte_wen[18] & ~rst_tri_en;
   assign bit_en[150] = word_wen[2] & byte_wen[18] & ~rst_tri_en;
   assign bit_en[151] = word_wen[3] & byte_wen[18] & ~rst_tri_en;
   assign bit_en[152] = word_wen[0] & byte_wen[19] & ~rst_tri_en;
   assign bit_en[153] = word_wen[1] & byte_wen[19] & ~rst_tri_en;
   assign bit_en[154] = word_wen[2] & byte_wen[19] & ~rst_tri_en;
   assign bit_en[155] = word_wen[3] & byte_wen[19] & ~rst_tri_en;
   assign bit_en[156] = word_wen[0] & byte_wen[19] & ~rst_tri_en;
   assign bit_en[157] = word_wen[1] & byte_wen[19] & ~rst_tri_en;
   assign bit_en[158] = word_wen[2] & byte_wen[19] & ~rst_tri_en;
   assign bit_en[159] = word_wen[3] & byte_wen[19] & ~rst_tri_en;
endmodule
module clk_mux (
    input       clk0_p,
    input       clk0_n,
    input       clk1_p,
    input       clk1_n,
    input       clk2,
    input [1:0] sel,
    output      clk_muxed
);
assign clk_muxed = clk0_p;
endmodule
module clk_se_to_diff (
    input   clk_se,
    output  clk_p,
    output  clk_n
);
assign clk_p = clk_se;
assign clk_n = 1'bx;
endmodule
 
 
 
 
 
 
 
 
 
 
 
 module pll_top ( 
   output clk_locked,
   output clk_out,
   input ref_clk,
   input rst,
   input bypass_en,
   input [4:0] rangeA
);
assign clk_out = ref_clk;
assign clk_locked = ~rst;
endmodule
  
          
      
    
         
module rtap(
    input wire clk,
    input wire rst_n,
    input wire [8-1:0] own_tileid,
    
    
    output wire tile_jtag_ucb_val,
    output wire [4-1:0] tile_jtag_ucb_data,
    
    input wire jtag_tiles_ucb_val,
    input wire [4-1:0] jtag_tiles_ucb_data,
    
    
    input wire [4-1:0] srams_rtap_data,
    output reg [4-1:0] rtap_srams_bist_command,
    output reg [4-1:0] rtap_srams_bist_data,
    
    
    output reg               rtap_arb_req_val,
    output reg [63:0]        rtap_arb_req_data,
    output reg [1:0]         rtap_arb_req_threadid,
    
    
    input wire [94-1:0] core_rtap_data,
    output reg rtap_core_val,
    output reg [1:0] rtap_core_threadid,
    output reg [4-1:0]  rtap_core_id,
    output reg [94-1:0] rtap_core_data,
    
    
    output reg rtap_config_req_val,
    output reg rtap_config_req_rw,
    output reg [63:0] rtap_config_write_req_data,
    output reg [15:8] rtap_config_req_address,
    input wire [63:0] config_rtap_read_res_data
    );
wire ucb_rx_val;
wire [128-1:0] ucb_rx_data;
reg ucb_tx_val;
reg [128-1:0] ucb_tx_data;
reg [(128/4)-1:0] ucb_tx_data_vec;
reg req_val;
reg [32-1:0] req_header;
reg [8-1:0] req_op;
reg [16-1:0] req_misc;
reg [6-1:0] req_tileid;
reg [2-1:0] req_threadid;
reg [32-1:0] req_address;
reg [16:0] req_address_index;
reg [8:0] req_address_sramid;
reg [8:0] req_address_bsel;
reg [63:0] req_data;
reg [4-1:0] res_op_next;
reg [4-1:0] res_op;
reg res_val;
reg sram_res_val;
reg sram_res_val_f;
always @ (posedge clk)
begin
    if (!rst_n)
        sram_res_val_f <= 1'b0;
    else
        sram_res_val_f <= sram_res_val;
end
reg [4-1:0] sram_req_op;
reg [4-1:0] sram_req_dataout;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        rtap_srams_bist_command <= 4'd0;
    end
    else
    begin
        rtap_srams_bist_command <= sram_req_op;
    end
    rtap_srams_bist_data <= sram_req_dataout;
end
reg [15:0] sram_req_address_reg;
reg [3:0] sram_req_sramid_reg;
reg [63:0] sram_data_reg;
reg [7:0] sram_req_bsel_reg;
reg [15:0] sram_req_address_reg_next;
reg [3:0] sram_req_sramid_reg_next;
reg [63:0] sram_data_reg_next;
reg [7:0] sram_req_bsel_reg_next;
reg sram_req_rw;
reg sram_req_rw_next;
reg judi_op_val;
reg [1:0] judi_op_threadid;
reg [4-1:0] judi_op_id;
reg [94-1:0] judi_op_data;
always @ (posedge clk)
begin
    if (!rst_n)
        rtap_core_val <= 1'b0;
    else
        rtap_core_val <= judi_op_val;
    rtap_core_data <= judi_op_data;
    rtap_core_threadid <= judi_op_threadid;
    rtap_core_id <= judi_op_id;
end
wire judi_op_val_f = rtap_core_val;
reg judi_op_val_ff;
always @ (posedge clk)
begin
    judi_op_val_ff <= judi_op_val_f;
end
reg [4-1:0] state;
reg [4-1:0] state_next;
reg [3:0] state_counter;
reg [3:0] state_counter_next;
reg [3:0] state_counter_minus_1;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        state <= 4'd0;
        res_op <= 0;
    end
    else
    begin
        state <= state_next;
        state_counter <= state_counter_next;
        res_op <= res_op_next;
    end
end
always @ *
begin
    req_data = ucb_rx_data[127:64];
    req_address = ucb_rx_data[63:32];
    req_header = ucb_rx_data[31:0];
    req_op = 0;
    req_tileid = req_header[23:18];
    req_threadid = req_header[17:16];
    req_misc = req_header[15:0];
    req_address_index = req_address[15:0];
    req_address_sramid = req_address[31:24];
    req_address_bsel = req_address[23:16];
    req_val = ucb_rx_val && (req_tileid == 6'b111111 || req_tileid == own_tileid);
    if (req_val)
        req_op = req_header[31:24];
    res_op_next = 0;
    
    sram_req_address_reg_next = sram_req_address_reg;
    sram_req_sramid_reg_next = sram_req_sramid_reg;
    sram_data_reg_next = sram_data_reg;
    sram_req_bsel_reg_next = sram_req_bsel_reg;
    sram_req_rw_next = sram_req_rw;
    sram_req_op = 0;
    sram_req_dataout = 0;
    sram_res_val = 1'b0;
    state_counter_minus_1 = state_counter - 1;
    state_counter_next = state_counter;
    state_next = 4'd0;
    case (state)
        4'd0:
        begin
            if (req_op == 8'd4 || req_op == 8'd5)
            begin
                
                sram_req_address_reg_next[15:0] = req_address_index[15:0];
                sram_req_sramid_reg_next[3:0] = req_address_sramid;
                sram_req_bsel_reg_next[7:0] = req_address_bsel;
                state_next = 4'd1;
                state_counter_next = 0; 
                if (req_op == 8'd4)
                    sram_req_rw_next = 1'b0;
                else
                begin
                    sram_req_rw_next = 1'b1;
                    sram_data_reg_next = req_data[63:0];
                end
            end
        end
        4'd1:
        begin
            
            sram_req_op = 4'd6;
            sram_req_dataout[3:0] = sram_req_sramid_reg[3:0];
            if (state_counter == 0)
            begin
                state_next = 4'd2;
                state_counter_next = 1; 
            end
            else
            begin
                state_next = state;
                state_counter_next = state_counter_minus_1;
            end
        end
        4'd2:
        begin
            
            sram_req_op = 4'd7;
            sram_req_dataout[3:0] = sram_req_bsel_reg[7:4];
            sram_req_bsel_reg_next = {sram_req_bsel_reg[3:0], 4'b0};
            if (state_counter == 0)
            begin
                state_next = 4'd3;
                state_counter_next = 3; 
            end
            else
            begin
                state_next = state;
                state_counter_next = state_counter_minus_1;
            end
        end
        4'd3:
        begin
            
            sram_req_op = 4'd5;
            sram_req_dataout[3:0] = sram_req_address_reg[15:12];
            sram_req_address_reg_next = {sram_req_address_reg[11:0], 4'b0};
            if (state_counter == 0)
            begin
                if (sram_req_rw == 1'b0)
                begin
                    state_next = 4'd4;
                end
                else
                    state_next = 4'd7;
                    state_counter_next = 15; 
            end
            else
            begin
                state_next = state;
                state_counter_next = state_counter_minus_1;
            end
        end
        4'd4:
        begin
            
            sram_req_op = 4'd1;
            state_next = 4'd5;
        end
        4'd5:
        begin
            
            sram_req_op = 0;
            state_next = 4'd9;
            
        end
        4'd9:
        begin
            
            sram_req_op = 4'd4;
            state_next = 4'd6;
            state_counter_next = 15; 
        end
        4'd6:
        begin
            
            sram_req_op = 4'd4;
            sram_req_dataout[3:0] = sram_data_reg[63:60]; 
            sram_data_reg_next = {sram_data_reg[59:0], srams_rtap_data[3:0]};
            if (state_counter == 0)
            begin
                state_next = 4'd0;
                
                sram_res_val = 1'b1;
            end
            else
            begin
                state_next = state;
                state_counter_next = state_counter_minus_1;
            end
        end
        4'd7:
        begin
            
            sram_req_op = 4'd4;
            sram_req_dataout[3:0] = sram_data_reg[63:60];
            sram_data_reg_next = {sram_data_reg[59:0], srams_rtap_data[3:0]};
            if (state_counter == 0)
            begin
                state_next = 4'd8;
            end
            else
            begin
                state_next = state;
                state_counter_next = state_counter_minus_1;
            end
        end
        4'd8:
        begin
            
            sram_req_op = 4'd2;
            
            sram_res_val = 1'b1;
            state_next = 4'd0;
        end
    endcase
    rtap_arb_req_val = 0;
    rtap_arb_req_data[63:0] = 0;
    rtap_arb_req_threadid[1:0] = 0;
    judi_op_val = 0;
    judi_op_threadid = 0;
    judi_op_id = 0;
    judi_op_data = 0;
    rtap_config_req_val = 0;
    rtap_config_req_rw = 0;
    rtap_config_req_address = 0;
    rtap_config_write_req_data = 0;
    case (req_op)
        
        
        
        
        
        
        
        8'd10:
        begin
            case (req_misc)
                16'd7:
                begin
                    res_op_next = 4'd4;
                    rtap_config_req_val = 1'b1;
                    rtap_config_req_rw = 1'b0;
                    rtap_config_req_address[15:8] = req_address;
                end
                16'd8:
                begin
                    
                    judi_op_threadid = req_threadid;
                    judi_op_val = 1'b1;
                    judi_op_id = 4'd5;
                end
                16'd9:
                begin
                    
                    judi_op_threadid = req_threadid;
                    judi_op_val = 1'b1;
                    judi_op_id = 4'd6;
                    judi_op_data = req_address;
                end
            endcase
        end
        8'd11:
        begin
            case (req_misc)
                16'd1:
                begin
                    
                    judi_op_threadid = req_threadid;
                    judi_op_val = 1'b1;
                    judi_op_id = 4'd3;
                    judi_op_data[47:0] = req_data[47:0];
                end
                16'd5:
                begin
                    
                    judi_op_data[47:0] = req_data[47:0];
                    judi_op_threadid = req_threadid;
                    judi_op_val = 1'b1;
                    judi_op_id = 4'd4;
                end
                16'd3:
                begin
                    
                    judi_op_threadid = req_threadid;
                    judi_op_val = 1'b1;
                    judi_op_id = 4'd2;
                    judi_op_data[4:0] = req_data[4:0];
                end
                16'd6:
                begin
                    
                    judi_op_threadid = req_threadid;
                    judi_op_val = 1'b1;
                    judi_op_id = 4'd1;
                    judi_op_data[13:0] = req_data[13:0];
                end
                16'd4:
                begin
                    res_op_next = 4'd1;
                    rtap_arb_req_val = 1'b1;
                    rtap_arb_req_data[63:0] = req_data[63:0];
                    rtap_arb_req_threadid[1:0] = req_threadid[1:0];
                end
                16'd7:
                begin
                    res_op_next = 4'd1;
                    rtap_config_req_val = 1'b1;
                    rtap_config_req_rw = 1'b1;
                    rtap_config_req_address[15:8] = req_address;
                    rtap_config_write_req_data = req_data;
                end
                16'd10:
                begin
                    
                    
                    judi_op_val = 1'b1;
                    judi_op_id = 4'd8;
                    judi_op_data[4:0] = req_data[4:0]; 
                end
                16'd11:
                begin
                    
                    
                    
                    
                    judi_op_val = 1'b1;
                    judi_op_id = 4'd7;
                    judi_op_data[47:0] = req_data[47:0]; 
                end
            endcase
        end
    endcase
end
always @ (posedge clk)
begin
    sram_req_address_reg <= sram_req_address_reg_next;
    sram_req_sramid_reg <= sram_req_sramid_reg_next;
    sram_data_reg <= sram_data_reg_next;
    sram_req_bsel_reg <= sram_req_bsel_reg_next;
    sram_req_rw <= sram_req_rw_next;
end
reg [128-1:0] res_data;
always @ *
begin
    res_val = 0;
    res_data = 0;
    
    if (judi_op_val_ff)
    begin
        res_val = 1'b1;
        res_data = core_rtap_data[94-1:0];
    end
    else
    if (sram_res_val_f)
    begin
        res_val = 1'b1;
        res_data = sram_data_reg;
    end
    else case (res_op)
        4'd1:
        begin
            res_val = 1'b1;
        end
        
        
        
        
        
        
        
        
        
        
        4'd4:
        begin
            res_val = 1'b1;
            res_data = config_rtap_read_res_data;
        end
    endcase
    ucb_tx_val = res_val;
    ucb_tx_data_vec = 32'hffffffff;
    ucb_tx_data = res_data;
end
rtap_ucb_receiver ucb_rx(
    .clk(clk),
    .rst_n(rst_n),
    .ucb_rx_val(ucb_rx_val),
    .ucb_rx_data(ucb_rx_data),
    .ucb_in_vld(jtag_tiles_ucb_val),
    .ucb_in_data(jtag_tiles_ucb_data)
    );
rtap_ucb_transmitter ucb_tx(
    .clk(clk),
    .rst_n(rst_n),
    .ucb_tx_val(ucb_tx_val),
    .ucb_tx_data(ucb_tx_data),
    .ucb_tx_data_vec(ucb_tx_data_vec),
    .ucb_out_val(tile_jtag_ucb_val),
    .ucb_out_data(tile_jtag_ucb_data)
    );
endmodule
  
          
      
    
         
module rtap_ucb_receiver(
    input wire clk,
    input wire rst_n,
    
    output wire ucb_rx_val,
    output wire [128-1:0] ucb_rx_data,
    
    
    input wire ucb_in_vld,
    
    input wire [4-1:0] ucb_in_data
    );
ucb_bus_in #(4, 128-64) ucb_in_tile0(
    .vld(ucb_in_vld),
    .data(ucb_in_data),
    .stall(),
    .clk(clk),
    .rst_l(rst_n),
    .indata_buf_vld(ucb_rx_val),
    .indata_buf(ucb_rx_data),
    .stall_a1(1'b0)
    );
endmodule
  
          
      
    
         
module rtap_ucb_transmitter(
    input wire clk,
    input wire rst_n,
    
    input wire ucb_tx_val,
    input wire [128-1:0] ucb_tx_data,
    input wire [(128/4)-1:0] ucb_tx_data_vec,
    
    
    output wire ucb_out_val,
    
    output wire [4-1:0] ucb_out_data
    );
ucb_bus_out #(4, 128-64) ucb_out(
    .vld(ucb_out_val),
    .data(ucb_out_data),
    .outdata_buf_busy(),
    .clk(clk),
    .rst_l(rst_n),
    .stall(1'b0),
    .outdata_buf_in(ucb_tx_data),
    .outdata_vec_in(ucb_tx_data_vec),
    .outdata_buf_wr(ucb_tx_val)
    );
endmodule
module axi2mem #(
    parameter int unsigned AXI_ID_WIDTH      = 10,
    parameter int unsigned AXI_ADDR_WIDTH    = 64,
    parameter int unsigned AXI_DATA_WIDTH    = 64,
    parameter int unsigned AXI_USER_WIDTH    = 10
)(
    input logic                         clk_i,    
    input logic                         rst_ni,  
    AXI_BUS.Slave                       slave,
    output logic                        req_o,
    output logic                        we_o,
    output logic [AXI_ADDR_WIDTH-1:0]   addr_o,
    output logic [AXI_DATA_WIDTH/8-1:0] be_o,
    output logic [AXI_DATA_WIDTH-1:0]   data_o,
    input  logic [AXI_DATA_WIDTH-1:0]   data_i
);
    
    
    
    
    typedef enum logic [1:0] { FIXED = 2'b00, INCR = 2'b01, WRAP = 2'b10} axi_burst_t;
    localparam LOG_NR_BYTES = $clog2(AXI_DATA_WIDTH/8);
    typedef struct packed {
        logic [AXI_ID_WIDTH-1:0]   id;
        logic [AXI_ADDR_WIDTH-1:0] addr;
        logic [7:0]                len;
        logic [2:0]                size;
        axi_burst_t                burst;
    } ax_req_t;
    
    enum logic [2:0] { IDLE, READ, WRITE, SEND_B, WAIT_WVALID }  state_d, state_q;
    ax_req_t                   ax_req_d, ax_req_q;
    logic [AXI_ADDR_WIDTH-1:0] req_addr_d, req_addr_q;
    logic [7:0]                cnt_d, cnt_q;
    function automatic logic [AXI_ADDR_WIDTH-1:0] get_wrap_bounadry (input logic [AXI_ADDR_WIDTH-1:0] unaligned_address, input logic [7:0] len);
        logic [AXI_ADDR_WIDTH-1:0] warp_address = '0;
        
        if (len == 4'b1)
            warp_address[AXI_ADDR_WIDTH-1:1+LOG_NR_BYTES] = unaligned_address[AXI_ADDR_WIDTH-1:1+LOG_NR_BYTES];
        else if (len == 4'b11)
            warp_address[AXI_ADDR_WIDTH-1:2+LOG_NR_BYTES] = unaligned_address[AXI_ADDR_WIDTH-1:2+LOG_NR_BYTES];
        else if (len == 4'b111)
            warp_address[AXI_ADDR_WIDTH-1:3+LOG_NR_BYTES] = unaligned_address[AXI_ADDR_WIDTH-3:2+LOG_NR_BYTES];
        else if (len == 4'b1111)
            warp_address[AXI_ADDR_WIDTH-1:4+LOG_NR_BYTES] = unaligned_address[AXI_ADDR_WIDTH-3:4+LOG_NR_BYTES];
        return warp_address;
    endfunction
    logic [AXI_ADDR_WIDTH-1:0] aligned_address;
    logic [AXI_ADDR_WIDTH-1:0] wrap_boundary;
    logic [AXI_ADDR_WIDTH-1:0] upper_wrap_boundary;
    logic [AXI_ADDR_WIDTH-1:0] cons_addr;
    always_comb begin
        
        aligned_address = {ax_req_q.addr[AXI_ADDR_WIDTH-1:LOG_NR_BYTES], {{LOG_NR_BYTES}{1'b0}}};
        wrap_boundary = get_wrap_bounadry(ax_req_q.addr, ax_req_q.len);
        
        upper_wrap_boundary = wrap_boundary + ((ax_req_q.len + 1) << LOG_NR_BYTES);
        
        cons_addr = aligned_address + (cnt_q << LOG_NR_BYTES);
        
        
        state_d    = state_q;
        ax_req_d   = ax_req_q;
        req_addr_d = req_addr_q;
        cnt_d      = cnt_q;
        
        data_o = slave.w_data;
        be_o   = slave.w_strb;
        we_o   = 1'b0;
        req_o  = 1'b0;
        addr_o = '0;
        
        
        slave.aw_ready = 1'b0;
        slave.ar_ready = 1'b0;
        
        slave.r_valid  = 1'b0;
        slave.r_data   = data_i;
        slave.r_resp   = '0;
        slave.r_last   = '0;
        slave.r_id     = ax_req_q.id;
        slave.r_user   = '0;
        
        slave.w_ready  = 1'b0;
        
        slave.b_valid  = 1'b0;
        slave.b_resp   = 1'b0;
        slave.b_id     = 1'b0;
        slave.b_user   = 1'b0;
        case (state_q)
            IDLE: begin
                
                
                
                
                if (slave.ar_valid) begin
                    slave.ar_ready = 1'b1;
                    
                    ax_req_d       = {slave.ar_id, slave.ar_addr, slave.ar_len, slave.ar_size, slave.ar_burst};
                    state_d        = READ;
                    
                    req_o          = 1'b1;
                    addr_o         = slave.ar_addr;
                    
                    req_addr_d     = slave.ar_addr;
                    
                    cnt_d          = 1;
                
                
                
                end else if (slave.aw_valid) begin
                    slave.aw_ready = 1'b1;
                    slave.w_ready  = 1'b1;
                    addr_o         = slave.aw_addr;
                    
                    ax_req_d       = {slave.aw_id, slave.aw_addr, slave.aw_len, slave.aw_size, slave.aw_burst};
                    
                    if (slave.w_valid) begin
                        req_o          = 1'b1;
                        we_o           = 1'b1;
                        state_d        = (slave.w_last) ? SEND_B : WRITE;
                        cnt_d          = 1;
                    
                    end else
                        state_d = WAIT_WVALID;
                end
            end
            
            WAIT_WVALID: begin
                slave.w_ready = 1'b1;
                addr_o = ax_req_q.addr;
                
                if (slave.w_valid) begin
                    req_o          = 1'b1;
                    we_o           = 1'b1;
                    state_d        = (slave.w_last) ? SEND_B : WRITE;
                    cnt_d          = 1;
                end
            end
            READ: begin
                
                req_o  = 1'b1;
                addr_o = req_addr_q;
                
                slave.r_valid = 1'b1;
                slave.r_data  = data_i;
                slave.r_id    = ax_req_q.id;
                slave.r_last  = (cnt_q == ax_req_q.len + 1);
                
                if (slave.r_ready) begin
                    
                    
                    
                    
                    case (ax_req_q.burst)
                        FIXED, INCR: addr_o = cons_addr;
                        WRAP:  begin
                            
                            if (cons_addr == upper_wrap_boundary) begin
                                addr_o = wrap_boundary;
                            
                            end else if (cons_addr > upper_wrap_boundary) begin
                                addr_o = ax_req_q.addr + ((cnt_q - ax_req_q.len) << LOG_NR_BYTES);
                            
                            end else begin
                                addr_o = cons_addr;
                            end
                        end
                    endcase
                    
                    
                    if (slave.r_last) begin
                        state_d = IDLE;
                        
                        req_o = 1'b0;
                    end
                    
                    req_addr_d = addr_o;
                    
                    cnt_d = cnt_q + 1;
                    
                end
            end
            
            WRITE: begin
                slave.w_ready = 1'b1;
                
                if (slave.w_valid) begin
                    req_o         = 1'b1;
                    we_o          = 1'b1;
                    
                    
                    
                    
                    case (ax_req_q.burst)
                        FIXED, INCR: addr_o = cons_addr;
                        WRAP:  begin
                            
                            if (cons_addr == upper_wrap_boundary) begin
                                addr_o = wrap_boundary;
                            
                            end else if (cons_addr > upper_wrap_boundary) begin
                                addr_o = ax_req_q.addr + ((cnt_q - ax_req_q.len) << LOG_NR_BYTES);
                            
                            end else begin
                                addr_o = cons_addr;
                            end
                        end
                    endcase
                    
                    req_addr_d = addr_o;
                    
                    cnt_d = cnt_q + 1;
                    if (slave.w_last)
                        state_d = SEND_B;
                end
            end
            
            SEND_B: begin
                slave.b_valid = 1'b1;
                slave.b_id    = ax_req_q.id;
                if (slave.b_ready)
                    state_d = IDLE;
            end
        endcase
    end
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (~rst_ni) begin
            state_q    <= IDLE;
            ax_req_q  <= '0;
            req_addr_q <= '0;
            cnt_q      <= '0;
        end else begin
            state_q    <= state_d;
            ax_req_q   <= ax_req_d;
            req_addr_q <= req_addr_d;
            cnt_q      <= cnt_d;
        end
    end
endmodule
module axi_mem_if
#(
    parameter int unsigned AXI4_ADDRESS_WIDTH = 64,
    parameter int unsigned AXI4_RDATA_WIDTH   = 64,
    parameter int unsigned AXI4_WDATA_WIDTH   = 64,
    parameter int unsigned AXI4_ID_WIDTH      = 16,
    parameter int unsigned AXI4_USER_WIDTH    = 10,
    parameter int unsigned AXI_NUMBYTES       = AXI4_WDATA_WIDTH/8,
    parameter int unsigned BUFF_DEPTH_SLAVE   = 4
)
(
    input logic                                     ACLK,
    input logic                                     ARESETn,
    input logic                                     test_en_i,
    
    input  logic [AXI4_ID_WIDTH-1:0]                AWID_i     ,
    input  logic [AXI4_ADDRESS_WIDTH-1:0]           AWADDR_i   ,
    input  logic [ 7:0]                             AWLEN_i    ,
    input  logic [ 2:0]                             AWSIZE_i   ,
    input  logic [ 1:0]                             AWBURST_i  ,
    input  logic                                    AWLOCK_i   ,
    input  logic [ 3:0]                             AWCACHE_i  ,
    input  logic [ 2:0]                             AWPROT_i   ,
    input  logic [ 3:0]                             AWREGION_i ,
    input  logic [ AXI4_USER_WIDTH-1:0]             AWUSER_i   ,
    input  logic [ 3:0]                             AWQOS_i    ,
    input  logic                                    AWVALID_i  ,
    output logic                                    AWREADY_o  ,
    
    input  logic [AXI_NUMBYTES-1:0][7:0]            WDATA_i    ,
    input  logic [AXI_NUMBYTES-1:0]                 WSTRB_i    ,
    input  logic                                    WLAST_i    ,
    input  logic [AXI4_USER_WIDTH-1:0]              WUSER_i    ,
    input  logic                                    WVALID_i   ,
    output logic                                    WREADY_o   ,
    
    output logic   [AXI4_ID_WIDTH-1:0]              BID_o      ,
    output logic   [ 1:0]                           BRESP_o    ,
    output logic                                    BVALID_o   ,
    output logic   [AXI4_USER_WIDTH-1:0]            BUSER_o    ,
    input  logic                                    BREADY_i   ,
    
    input  logic [AXI4_ID_WIDTH-1:0]                ARID_i     ,
    input  logic [AXI4_ADDRESS_WIDTH-1:0]           ARADDR_i   ,
    input  logic [ 7:0]                             ARLEN_i    ,
    input  logic [ 2:0]                             ARSIZE_i   ,
    input  logic [ 1:0]                             ARBURST_i  ,
    input  logic                                    ARLOCK_i   ,
    input  logic [ 3:0]                             ARCACHE_i  ,
    input  logic [ 2:0]                             ARPROT_i   ,
    input  logic [ 3:0]                             ARREGION_i ,
    input  logic [ AXI4_USER_WIDTH-1:0]             ARUSER_i   ,
    input  logic [ 3:0]                             ARQOS_i    ,
    input  logic                                    ARVALID_i  ,
    output logic                                    ARREADY_o  ,
    
    output  logic [AXI4_ID_WIDTH-1:0]               RID_o      ,
    output  logic [AXI4_RDATA_WIDTH-1:0]            RDATA_o    ,
    output  logic [ 1:0]                            RRESP_o    ,
    output  logic                                   RLAST_o    ,
    output  logic [AXI4_USER_WIDTH-1:0]             RUSER_o    ,
    output  logic                                   RVALID_o   ,
    input   logic                                   RREADY_i   ,
    
    output logic                                    CEN        ,
    output logic                                    WEN        ,
    output logic  [AXI4_ADDRESS_WIDTH-1:0]          A          ,
    output logic  [AXI4_WDATA_WIDTH-1:0]            D          ,
    output logic  [AXI_NUMBYTES-1:0]                BE         ,
    input  logic  [AXI4_RDATA_WIDTH-1:0]            Q
);
    
    localparam ADDRESS_BITS= $clog2(AXI4_WDATA_WIDTH/8);
  
  
  
  
  logic [AXI4_ID_WIDTH-1:0]                         AWID       ;
  logic [AXI4_ADDRESS_WIDTH-1:0]                    AWADDR     ;
  logic [ 7:0]                                      AWLEN      ;
  logic [ 2:0]                                      AWSIZE     ;
  logic [ 1:0]                                      AWBURST    ;
  logic                                             AWLOCK     ;
  logic [ 3:0]                                      AWCACHE    ;
  logic [ 2:0]                                      AWPROT     ;
  logic [ 3:0]                                      AWREGION   ;
  logic [ AXI4_USER_WIDTH-1:0]                      AWUSER     ;
  logic [ 3:0]                                      AWQOS      ;
  logic                                             AWVALID    ;
  logic                                             AWREADY    ;
  
  logic [AXI_NUMBYTES-1:0][7:0]                     WDATA      ;
  logic [AXI_NUMBYTES-1:0]                          WSTRB      ;
  logic                                             WLAST      ;
  logic [AXI4_USER_WIDTH-1:0]                       WUSER      ;
  logic                                             WVALID     ;
  logic                                             WREADY     ;
  
  logic   [AXI4_ID_WIDTH-1:0]                       BID        ;
  logic   [ 1:0]                                    BRESP      ;
  logic                                             BVALID     ;
  logic   [AXI4_USER_WIDTH-1:0]                     BUSER      ;
  logic                                             BREADY     ;
  
  logic [AXI4_ID_WIDTH-1:0]                         ARID       ;
  logic [AXI4_ADDRESS_WIDTH-1:0]                    ARADDR     ;
  logic [ 7:0]                                      ARLEN      ;
  logic [ 2:0]                                      ARSIZE     ;
  logic [ 1:0]                                      ARBURST    ;
  logic                                             ARLOCK     ;
  logic [ 3:0]                                      ARCACHE    ;
  logic [ 2:0]                                      ARPROT     ;
  logic [ 3:0]                                      ARREGION   ;
  logic [ AXI4_USER_WIDTH-1:0]                      ARUSER     ;
  logic [ 3:0]                                      ARQOS      ;
  logic                                             ARVALID    ;
  logic                                             ARREADY    ;
  
  logic [AXI4_ID_WIDTH-1:0]                         RID        ;
  logic [AXI4_RDATA_WIDTH-1:0]                      RDATA      ;
  logic [ 1:0]                                      RRESP      ;
  logic                                             RLAST      ;
  logic [AXI4_USER_WIDTH-1:0]                       RUSER      ;
  logic                                             RVALID     ;
  logic                                             RREADY     ;
  enum logic [3:0] { IDLE,
                     SINGLE_RD, BURST_RD, WRAP_RD,
                     BURST_WR, SINGLE_WR, WRAP_WR,
                     WAIT_WDATA_BURST,
                     WAIT_WDATA_SINGLE,
                     WAIT_WDATA_BURST_WRAP,
                     BURST_RESP
                    } CS , NS;
  logic [8:0]                      CountBurstCS;
  logic [8:0]                      CountBurstNS;
  logic [AXI4_ADDRESS_WIDTH-1:0]   address;
  logic [AXI4_ADDRESS_WIDTH-1:0]   address_q;
  logic                            read_req;
  logic                            sample_AR;
  logic [AXI4_ADDRESS_WIDTH-1:0]   ARADDR_Q;
  logic [7:0]                      ARLEN_Q;
  logic [63:0]                     arlen_fixed_q;
  logic                            decr_ARLEN;
  logic [AXI4_ID_WIDTH-1:0]        ARID_Q;
  logic [ AXI4_USER_WIDTH-1:0]     ARUSER_Q;
  logic                            write_req;
  logic                            sample_AW;
  logic [AXI4_ADDRESS_WIDTH-1:0]   AWADDR_Q;
  logic [7:0]                      AWLEN_Q;
  logic [63:0]                     awlen_fixed_q;
  logic                            decr_AWLEN;
  logic [AXI4_ID_WIDTH-1:0]        AWID_Q;
  logic [ AXI4_USER_WIDTH-1:0]     AWUSER_Q;
  logic                            RR_FLAG;
  logic [2:0]                      ar_size_q;
  logic [2:0]                      aw_size_q;
   
   axi_aw_buffer #(
       .ID_WIDTH     ( AXI4_ID_WIDTH      ),
       .ADDR_WIDTH   ( AXI4_ADDRESS_WIDTH ),
       .USER_WIDTH   ( AXI4_USER_WIDTH    ),
       .BUFFER_DEPTH ( BUFF_DEPTH_SLAVE   )
   ) slave_aw_buffer_i (
      .clk_i           ( ACLK        ),
      .rst_ni          ( ARESETn     ),
      .test_en_i       ( test_en_i   ),
      .slave_valid_i   ( AWVALID_i   ),
      .slave_addr_i    ( AWADDR_i    ),
      .slave_prot_i    ( AWPROT_i    ),
      .slave_region_i  ( AWREGION_i  ),
      .slave_len_i     ( AWLEN_i     ),
      .slave_size_i    ( AWSIZE_i    ),
      .slave_burst_i   ( AWBURST_i   ),
      .slave_lock_i    ( AWLOCK_i    ),
      .slave_cache_i   ( AWCACHE_i   ),
      .slave_qos_i     ( AWQOS_i     ),
      .slave_id_i      ( AWID_i      ),
      .slave_user_i    ( AWUSER_i    ),
      .slave_ready_o   ( AWREADY_o   ),
      .master_valid_o  ( AWVALID     ),
      .master_addr_o   ( AWADDR      ),
      .master_prot_o   ( AWPROT      ),
      .master_region_o ( AWREGION    ),
      .master_len_o    ( AWLEN       ),
      .master_size_o   ( AWSIZE      ),
      .master_burst_o  ( AWBURST     ),
      .master_lock_o   ( AWLOCK      ),
      .master_cache_o  ( AWCACHE     ),
      .master_qos_o    ( AWQOS       ),
      .master_id_o     ( AWID        ),
      .master_user_o   ( AWUSER      ),
      .master_ready_i  ( AWREADY     )
   );
   
   axi_ar_buffer #(
       .ID_WIDTH     ( AXI4_ID_WIDTH      ),
       .ADDR_WIDTH   ( AXI4_ADDRESS_WIDTH ),
       .USER_WIDTH   ( AXI4_USER_WIDTH    ),
       .BUFFER_DEPTH ( BUFF_DEPTH_SLAVE   )
   ) slave_ar_buffer_i (
      .clk_i           ( ACLK       ),
      .rst_ni          ( ARESETn    ),
      .test_en_i       ( test_en_i  ),
      .slave_valid_i   ( ARVALID_i  ),
      .slave_addr_i    ( ARADDR_i   ),
      .slave_prot_i    ( ARPROT_i   ),
      .slave_region_i  ( ARREGION_i ),
      .slave_len_i     ( ARLEN_i    ),
      .slave_size_i    ( ARSIZE_i   ),
      .slave_burst_i   ( ARBURST_i  ),
      .slave_lock_i    ( ARLOCK_i   ),
      .slave_cache_i   ( ARCACHE_i  ),
      .slave_qos_i     ( ARQOS_i    ),
      .slave_id_i      ( ARID_i     ),
      .slave_user_i    ( ARUSER_i   ),
      .slave_ready_o   ( ARREADY_o  ),
      .master_valid_o  ( ARVALID    ),
      .master_addr_o   ( ARADDR     ),
      .master_prot_o   ( ARPROT     ),
      .master_region_o ( ARREGION   ),
      .master_len_o    ( ARLEN      ),
      .master_size_o   ( ARSIZE     ),
      .master_burst_o  ( ARBURST    ),
      .master_lock_o   ( ARLOCK     ),
      .master_cache_o  ( ARCACHE    ),
      .master_qos_o    ( ARQOS      ),
      .master_id_o     ( ARID       ),
      .master_user_o   ( ARUSER     ),
      .master_ready_i  ( ARREADY    )
   );
   axi_w_buffer #(
       .DATA_WIDTH(AXI4_WDATA_WIDTH),
       .USER_WIDTH(AXI4_USER_WIDTH),
       .BUFFER_DEPTH(BUFF_DEPTH_SLAVE)
   ) slave_w_buffer_i (
        .clk_i          ( ACLK      ),
        .rst_ni         ( ARESETn   ),
        .test_en_i      ( test_en_i ),
        .slave_valid_i  ( WVALID_i  ),
        .slave_data_i   ( WDATA_i   ),
        .slave_strb_i   ( WSTRB_i   ),
        .slave_user_i   ( WUSER_i   ),
        .slave_last_i   ( WLAST_i   ),
        .slave_ready_o  ( WREADY_o  ),
        .master_valid_o ( WVALID    ),
        .master_data_o  ( WDATA     ),
        .master_strb_o  ( WSTRB     ),
        .master_user_o  ( WUSER     ),
        .master_last_o  ( WLAST     ),
        .master_ready_i ( WREADY    )
    );
   axi_r_buffer #(
        .ID_WIDTH(AXI4_ID_WIDTH),
        .DATA_WIDTH(AXI4_RDATA_WIDTH),
        .USER_WIDTH(AXI4_USER_WIDTH),
        .BUFFER_DEPTH(BUFF_DEPTH_SLAVE)
   ) slave_r_buffer_i (
        .clk_i          ( ACLK       ),
        .rst_ni         ( ARESETn    ),
        .test_en_i      ( test_en_i  ),
        .slave_valid_i  ( RVALID     ),
        .slave_data_i   ( RDATA      ),
        .slave_resp_i   ( RRESP      ),
        .slave_user_i   ( RUSER      ),
        .slave_id_i     ( RID        ),
        .slave_last_i   ( RLAST      ),
        .slave_ready_o  ( RREADY     ),
        .master_valid_o ( RVALID_o   ),
        .master_data_o  ( RDATA_o    ),
        .master_resp_o  ( RRESP_o    ),
        .master_user_o  ( RUSER_o    ),
        .master_id_o    ( RID_o      ),
        .master_last_o  ( RLAST_o    ),
        .master_ready_i ( RREADY_i   )
   );
   axi_b_buffer #(
        .ID_WIDTH(AXI4_ID_WIDTH),
        .USER_WIDTH(AXI4_USER_WIDTH),
        .BUFFER_DEPTH(BUFF_DEPTH_SLAVE)
   ) slave_b_buffer_i (
        .clk_i          ( ACLK      ),
        .rst_ni         ( ARESETn   ),
        .test_en_i      ( test_en_i ),
        .slave_valid_i  ( BVALID    ),
        .slave_resp_i   ( BRESP     ),
        .slave_id_i     ( BID       ),
        .slave_user_i   ( BUSER     ),
        .slave_ready_o  ( BREADY    ),
        .master_valid_o ( BVALID_o  ),
        .master_resp_o  ( BRESP_o   ),
        .master_id_o    ( BID_o     ),
        .master_user_o  ( BUSER_o   ),
        .master_ready_i ( BREADY_i  )
   );
    
    always_ff @(posedge ACLK, negedge ARESETn) begin
        if (ARESETn == 1'b0)
            RR_FLAG <= 1'b0;
        else
            RR_FLAG <= ~RR_FLAG;
    end
    
    assign BE    = WSTRB;
    assign RDATA = Q;
    assign D     = WDATA;
    assign A   = address;
    assign WEN = (write_req) ? 1'b0 : 1'b1;
    always_comb begin
        CEN = ~(  write_req | read_req);
    end
    always_comb begin
        CountBurstNS   = CountBurstCS;
        AWREADY        = 1'b0;
        WREADY         = 1'b0;
        address        = '0;
        write_req      = 1'b0;
        sample_AW      = 1'b0;
        decr_AWLEN     = 1'b0;
        BID            = '0;
        BRESP          = 2'b00;
        BUSER          = '0;
        BVALID         = 1'b0;
        ARREADY        = 1'b0;
        read_req       = 1'b0;
        sample_AR      = 1'b0;
        decr_ARLEN     = 1'b0;
        RRESP          = 2'b00;
        RUSER          = '0;
        RLAST          = 1'b0;
        RID            = '0;
        
        address        = address_q;
        NS = CS;
        case (CS)
            IDLE: begin
                case (RR_FLAG)
                    1'b0: begin 
                        if (ARVALID == 1'b1) begin
                            sample_AR      = 1'b1;
                            read_req       = 1'b1;
                            address        = ARADDR;
                            ARREADY        = 1'b1;
                            if (ARLEN == 0) begin
                                NS = SINGLE_RD;
                                CountBurstNS   = '0;
                            end else  begin
                                NS           = (ARBURST == 2'b01) ? BURST_RD : WRAP_RD;
                                CountBurstNS = CountBurstCS + 1'b1;
                            end
                        end else begin
                            if (AWVALID) begin
                                AWREADY   = 1'b1;
                                sample_AW = 1'b1;
                                WREADY    = 1'b1;
                                if (WVALID) begin
                                    write_req = 1'b1;
                                    address   =  AWADDR;
                                    decr_AWLEN = 1'b1;
                                    if (AWLEN == 0) begin
                                          NS            = SINGLE_WR;
                                          CountBurstNS  = 0;
                                    end else begin
                                        NS            = (AWBURST == 2'b01) ? BURST_WR : WRAP_WR;
                                        CountBurstNS  = 1;
                                    end
                                end else begin 
                                    write_req  = 1'b0;
                                    address    = '0;
                                    if (AWLEN == 0) begin
                                        NS           =  WAIT_WDATA_SINGLE;
                                        CountBurstNS = 0;
                                    end else begin
                                        NS           =  (AWBURST == 2'b01) ? WAIT_WDATA_BURST : WAIT_WDATA_BURST_WRAP;
                                        CountBurstNS = 0;
                                    end
                                end
                            end else begin
                                NS = IDLE;
                            end
                        end
                    end
                    1'b1: begin
                        if (AWVALID) begin
                            AWREADY         = 1'b1;
                            sample_AW       = 1'b1;
                            WREADY          = 1'b1;
                            if (WVALID) begin
                                write_req       = 1'b1;
                                address         =  AWADDR;
                                decr_AWLEN      = 1'b1;
                                if (AWLEN == 0) begin
                                    NS              = SINGLE_WR;
                                    CountBurstNS    = 0;
                                end else begin
                                    NS              = (AWBURST == 2'b01) ? BURST_WR : WRAP_WR;
                                    CountBurstNS    = 1;
                                end
                            end else begin 
                                write_req  = 1'b0;
                                address    = '0;
                                if (AWLEN == 0) begin
                                    NS           =  WAIT_WDATA_SINGLE;
                                    CountBurstNS = 0;
                                end else begin
                                    NS           =  (AWBURST == 2'b01) ? WAIT_WDATA_BURST : WAIT_WDATA_BURST_WRAP;
                                    CountBurstNS = 0;
                                end
                            end
                        end else if (ARVALID) begin
                            sample_AR      = 1'b1;
                            read_req       = 1'b1;
                            address        = ARADDR;
                            ARREADY        = 1'b1;
                            if (ARLEN == 0) begin
                                NS = SINGLE_RD;
                                CountBurstNS   = '0;
                            end else begin
                                NS             = (ARBURST == 2'b01) ? BURST_RD : WRAP_RD;
                                CountBurstNS   = CountBurstCS + 1'b1;
                            end
                        end else begin
                            NS = IDLE;
                        end
                    end
                endcase
            end
            SINGLE_RD: begin
                RRESP  = 2'b00;
                RID    = ARID_Q;
                RUSER  = ARUSER_Q;
                RLAST  = 1'b1;
                
                if (RREADY) begin
                    NS             = IDLE;
                    CountBurstNS   = '0;
                end else begin
                    NS             = SINGLE_RD;
                    read_req       = 1'b1;
                    address        = ARADDR_Q;
                    CountBurstNS   = '0;
                end
            end
            BURST_RD, WRAP_RD:  begin
                automatic logic [AXI4_ADDRESS_WIDTH-1:0] aligned_address = ARADDR_Q & ~{{{AXI4_ADDRESS_WIDTH - 3}{1'b0}}, ar_size_q};
                automatic logic [AXI4_ADDRESS_WIDTH-1:0] wrap_boundary = aligned_address + (1 << ar_size_q) * (arlen_fixed_q + 1);
                automatic logic [AXI4_ADDRESS_WIDTH-1:0] addr = ARADDR_Q + (CountBurstCS << ADDRESS_BITS);
                RRESP   = 2'b00;
                RID     = ARID_Q;
                RUSER   = ARUSER_Q;
                ARREADY = 1'b0;
                if (RREADY) begin
                    if (ARLEN_Q > 0) begin
                        read_req      = 1'b1; 
                        decr_ARLEN    = 1'b1;
                        CountBurstNS  = CountBurstCS + 1'b1;
                        address = addr;
                        if (CS == WRAP_RD) begin
                            
                            if (addr == wrap_boundary)
                                CountBurstNS = 0;
                        end
                        RLAST         = 1'b0;
                    end else begin 
                        RLAST         = 1'b1;
                        NS            = IDLE;
                        CountBurstNS  = '0;
                    end
                end else begin 
                    read_req     = 1'b1; 
                    decr_ARLEN   = 1'b0;
                    ARREADY      = 1'b0;
                    address      = address_q;
                end
            end
            SINGLE_WR: begin
                BID          = AWID_Q;
                BRESP        = 2'b00;
                BUSER        = AWUSER_Q;
                BVALID       = 1'b1;
                AWREADY      = 1'b0;
                CountBurstNS = '0;
                if (BREADY)  begin
                    NS = IDLE;
                end else begin
                    NS = SINGLE_WR;
                end
            end
            BURST_WR, WRAP_WR: begin
                automatic logic [AXI4_ADDRESS_WIDTH-1:0] aligned_address = AWADDR_Q & ~{{{AXI4_ADDRESS_WIDTH - 3}{1'b0}}, aw_size_q};
                automatic logic [AXI4_ADDRESS_WIDTH-1:0] wrap_boundary = aligned_address + (1 << aw_size_q) * (awlen_fixed_q + 1);
                automatic logic [AXI4_ADDRESS_WIDTH-1:0] addr = AWADDR_Q + (CountBurstCS << ADDRESS_BITS);
                WREADY   = 1'b1;
                AWREADY  = 1'b0;
                address = addr;
                if (CS == WRAP_WR) begin
                    
                    if (addr == wrap_boundary)
                        CountBurstNS = 0;
                end
                if (WVALID) begin
                    write_req = 1'b1; 
                      if (AWLEN_Q > 0) begin
                          decr_AWLEN   = 1'b1;
                          CountBurstNS = CountBurstCS + 1'b1;
                      end else begin
                          decr_AWLEN   = 1'b0;
                          NS           = BURST_RESP;
                    end
                end else begin
                    write_req  = 1'b0; 
                    decr_AWLEN = 1'b0;
                end
            end
            BURST_RESP: begin
                BVALID       = 1'b1;
                BID          = AWID_Q;
                BRESP        = 2'b00;
                BUSER        = AWUSER_Q;
                AWREADY      = 1'b0;
                CountBurstNS = '0;
                if (BREADY) begin
                    NS = IDLE;
                end else begin 
                    NS = BURST_RESP;
                end
            end
            WAIT_WDATA_BURST, WAIT_WDATA_BURST_WRAP: begin
                AWREADY  = 1'b0;
                WREADY   = 1'b1;
                address  =  AWADDR_Q;
                if (WVALID) begin
                    write_req    = 1'b1;
                    NS           = (CS == WAIT_WDATA_BURST) ? BURST_WR : WRAP_WR;
                    CountBurstNS = 1;
                    decr_AWLEN   = 1'b1;
                end else begin
                    write_req    = 1'b0;
                    CountBurstNS = '0;
                end
            end
            WAIT_WDATA_SINGLE: begin
                AWREADY          = 1'b0;
                WREADY           = 1'b1;
                CountBurstNS     = '0;
                decr_AWLEN       =  1'b0;
                address          =  AWADDR_Q;
                if (WVALID) begin
                    write_req        =  1'b1;
                    NS               =  BURST_RESP;
                end else begin
                    NS = WAIT_WDATA_SINGLE; 
                end
            end
            default:
              NS = CS;
        endcase
    end
    
    always_ff @(posedge ACLK, negedge ARESETn) begin
        if (ARESETn == 1'b0) begin
            CS           <= IDLE;
            CountBurstCS <= '0;
            
            ARLEN_Q       <= '0;
            ARADDR_Q      <= '0;
            ARID_Q        <= '0;
            ARUSER_Q      <= '0;
            ar_size_q     <= '0;
            RVALID        <= 1'b0;
            
            AWADDR_Q      <= '0;
            AWID_Q        <= '0;
            AWUSER_Q      <= '0;
            AWLEN_Q       <= '0;
            arlen_fixed_q <= '0;
            awlen_fixed_q <= '0;
            aw_size_q     <= '0;
            address_q     <= '0;
        end else begin
            CS           <= NS;
            address_q    <= address;
            CountBurstCS <= CountBurstNS;
            RVALID       <= read_req;
            if (sample_AR) begin
                ARLEN_Q            <=  ARLEN;
                ARID_Q             <=  ARID;
                ARADDR_Q           <=  ARADDR;
                ARUSER_Q           <=  ARUSER;
                arlen_fixed_q      <=  ARLEN;
                ar_size_q          <=  ARSIZE;
            end else begin
                if (decr_ARLEN)
                  ARLEN_Q  <=  ARLEN_Q - 1'b1;
            end
            if (sample_AW) begin
                AWADDR_Q  <=  AWADDR;
                AWID_Q    <=  AWID;
                AWUSER_Q  <=  AWUSER;
                aw_size_q <= AWSIZE;
                awlen_fixed_q <= AWLEN;
            end
            case({sample_AW,decr_AWLEN})
              2'b00: AWLEN_Q  <=  AWLEN_Q;
              2'b01: AWLEN_Q  <=  AWLEN_Q - 1'b1;
              2'b10: AWLEN_Q  <=  AWLEN;
              2'b11: AWLEN_Q  <=  AWLEN   - 1'b1;
            endcase
          end
        end
endmodule
module   axi_mem_if_var_latency
#(
    parameter AXI4_ADDRESS_WIDTH = 32,
    parameter AXI4_RDATA_WIDTH   = 64,
    parameter AXI4_WDATA_WIDTH   = 64,
    parameter AXI4_ID_WIDTH      = 16,
    parameter AXI4_USER_WIDTH    = 10,
    parameter AXI_NUMBYTES       = AXI4_WDATA_WIDTH/8,
    parameter MEM_ADDR_WIDTH     = 13,
    parameter BUFF_DEPTH_SLAVE   = 4,
    parameter LATENCY_AW         = 50,
    parameter LATENCY_AR         = 50,
    parameter LATENCY_R          = 50,
    parameter LATENCY_B          = 50,
    parameter LATENCY_W          = 50
)
(
    input logic                                     ACLK,
    input logic                                     ARESETn,
    
    
    
    
    input  logic [AXI4_ID_WIDTH-1:0]                AWID_i     ,
    input  logic [AXI4_ADDRESS_WIDTH-1:0]           AWADDR_i   ,
    input  logic [ 7:0]                             AWLEN_i    ,
    input  logic [ 2:0]                             AWSIZE_i   ,
    input  logic [ 1:0]                             AWBURST_i  ,
    input  logic                                    AWLOCK_i   ,
    input  logic [ 3:0]                             AWCACHE_i  ,
    input  logic [ 2:0]                             AWPROT_i   ,
    input  logic [ 3:0]                             AWREGION_i ,
    input  logic [ AXI4_USER_WIDTH-1:0]             AWUSER_i   ,
    input  logic [ 3:0]                             AWQOS_i    ,
    input  logic                                    AWVALID_i  ,
    output logic                                    AWREADY_o  ,
    
    
    input  logic [AXI_NUMBYTES-1:0][7:0]            WDATA_i    ,
    input  logic [AXI_NUMBYTES-1:0]                 WSTRB_i    ,
    input  logic                                    WLAST_i    ,
    input  logic [AXI4_USER_WIDTH-1:0]              WUSER_i    ,
    input  logic                                    WVALID_i   ,
    output logic                                    WREADY_o   ,
    
    
    output logic   [AXI4_ID_WIDTH-1:0]              BID_o      ,
    output logic   [ 1:0]                           BRESP_o    ,
    output logic                                    BVALID_o   ,
    output logic   [AXI4_USER_WIDTH-1:0]            BUSER_o    ,
    input  logic                                    BREADY_i   ,
    
    
    input  logic [AXI4_ID_WIDTH-1:0]                ARID_i     ,
    input  logic [AXI4_ADDRESS_WIDTH-1:0]           ARADDR_i   ,
    input  logic [ 7:0]                             ARLEN_i    ,
    input  logic [ 2:0]                             ARSIZE_i   ,
    input  logic [ 1:0]                             ARBURST_i  ,
    input  logic                                    ARLOCK_i   ,
    input  logic [ 3:0]                             ARCACHE_i  ,
    input  logic [ 2:0]                             ARPROT_i   ,
    input  logic [ 3:0]                             ARREGION_i ,
    input  logic [ AXI4_USER_WIDTH-1:0]             ARUSER_i   ,
    input  logic [ 3:0]                             ARQOS_i    ,
    input  logic                                    ARVALID_i  ,
    output logic                                    ARREADY_o  ,
    
    
    output  logic [AXI4_ID_WIDTH-1:0]               RID_o      ,
    output  logic [AXI4_RDATA_WIDTH-1:0]            RDATA_o    ,
    output  logic [ 1:0]                            RRESP_o    ,
    output  logic                                   RLAST_o    ,
    output  logic [AXI4_USER_WIDTH-1:0]             RUSER_o    ,
    output  logic                                   RVALID_o   ,
    input   logic                                   RREADY_i   ,
    
    output logic                                    CEN        ,
    output logic                                    WEN        ,
    output logic  [MEM_ADDR_WIDTH-1:0]              A          ,
    output logic  [AXI4_WDATA_WIDTH-1:0]            D          ,
    output logic  [AXI_NUMBYTES-1:0]                BE         ,
    input  logic  [AXI4_RDATA_WIDTH-1:0]            Q
);
  
  
  
  
  logic [LATENCY_AW-1:0][AXI4_ID_WIDTH-1:0]             AWID       ;
  logic [LATENCY_AW-1:0][AXI4_ADDRESS_WIDTH-1:0]        AWADDR     ;
  logic [LATENCY_AW-1:0][ 7:0]                          AWLEN      ;
  logic [LATENCY_AW-1:0][ 2:0]                          AWSIZE     ;
  logic [LATENCY_AW-1:0][ 1:0]                          AWBURST    ;
  logic [LATENCY_AW-1:0]                                AWLOCK     ;
  logic [LATENCY_AW-1:0][ 3:0]                          AWCACHE    ;
  logic [LATENCY_AW-1:0][ 2:0]                          AWPROT     ;
  logic [LATENCY_AW-1:0][ 3:0]                          AWREGION   ;
  logic [LATENCY_AW-1:0][ AXI4_USER_WIDTH-1:0]          AWUSER     ;
  logic [LATENCY_AW-1:0][ 3:0]                          AWQOS      ;
  logic [LATENCY_AW-1:0]                                AWVALID    ;
  logic                                                 AWREADY    ;
  logic                                                 AWREADY_int;
  
  
  logic [LATENCY_W-1:0][AXI_NUMBYTES-1:0][7:0]          WDATA      ;
  logic [LATENCY_W-1:0][AXI_NUMBYTES-1:0]               WSTRB      ;
  logic [LATENCY_W-1:0]                                 WLAST      ;
  logic [LATENCY_W-1:0][AXI4_USER_WIDTH-1:0]            WUSER      ;
  logic [LATENCY_W-1:0]                                 WVALID     ;
  logic                                                 WREADY     ;
  logic                                                 WREADY_int ;
  
  
  logic [LATENCY_B-1:0][AXI4_ID_WIDTH-1:0]             BID         ;
  logic [LATENCY_B-1:0][ 1:0]                          BRESP       ;
  logic [LATENCY_B-1:0]                                BVALID      ;
  logic [LATENCY_B-1:0] [AXI4_USER_WIDTH-1:0]          BUSER       ;
  logic                                                BREADY      ;
  logic [AXI4_ID_WIDTH-1:0]                            BID_int     ;
  logic [ 1:0]                                         BRESP_int   ;
  logic                                                BVALID_int  ;
  logic [AXI4_USER_WIDTH-1:0]                          BUSER_int   ;
  
  
  logic [LATENCY_AR-1:0][AXI4_ID_WIDTH-1:0]            ARID       ;
  logic [LATENCY_AR-1:0][AXI4_ADDRESS_WIDTH-1:0]       ARADDR     ;
  logic [LATENCY_AR-1:0][ 7:0]                         ARLEN      ;
  logic [LATENCY_AR-1:0][ 2:0]                         ARSIZE     ;
  logic [LATENCY_AR-1:0][ 1:0]                         ARBURST    ;
  logic [LATENCY_AR-1:0]                               ARLOCK     ;
  logic [LATENCY_AR-1:0][ 3:0]                         ARCACHE    ;
  logic [LATENCY_AR-1:0][ 2:0]                         ARPROT     ;
  logic [LATENCY_AR-1:0][ 3:0]                         ARREGION   ;
  logic [LATENCY_AR-1:0][ AXI4_USER_WIDTH-1:0]         ARUSER     ;
  logic [LATENCY_AR-1:0][ 3:0]                         ARQOS      ;
  logic [LATENCY_AR-1:0]                               ARVALID    ;
  logic                                                ARREADY    ;
  logic                                                ARREADY_int;
  
  
  logic [LATENCY_R-1:0][AXI4_ID_WIDTH-1:0]             RID        ;
  logic [LATENCY_R-1:0][AXI4_RDATA_WIDTH-1:0]          RDATA      ;
  logic [LATENCY_R-1:0][ 1:0]                          RRESP      ;
  logic [LATENCY_R-1:0]                                RLAST      ;
  logic [LATENCY_R-1:0][AXI4_USER_WIDTH-1:0]           RUSER      ;
  logic [LATENCY_R-1:0]                                RVALID     ;
  logic                                                RREADY     ;
  logic [AXI4_ID_WIDTH-1:0]                            RID_int    ;
  logic [AXI4_RDATA_WIDTH-1:0]                         RDATA_int  ;
  logic [ 1:0]                                         RRESP_int  ;
  logic                                                RLAST_int  ;
  logic [AXI4_USER_WIDTH-1:0]                          RUSER_int  ;
  logic                                                RVALID_int ;
  
  
  
  int unsigned i,j,k,l,m;
    always_ff @(posedge ACLK, negedge ARESETn)
    begin
      if(ARESETn == 1'b0)
      begin
           for(i=0;i<LATENCY_AW;i++)
           begin
              AWID[i]    <= '0;
              AWADDR[i]  <= '0;
              AWLEN[i]   <= '0;
              AWSIZE[i]  <= '0;
              AWBURST[i] <= '0;
              AWLOCK[i]  <= '0;
              AWCACHE[i] <= '0;
              AWPROT[i]  <= '0;
              AWREGION[i]<= '0;
              AWUSER[i]  <= '0;
              AWQOS[i]   <= '0;
              AWVALID[i] <= '0;
           end
      end
      else
      begin
           if(AWREADY)
           begin
              AWID[0]    <=   AWID_i    ;
              AWADDR[0]  <=   AWADDR_i  ;
              AWLEN[0]   <=   AWLEN_i   ;
              AWSIZE[0]  <=   AWSIZE_i  ;
              AWBURST[0] <=   AWBURST_i ;
              AWLOCK[0]  <=   AWLOCK_i  ;
              AWCACHE[0] <=   AWCACHE_i ;
              AWPROT[0]  <=   AWPROT_i  ;
              AWREGION[0]<=   AWREGION_i;
              AWUSER[0]  <=   AWUSER_i  ;
              AWQOS[0]   <=   AWQOS_i   ;
              AWVALID[0] <=   AWVALID_i ;
              AWID[LATENCY_AW-1:1]    <=   AWID[LATENCY_AW-2:0]    ;
              AWADDR[LATENCY_AW-1:1]  <=   AWADDR[LATENCY_AW-2:0]  ;
              AWLEN[LATENCY_AW-1:1]   <=   AWLEN[LATENCY_AW-2:0]   ;
              AWSIZE[LATENCY_AW-1:1]  <=   AWSIZE[LATENCY_AW-2:0]  ;
              AWBURST[LATENCY_AW-1:1] <=   AWBURST[LATENCY_AW-2:0] ;
              AWLOCK[LATENCY_AW-1:1]  <=   AWLOCK[LATENCY_AW-2:0]  ;
              AWCACHE[LATENCY_AW-1:1] <=   AWCACHE[LATENCY_AW-2:0] ;
              AWPROT[LATENCY_AW-1:1]  <=   AWPROT[LATENCY_AW-2:0]  ;
              AWREGION[LATENCY_AW-1:1]<=   AWREGION[LATENCY_AW-2:0];
              AWUSER[LATENCY_AW-1:1]  <=   AWUSER[LATENCY_AW-2:0]  ;
              AWQOS[LATENCY_AW-1:1]   <=   AWQOS[LATENCY_AW-2:0]   ;
              AWVALID[LATENCY_AW-1:1] <=   AWVALID[LATENCY_AW-2:0] ;
           end
      end
    end
    always_ff @(posedge ACLK, negedge ARESETn)
    begin
      if(ARESETn == 1'b0)
      begin
           for(j=0;j<LATENCY_AR;j++)
           begin
              ARID[j]    <= '0;
              ARADDR[j]  <= '0;
              ARLEN[j]   <= '0;
              ARSIZE[j]  <= '0;
              ARBURST[j] <= '0;
              ARLOCK[j]  <= '0;
              ARCACHE[j] <= '0;
              ARPROT[j]  <= '0;
              ARREGION[j]<= '0;
              ARUSER[j]  <= '0;
              ARQOS[j]   <= '0;
              ARVALID[j] <= '0;
           end
      end
      else
      begin
           if(ARREADY)
           begin
              ARID[0]    <=   ARID_i    ;
              ARADDR[0]  <=   ARADDR_i  ;
              ARLEN[0]   <=   ARLEN_i   ;
              ARSIZE[0]  <=   ARSIZE_i  ;
              ARBURST[0] <=   ARBURST_i ;
              ARLOCK[0]  <=   ARLOCK_i  ;
              ARCACHE[0] <=   ARCACHE_i ;
              ARPROT[0]  <=   ARPROT_i  ;
              ARREGION[0]<=   ARREGION_i;
              ARUSER[0]  <=   ARUSER_i  ;
              ARQOS[0]   <=   ARQOS_i   ;
              ARVALID[0] <=   ARVALID_i ;
              ARID[LATENCY_AR-1:1]    <=   ARID[LATENCY_AR-2:0]    ;
              ARADDR[LATENCY_AR-1:1]  <=   ARADDR[LATENCY_AR-2:0]  ;
              ARLEN[LATENCY_AR-1:1]   <=   ARLEN[LATENCY_AR-2:0]   ;
              ARSIZE[LATENCY_AR-1:1]  <=   ARSIZE[LATENCY_AR-2:0]  ;
              ARBURST[LATENCY_AR-1:1] <=   ARBURST[LATENCY_AR-2:0] ;
              ARLOCK[LATENCY_AR-1:1]  <=   ARLOCK[LATENCY_AR-2:0]  ;
              ARCACHE[LATENCY_AR-1:1] <=   ARCACHE[LATENCY_AR-2:0] ;
              ARPROT[LATENCY_AR-1:1]  <=   ARPROT[LATENCY_AR-2:0]  ;
              ARREGION[LATENCY_AR-1:1]<=   ARREGION[LATENCY_AR-2:0];
              ARUSER[LATENCY_AR-1:1]  <=   ARUSER[LATENCY_AR-2:0]  ;
              ARQOS[LATENCY_AR-1:1]   <=   ARQOS[LATENCY_AR-2:0]   ;
              ARVALID[LATENCY_AR-1:1] <=   ARVALID[LATENCY_AR-2:0] ;
           end
      end
    end
    assign RID_o    = RID   [LATENCY_R-1];
    assign RDATA_o  = RDATA [LATENCY_R-1];
    assign RRESP_o  = RRESP [LATENCY_R-1];
    assign RLAST_o  = RLAST [LATENCY_R-1];
    assign RUSER_o  = RUSER [LATENCY_R-1];
    assign RVALID_o = RVALID[LATENCY_R-1];
    
    always_ff @(posedge ACLK, negedge ARESETn)
    begin
      if(ARESETn == 1'b0)
      begin
           for(k=0;k<LATENCY_R;k++)
           begin
              RID[k]    <= '0;
              RDATA[k]  <= '0;
              RRESP[k]  <= '0;
              RLAST[k]  <= '0;
              RUSER[k]  <= '0;
              RVALID[k] <= '0;
           end
      end
      else
      begin
           if(RREADY)
           begin
              RID[0]    <= RID_int    ;
              RDATA[0]  <= RDATA_int  ;
              RRESP[0]  <= RRESP_int  ;
              RLAST[0]  <= RLAST_int  ;
              RUSER[0]  <= RUSER_int  ;
              RVALID[0] <= RVALID_int ;
              RID[LATENCY_R-1:1]      <= RID[LATENCY_R-2:0]   ;
              RDATA[LATENCY_R-1:1]    <= RDATA[LATENCY_R-2:0] ;
              RRESP[LATENCY_R-1:1]    <= RRESP[LATENCY_R-2:0] ;
              RLAST[LATENCY_R-1:1]    <= RLAST[LATENCY_R-2:0] ;
              RUSER[LATENCY_R-1:1]    <= RUSER[LATENCY_R-2:0] ;
              RVALID[LATENCY_R-1:1]   <= RVALID[LATENCY_R-2:0];
           end
      end
    end
    assign BID_o    = BID   [LATENCY_B-1];
    assign BRESP_o  = BRESP [LATENCY_B-1];
    assign BUSER_o  = BUSER [LATENCY_B-1];
    assign BVALID_o = BVALID[LATENCY_B-1];
    
    always_ff @(posedge ACLK, negedge ARESETn)
    begin
      if(ARESETn == 1'b0)
      begin
           for(l=0;l<LATENCY_B;l++)
           begin
              BID[l]    <= '0;
              BRESP[l]  <= '0;
              BUSER[l]  <= '0;
              BVALID[l] <= '0;
           end
      end
      else
      begin
           if(BREADY)
           begin
              BID[0]    <=  BID_int;
              BRESP[0]  <=  BRESP_int;
              BUSER[0]  <=  BUSER_int;
              BVALID[0] <=  BVALID_int;
              BID[LATENCY_B-1:1]      <= BID[LATENCY_B-2:0]   ;
              BRESP[LATENCY_B-1:1]    <= BRESP[LATENCY_B-2:0] ;
              BUSER[LATENCY_B-1:1]    <= BUSER[LATENCY_B-2:0] ;
              BVALID[LATENCY_B-1:1]   <= BVALID[LATENCY_B-2:0];
           end
      end
    end
    
    
    always_ff @(posedge ACLK, negedge ARESETn)
    begin
      if(ARESETn == 1'b0)
      begin
           for(m=0;m<LATENCY_W;m++)
           begin
              WDATA[m]   <= '0;
              WSTRB[m]   <= '0;
              WLAST[m]   <= '0;
              WUSER[m]   <= '0;
              WVALID[m]  <= '0;
           end
      end
      else
      begin
           if(WREADY)
           begin
              WDATA[0]   <= WDATA_i ;
              WSTRB[0]   <= WSTRB_i ;
              WLAST[0]   <= WLAST_i ;
              WUSER[0]   <= WUSER_i ;
              WVALID[0]  <= WVALID_i;
              WDATA [LATENCY_W-1:1]  <= WDATA [LATENCY_W-2:0];
              WSTRB [LATENCY_W-1:1]  <= WSTRB [LATENCY_W-2:0];
              WLAST [LATENCY_W-1:1]  <= WLAST [LATENCY_W-2:0];
              WUSER [LATENCY_W-1:1]  <= WUSER [LATENCY_W-2:0];
              WVALID[LATENCY_W-1:1]  <= WVALID[LATENCY_W-2:0];
           end
      end
    end
    assign  AWREADY    =   AWREADY_int | ~AWVALID[LATENCY_AW-1];
    assign  ARREADY    =   ARREADY_int | ~ARVALID[LATENCY_AR-1];
    assign  WREADY     =   WREADY_int  | ~WVALID[LATENCY_W-1];
    assign  AWREADY_o =   AWREADY;
    assign  ARREADY_o =   ARREADY;
    assign  RREADY    =   RREADY_i | ~RVALID[LATENCY_R-1];
    assign  BREADY    =   BREADY_i | ~BVALID[LATENCY_B-1];
    assign  WREADY_o  =   WREADY;
    axi_mem_if
    #(
        .AXI4_ADDRESS_WIDTH(AXI4_ADDRESS_WIDTH),
        .AXI4_RDATA_WIDTH(AXI4_RDATA_WIDTH),
        .AXI4_WDATA_WIDTH(AXI4_WDATA_WIDTH),
        .AXI4_ID_WIDTH(AXI4_ID_WIDTH),
        .AXI4_USER_WIDTH(AXI4_USER_WIDTH),
        .MEM_ADDR_WIDTH(MEM_ADDR_WIDTH),
        .BUFF_DEPTH_SLAVE(BUFF_DEPTH_SLAVE)
    )
    axi_mem_if_i
    (
        .ACLK(ACLK),
        .ARESETn(ARESETn),
        .AWVALID_i  ( AWVALID[LATENCY_AW-1]  ),
        .AWADDR_i   ( AWADDR[LATENCY_AW-1]   ),
        .AWPROT_i   ( AWPROT[LATENCY_AW-1]   ),
        .AWREGION_i ( AWREGION[LATENCY_AW-1] ),
        .AWLEN_i    ( AWLEN[LATENCY_AW-1]    ),
        .AWSIZE_i   ( AWSIZE[LATENCY_AW-1]   ),
        .AWBURST_i  ( AWBURST[LATENCY_AW-1]  ),
        .AWLOCK_i   ( AWLOCK[LATENCY_AW-1]   ),
        .AWCACHE_i  ( AWCACHE[LATENCY_AW-1]  ),
        .AWQOS_i    ( AWQOS[LATENCY_AW-1]    ),
        .AWID_i     ( AWID[LATENCY_AW-1]     ),
        .AWUSER_i   ( AWUSER[LATENCY_AW-1]   ),
        .AWREADY_o  ( AWREADY_int            ),
        .ARVALID_i  ( ARVALID[LATENCY_AR-1]  ),
        .ARADDR_i   ( ARADDR[LATENCY_AR-1]   ),
        .ARPROT_i   ( ARPROT[LATENCY_AR-1]   ),
        .ARREGION_i ( ARREGION[LATENCY_AR-1] ),
        .ARLEN_i    ( ARLEN[LATENCY_AR-1]    ),
        .ARSIZE_i   ( ARSIZE[LATENCY_AR-1]   ),
        .ARBURST_i  ( ARBURST[LATENCY_AR-1]  ),
        .ARLOCK_i   ( ARLOCK[LATENCY_AR-1]   ),
        .ARCACHE_i  ( ARCACHE[LATENCY_AR-1]  ),
        .ARQOS_i    ( ARQOS[LATENCY_AR-1]    ),
        .ARID_i     ( ARID[LATENCY_AR-1]     ),
        .ARUSER_i   ( ARUSER[LATENCY_AR-1]   ),
        .ARREADY_o  ( ARREADY_int            ),
        .RVALID_o   ( RVALID_int             ),
        .RDATA_o    ( RDATA_int              ),
        .RRESP_o    ( RRESP_int              ),
        .RLAST_o    ( RLAST_int              ),
        .RID_o      ( RID_int                ),
        .RUSER_o    ( RUSER_int              ),
        .RREADY_i   ( RREADY                 ),
        .WVALID_i   ( WVALID[LATENCY_W-1]    ),
        .WDATA_i    ( WDATA[LATENCY_W-1]     ),
        .WSTRB_i    ( WSTRB[LATENCY_W-1]     ),
        .WLAST_i    ( WLAST[LATENCY_W-1]     ),
        .WUSER_i    ( WUSER[LATENCY_W-1]     ),
        .WREADY_o   ( WREADY_int             ),
        .BVALID_o  ( BVALID_int              ),
        .BRESP_o   ( BRESP_int               ),
        .BID_o     ( BID_int                 ),
        .BUSER_o   ( BUSER_int               ),
        .BREADY_i  ( BREADY                  ),
        .CEN       ( CEN                     ),
        .WEN       ( WEN                     ),
        .A         ( A                       ),
        .D         ( D                       ),
        .BE        ( BE                      ),
        .Q         ( Q                       )
    );
 endmodule
module axi_mem_if_wrap #(
    parameter AXI4_ADDRESS_WIDTH = 64,
    parameter AXI4_RDATA_WIDTH   = 64,
    parameter AXI4_WDATA_WIDTH   = 64,
    parameter AXI4_ID_WIDTH      = 16,
    parameter AXI4_USER_WIDTH    = 10,
    parameter AXI_NUMBYTES       = AXI4_WDATA_WIDTH/8,
    parameter BUFF_DEPTH_SLAVE   = 4
)(
    input logic                            clk_i,          
    input logic                            rst_ni,         
    input logic                            test_en_i,
    AXI_BUS.Slave                          slave,
    output logic                           CEN,
    output logic                           WEN,
    output logic  [AXI4_ADDRESS_WIDTH-1:0] A,
    output logic  [AXI4_WDATA_WIDTH-1:0]   D,
    output logic  [AXI_NUMBYTES-1:0]       BE,
    input  logic  [AXI4_RDATA_WIDTH-1:0]   Q
);
    axi_mem_if #(
        .AXI4_ADDRESS_WIDTH ( AXI4_ADDRESS_WIDTH ),
        .AXI4_RDATA_WIDTH   ( AXI4_RDATA_WIDTH   ),
        .AXI4_WDATA_WIDTH   ( AXI4_WDATA_WIDTH   ),
        .AXI4_ID_WIDTH      ( AXI4_ID_WIDTH      ),
        .AXI4_USER_WIDTH    ( AXI4_USER_WIDTH    ),
        .AXI_NUMBYTES       ( AXI_NUMBYTES       ),
        .BUFF_DEPTH_SLAVE   ( BUFF_DEPTH_SLAVE   )
    ) axi_mem_if_i (
        .ACLK       (  clk_i            ),
        .test_en_i  (  test_en_i        ),
        .ARESETn    (  rst_ni           ),
        .AWID_i     (  slave.aw_id      ),
        .AWADDR_i   (  slave.aw_addr    ),
        .AWLEN_i    (  slave.aw_len     ),
        .AWSIZE_i   (  slave.aw_size    ),
        .AWBURST_i  (  slave.aw_burst   ),
        .AWLOCK_i   (  slave.aw_lock    ),
        .AWCACHE_i  (  slave.aw_cache   ),
        .AWPROT_i   (  slave.aw_prot    ),
        .AWREGION_i (  slave.aw_region  ),
        .AWUSER_i   (  slave.aw_user    ),
        .AWQOS_i    (  slave.aw_qos     ),
        .AWVALID_i  (  slave.aw_valid   ),
        .AWREADY_o  (  slave.aw_ready   ),
        .WDATA_i    (  slave.w_data     ),
        .WSTRB_i    (  slave.w_strb     ),
        .WLAST_i    (  slave.w_last     ),
        .WUSER_i    (  slave.w_user     ),
        .WVALID_i   (  slave.w_valid    ),
        .WREADY_o   (  slave.w_ready    ),
        .BID_o      (  slave.b_id       ),
        .BRESP_o    (  slave.b_resp     ),
        .BVALID_o   (  slave.b_valid    ),
        .BUSER_o    (  slave.b_user     ),
        .BREADY_i   (  slave.b_ready    ),
        .ARID_i     (  slave.ar_id      ),
        .ARADDR_i   (  slave.ar_addr    ),
        .ARLEN_i    (  slave.ar_len     ),
        .ARSIZE_i   (  slave.ar_size    ),
        .ARBURST_i  (  slave.ar_burst   ),
        .ARLOCK_i   (  slave.ar_lock    ),
        .ARCACHE_i  (  slave.ar_cache   ),
        .ARPROT_i   (  slave.ar_prot    ),
        .ARREGION_i (  slave.ar_region  ),
        .ARUSER_i   (  slave.ar_user    ),
        .ARQOS_i    (  slave.ar_qos     ),
        .ARVALID_i  (  slave.ar_valid   ),
        .ARREADY_o  (  slave.ar_ready   ),
        .RID_o      (  slave.r_id       ),
        .RDATA_o    (  slave.r_data     ),
        .RRESP_o    (  slave.r_resp     ),
        .RLAST_o    (  slave.r_last     ),
        .RUSER_o    (  slave.r_user     ),
        .RVALID_o   (  slave.r_valid    ),
        .RREADY_i   (  slave.r_ready    ),
        .*
    );
endmodule
package riscv;
    
    
    
    typedef enum logic [3:0] {
       ModeOff  = 0,
       ModeSv32 = 1,
       ModeSv39 = 8,
       ModeSv48 = 9,
       ModeSv57 = 10,
       ModeSv64 = 11
    } vm_mode_t;
    localparam XLEN = 64;
    
    
    localparam VLEN       = (XLEN == 32) ? 32 : 64;    
    localparam PLEN       = (XLEN == 32) ? 34 : 56;    
    localparam IS_XLEN32  = (XLEN == 32) ? 1'b1 : 1'b0;
    localparam IS_XLEN64  = (XLEN == 32) ? 1'b0 : 1'b1;
    localparam ModeW      = (XLEN == 32) ? 1 : 4;
    localparam ASIDW      = (XLEN == 32) ? 9 : 16;
    localparam PPNW       = (XLEN == 32) ? 22 : 44;
    localparam vm_mode_t MODE_SV = (XLEN == 32) ? ModeSv32 : ModeSv39;
    localparam SV         = (MODE_SV == ModeSv32) ? 32 : 39;
    localparam VPN2       = (VLEN-31 < 8) ? VLEN-31 : 8;
    localparam  FPU_EN     = 1'b1; 
  
    typedef logic [XLEN-1:0] xlen_t;
    
    
    
    typedef enum logic[1:0] {
      PRIV_LVL_M = 2'b11,
      PRIV_LVL_S = 2'b01,
      PRIV_LVL_U = 2'b00
    } priv_lvl_t;
    
    typedef enum logic [1:0] {
        XLEN_32  = 2'b01,
        XLEN_64  = 2'b10,
        XLEN_128 = 2'b11
    } xlen_e;
    typedef enum logic [1:0] {
        Off     = 2'b00,
        Initial = 2'b01,
        Clean   = 2'b10,
        Dirty   = 2'b11
    } xs_t;
    typedef struct packed {
        logic         sd;     
        logic [62:36] wpri4;  
        xlen_e        sxl;    
        xlen_e        uxl;    
        logic [8:0]   wpri3;  
        logic         tsr;    
        logic         tw;     
        logic         tvm;    
        logic         mxr;    
        logic         sum;    
        logic         mprv;   
        xs_t          xs;     
        xs_t          fs;     
        priv_lvl_t    mpp;    
        logic [1:0]   wpri2;  
        logic         spp;    
        logic         mpie;   
        logic         wpri1;  
        logic         spie;   
        logic         upie;   
        logic         mie;    
        logic         wpri0;  
        logic         sie;    
        logic         uie;    
    } status_rv_t;
    typedef struct packed {
        logic [ModeW-1:0] mode;
        logic [ASIDW-1:0] asid;
        logic [PPNW-1:0]  ppn;
    } satp_t;
    
    
    
    typedef struct packed {
        logic [31:25] funct7;
        logic [24:20] rs2;
        logic [19:15] rs1;
        logic [14:12] funct3;
        logic [11:7]  rd;
        logic [6:0]   opcode;
    } rtype_t;
    typedef struct packed {
        logic [31:27] rs3;
        logic [26:25] funct2;
        logic [24:20] rs2;
        logic [19:15] rs1;
        logic [14:12] funct3;
        logic [11:7]  rd;
        logic [6:0]   opcode;
    } r4type_t;
    typedef struct packed {
        logic [31:27] funct5;
        logic [26:25] fmt;
        logic [24:20] rs2;
        logic [19:15] rs1;
        logic [14:12] rm;
        logic [11:7]  rd;
        logic [6:0]   opcode;
    } rftype_t; 
    typedef struct packed {
        logic [31:30] funct2;
        logic [29:25] vecfltop;
        logic [24:20] rs2;
        logic [19:15] rs1;
        logic [14:14] repl;
        logic [13:12] vfmt;
        logic [11:7]  rd;
        logic [6:0]   opcode;
    } rvftype_t; 
    typedef struct packed {
        logic [31:20] imm;
        logic [19:15] rs1;
        logic [14:12] funct3;
        logic [11:7]  rd;
        logic [6:0]   opcode;
    } itype_t;
    typedef struct packed {
        logic [31:25] imm;
        logic [24:20] rs2;
        logic [19:15] rs1;
        logic [14:12] funct3;
        logic [11:7]  imm0;
        logic [6:0]   opcode;
    } stype_t;
    typedef struct packed {
        logic [31:12] funct3;
        logic [11:7]  rd;
        logic [6:0]   opcode;
    } utype_t;
    
    typedef struct packed {
        logic [31:27] funct5;
        logic         aq;
        logic         rl;
        logic [24:20] rs2;
        logic [19:15] rs1;
        logic [14:12] funct3;
        logic [11:7]  rd;
        logic [6:0]   opcode;
    } atype_t;
    typedef union packed {
        logic [31:0]   instr;
        rtype_t        rtype;
        r4type_t       r4type;
        rftype_t       rftype;
        rvftype_t      rvftype;
        itype_t        itype;
        stype_t        stype;
        utype_t        utype;
        atype_t        atype;
    } instruction_t;
    
    
    
    
    
    localparam OpcodeLoad      = 7'b00_000_11;
    localparam OpcodeLoadFp    = 7'b00_001_11;
    localparam OpcodeCustom0   = 7'b00_010_11;
    localparam OpcodeMiscMem   = 7'b00_011_11;
    localparam OpcodeOpImm     = 7'b00_100_11;
    localparam OpcodeAuipc     = 7'b00_101_11;
    localparam OpcodeOpImm32   = 7'b00_110_11;
    
    localparam OpcodeStore     = 7'b01_000_11;
    localparam OpcodeStoreFp   = 7'b01_001_11;
    localparam OpcodeCustom1   = 7'b01_010_11;
    localparam OpcodeAmo       = 7'b01_011_11;
    localparam OpcodeOp        = 7'b01_100_11;
    localparam OpcodeLui       = 7'b01_101_11;
    localparam OpcodeOp32      = 7'b01_110_11;
    
    localparam OpcodeMadd      = 7'b10_000_11;
    localparam OpcodeMsub      = 7'b10_001_11;
    localparam OpcodeNmsub     = 7'b10_010_11;
    localparam OpcodeNmadd     = 7'b10_011_11;
    localparam OpcodeOpFp      = 7'b10_100_11;
    localparam OpcodeRsrvd1    = 7'b10_101_11;
    localparam OpcodeCustom2   = 7'b10_110_11;
    
    localparam OpcodeBranch    = 7'b11_000_11;
    localparam OpcodeJalr      = 7'b11_001_11;
    localparam OpcodeRsrvd2    = 7'b11_010_11;
    localparam OpcodeJal       = 7'b11_011_11;
    localparam OpcodeSystem    = 7'b11_100_11;
    localparam OpcodeRsrvd3    = 7'b11_101_11;
    localparam OpcodeCustom3   = 7'b11_110_11;
    
    
    localparam OpcodeC0             = 2'b00;
    localparam OpcodeC0Addi4spn     = 3'b000;
    localparam OpcodeC0Fld          = 3'b001;
    localparam OpcodeC0Lw           = 3'b010;
    localparam OpcodeC0Ld           = 3'b011;
    localparam OpcodeC0Rsrvd        = 3'b100;
    localparam OpcodeC0Fsd          = 3'b101;
    localparam OpcodeC0Sw           = 3'b110;
    localparam OpcodeC0Sd           = 3'b111;
    
    localparam OpcodeC1             = 2'b01;
    localparam OpcodeC1Addi         = 3'b000;
    localparam OpcodeC1Addiw        = 3'b001; 
    localparam OpcodeC1Jal          = 3'b001; 
    localparam OpcodeC1Li           = 3'b010;
    localparam OpcodeC1LuiAddi16sp  = 3'b011;
    localparam OpcodeC1MiscAlu      = 3'b100;
    localparam OpcodeC1J            = 3'b101;
    localparam OpcodeC1Beqz         = 3'b110;
    localparam OpcodeC1Bnez         = 3'b111;
    
    localparam OpcodeC2             = 2'b10;
    localparam OpcodeC2Slli         = 3'b000;
    localparam OpcodeC2Fldsp        = 3'b001;
    localparam OpcodeC2Lwsp         = 3'b010;
    localparam OpcodeC2Ldsp         = 3'b011;
    localparam OpcodeC2JalrMvAdd    = 3'b100;
    localparam OpcodeC2Fsdsp        = 3'b101;
    localparam OpcodeC2Swsp         = 3'b110;
    localparam OpcodeC2Sdsp         = 3'b111;
    
    
    
    
    typedef struct packed {
        logic [9:0]  reserved;
        logic [44-1:0] ppn; 
        logic [1:0]  rsw;
        logic d;
        logic a;
        logic g;
        logic u;
        logic x;
        logic w;
        logic r;
        logic v;
    } pte_t;
    
    typedef struct packed {
        logic [22-1:0] ppn; 
        logic [1:0]  rsw;
        logic d;
        logic a;
        logic g;
        logic u;
        logic x;
        logic w;
        logic r;
        logic v;
    } pte_sv32_t;
    
    
    
    localparam logic [XLEN-1:0] INSTR_ADDR_MISALIGNED = 0;
    localparam logic [XLEN-1:0] INSTR_ACCESS_FAULT    = 1;  
    localparam logic [XLEN-1:0] ILLEGAL_INSTR         = 2;
    localparam logic [XLEN-1:0] BREAKPOINT            = 3;
    localparam logic [XLEN-1:0] LD_ADDR_MISALIGNED    = 4;
    localparam logic [XLEN-1:0] LD_ACCESS_FAULT       = 5;  
    localparam logic [XLEN-1:0] ST_ADDR_MISALIGNED    = 6;
    localparam logic [XLEN-1:0] ST_ACCESS_FAULT       = 7;  
    localparam logic [XLEN-1:0] ENV_CALL_UMODE        = 8;  
    localparam logic [XLEN-1:0] ENV_CALL_SMODE        = 9;  
    localparam logic [XLEN-1:0] ENV_CALL_MMODE        = 11; 
    localparam logic [XLEN-1:0] INSTR_PAGE_FAULT      = 12; 
    localparam logic [XLEN-1:0] LOAD_PAGE_FAULT       = 13; 
    localparam logic [XLEN-1:0] STORE_PAGE_FAULT      = 15; 
    localparam logic [XLEN-1:0] DEBUG_REQUEST         = 24; 
    localparam int unsigned IRQ_S_SOFT  = 1;
    localparam int unsigned IRQ_M_SOFT  = 3;
    localparam int unsigned IRQ_S_TIMER = 5;
    localparam int unsigned IRQ_M_TIMER = 7;
    localparam int unsigned IRQ_S_EXT   = 9;
    localparam int unsigned IRQ_M_EXT   = 11;
    localparam logic [XLEN-1:0] MIP_SSIP = 1 << IRQ_S_SOFT;
    localparam logic [XLEN-1:0] MIP_MSIP = 1 << IRQ_M_SOFT;
    localparam logic [XLEN-1:0] MIP_STIP = 1 << IRQ_S_TIMER;
    localparam logic [XLEN-1:0] MIP_MTIP = 1 << IRQ_M_TIMER;
    localparam logic [XLEN-1:0] MIP_SEIP = 1 << IRQ_S_EXT;
    localparam logic [XLEN-1:0] MIP_MEIP = 1 << IRQ_M_EXT;
    localparam logic [XLEN-1:0] S_SW_INTERRUPT    = (1 << (XLEN-1)) | IRQ_S_SOFT;
    localparam logic [XLEN-1:0] M_SW_INTERRUPT    = (1 << (XLEN-1)) | IRQ_M_SOFT;
    localparam logic [XLEN-1:0] S_TIMER_INTERRUPT = (1 << (XLEN-1)) | IRQ_S_TIMER;
    localparam logic [XLEN-1:0] M_TIMER_INTERRUPT = (1 << (XLEN-1)) | IRQ_M_TIMER;
    localparam logic [XLEN-1:0] S_EXT_INTERRUPT   = (1 << (XLEN-1)) | IRQ_S_EXT;
    localparam logic [XLEN-1:0] M_EXT_INTERRUPT   = (1 << (XLEN-1)) | IRQ_M_EXT;
    
    
    
    typedef enum logic [11:0] {
        
        CSR_FFLAGS         = 12'h001,
        CSR_FRM            = 12'h002,
        CSR_FCSR           = 12'h003,
        CSR_FTRAN          = 12'h800,
        
        CSR_SSTATUS        = 12'h100,
        CSR_SIE            = 12'h104,
        CSR_STVEC          = 12'h105,
        CSR_SCOUNTEREN     = 12'h106,
        CSR_SSCRATCH       = 12'h140,
        CSR_SEPC           = 12'h141,
        CSR_SCAUSE         = 12'h142,
        CSR_STVAL          = 12'h143,
        CSR_SIP            = 12'h144,
        CSR_SATP           = 12'h180,
        
        CSR_MSTATUS        = 12'h300,
        CSR_MISA           = 12'h301,
        CSR_MEDELEG        = 12'h302,
        CSR_MIDELEG        = 12'h303,
        CSR_MIE            = 12'h304,
        CSR_MTVEC          = 12'h305,
        CSR_MCOUNTEREN     = 12'h306,
        CSR_MSCRATCH       = 12'h340,
        CSR_MEPC           = 12'h341,
        CSR_MCAUSE         = 12'h342,
        CSR_MTVAL          = 12'h343,
        CSR_MIP            = 12'h344,
        CSR_PMPCFG0        = 12'h3A0,
        CSR_PMPCFG1        = 12'h3A1,
        CSR_PMPCFG2        = 12'h3A2,
        CSR_PMPCFG3        = 12'h3A3,
        CSR_PMPADDR0       = 12'h3B0,
        CSR_PMPADDR1       = 12'h3B1,
        CSR_PMPADDR2       = 12'h3B2,
        CSR_PMPADDR3       = 12'h3B3,
        CSR_PMPADDR4       = 12'h3B4,
        CSR_PMPADDR5       = 12'h3B5,
        CSR_PMPADDR6       = 12'h3B6,
        CSR_PMPADDR7       = 12'h3B7,
        CSR_PMPADDR8       = 12'h3B8,
        CSR_PMPADDR9       = 12'h3B9,
        CSR_PMPADDR10      = 12'h3BA,
        CSR_PMPADDR11      = 12'h3BB,
        CSR_PMPADDR12      = 12'h3BC,
        CSR_PMPADDR13      = 12'h3BD,
        CSR_PMPADDR14      = 12'h3BE,
        CSR_PMPADDR15      = 12'h3BF,
        CSR_MVENDORID      = 12'hF11,
        CSR_MARCHID        = 12'hF12,
        CSR_MIMPID         = 12'hF13,
        CSR_MHARTID        = 12'hF14,
        CSR_MCYCLE         = 12'hB00,
        CSR_MINSTRET       = 12'hB02,
        
        CSR_ML1_ICACHE_MISS = 12'hB03,  
        CSR_ML1_DCACHE_MISS = 12'hB04,  
        CSR_MITLB_MISS      = 12'hB05,  
        CSR_MDTLB_MISS      = 12'hB06,  
        CSR_MLOAD           = 12'hB07,  
        CSR_MSTORE          = 12'hB08,  
        CSR_MEXCEPTION      = 12'hB09,  
        CSR_MEXCEPTION_RET  = 12'hB0A,  
        CSR_MBRANCH_JUMP    = 12'hB0B,  
        CSR_MCALL           = 12'hB0C,  
        CSR_MRET            = 12'hB0D,  
        CSR_MMIS_PREDICT    = 12'hB0E,  
        CSR_MSB_FULL        = 12'hB0F,  
        CSR_MIF_EMPTY       = 12'hB10,  
        CSR_MHPM_COUNTER_17 = 12'hB11,  
        CSR_MHPM_COUNTER_18 = 12'hB12,  
        CSR_MHPM_COUNTER_19 = 12'hB13,  
        CSR_MHPM_COUNTER_20 = 12'hB14,  
        CSR_MHPM_COUNTER_21 = 12'hB15,  
        CSR_MHPM_COUNTER_22 = 12'hB16,  
        CSR_MHPM_COUNTER_23 = 12'hB17,  
        CSR_MHPM_COUNTER_24 = 12'hB18,  
        CSR_MHPM_COUNTER_25 = 12'hB19,  
        CSR_MHPM_COUNTER_26 = 12'hB1A,  
        CSR_MHPM_COUNTER_27 = 12'hB1B,  
        CSR_MHPM_COUNTER_28 = 12'hB1C,  
        CSR_MHPM_COUNTER_29 = 12'hB1D,  
        CSR_MHPM_COUNTER_30 = 12'hB1E,  
        CSR_MHPM_COUNTER_31 = 12'hB1F,  
        
        CSR_DCACHE         = 12'h701,
        CSR_ICACHE         = 12'h700,
        
        CSR_TSELECT        = 12'h7A0,
        CSR_TDATA1         = 12'h7A1,
        CSR_TDATA2         = 12'h7A2,
        CSR_TDATA3         = 12'h7A3,
        CSR_TINFO          = 12'h7A4,
        
        CSR_DCSR           = 12'h7b0,
        CSR_DPC            = 12'h7b1,
        CSR_DSCRATCH0      = 12'h7b2, 
        CSR_DSCRATCH1      = 12'h7b3, 
        
        CSR_CYCLE          = 12'hC00,
        CSR_TIME           = 12'hC01,
        CSR_INSTRET        = 12'hC02,
        
        CSR_L1_ICACHE_MISS = 12'hC03,  
        CSR_L1_DCACHE_MISS = 12'hC04,  
        CSR_ITLB_MISS      = 12'hC05,  
        CSR_DTLB_MISS      = 12'hC06,  
        CSR_LOAD           = 12'hC07,  
        CSR_STORE          = 12'hC08,  
        CSR_EXCEPTION      = 12'hC09,  
        CSR_EXCEPTION_RET  = 12'hC0A,  
        CSR_BRANCH_JUMP    = 12'hC0B,  
        CSR_CALL           = 12'hC0C,  
        CSR_RET            = 12'hC0D,  
        CSR_MIS_PREDICT    = 12'hC0E,  
        CSR_SB_FULL        = 12'hC0F,  
        CSR_IF_EMPTY       = 12'hC10,  
        CSR_HPM_COUNTER_17 = 12'hC11,  
        CSR_HPM_COUNTER_18 = 12'hC12,  
        CSR_HPM_COUNTER_19 = 12'hC13,  
        CSR_HPM_COUNTER_20 = 12'hC14,  
        CSR_HPM_COUNTER_21 = 12'hC15,  
        CSR_HPM_COUNTER_22 = 12'hC16,  
        CSR_HPM_COUNTER_23 = 12'hC17,  
        CSR_HPM_COUNTER_24 = 12'hC18,  
        CSR_HPM_COUNTER_25 = 12'hC19,  
        CSR_HPM_COUNTER_26 = 12'hC1A,  
        CSR_HPM_COUNTER_27 = 12'hC1B,  
        CSR_HPM_COUNTER_28 = 12'hC1C,  
        CSR_HPM_COUNTER_29 = 12'hC1D,  
        CSR_HPM_COUNTER_30 = 12'hC1E,  
        CSR_HPM_COUNTER_31 = 12'hC1F  
    } csr_reg_t;
    localparam logic [63:0] SSTATUS_UIE  = 'h00000001;
    localparam logic [63:0] SSTATUS_SIE  = 'h00000002;
    localparam logic [63:0] SSTATUS_SPIE = 'h00000020;
    localparam logic [63:0] SSTATUS_SPP  = 'h00000100;
    localparam logic [63:0] SSTATUS_FS   = 'h00006000;
    localparam logic [63:0] SSTATUS_XS   = 'h00018000;
    localparam logic [63:0] SSTATUS_SUM  = 'h00040000;
    localparam logic [63:0] SSTATUS_MXR  = 'h00080000;
    localparam logic [63:0] SSTATUS_UPIE = 'h00000010;
    localparam logic [63:0] SSTATUS_UXL  = 64'h0000000300000000;
    localparam logic [63:0] SSTATUS_SD   = {IS_XLEN64, 31'h00000000, ~IS_XLEN64, 31'h00000000};
    localparam logic [63:0] MSTATUS_UIE  = 'h00000001;
    localparam logic [63:0] MSTATUS_SIE  = 'h00000002;
    localparam logic [63:0] MSTATUS_HIE  = 'h00000004;
    localparam logic [63:0] MSTATUS_MIE  = 'h00000008;
    localparam logic [63:0] MSTATUS_UPIE = 'h00000010;
    localparam logic [63:0] MSTATUS_SPIE = 'h00000020;
    localparam logic [63:0] MSTATUS_HPIE = 'h00000040;
    localparam logic [63:0] MSTATUS_MPIE = 'h00000080;
    localparam logic [63:0] MSTATUS_SPP  = 'h00000100;
    localparam logic [63:0] MSTATUS_HPP  = 'h00000600;
    localparam logic [63:0] MSTATUS_MPP  = 'h00001800;
    localparam logic [63:0] MSTATUS_FS   = 'h00006000;
    localparam logic [63:0] MSTATUS_XS   = 'h00018000;
    localparam logic [63:0] MSTATUS_MPRV = 'h00020000;
    localparam logic [63:0] MSTATUS_SUM  = 'h00040000;
    localparam logic [63:0] MSTATUS_MXR  = 'h00080000;
    localparam logic [63:0] MSTATUS_TVM  = 'h00100000;
    localparam logic [63:0] MSTATUS_TW   = 'h00200000;
    localparam logic [63:0] MSTATUS_TSR  = 'h00400000;
    localparam logic [63:0] MSTATUS_UXL  = {30'h0000000, IS_XLEN64, IS_XLEN64, 32'h00000000};
    localparam logic [63:0] MSTATUS_SXL  = {28'h0000000, IS_XLEN64, IS_XLEN64, 34'h00000000};
    localparam logic [63:0] MSTATUS_SD   = {IS_XLEN64, 31'h00000000, ~IS_XLEN64, 31'h00000000};
    typedef enum logic [2:0] {
        CSRRW  = 3'h1,
        CSRRS  = 3'h2,
        CSRRC  = 3'h3,
        CSRRWI = 3'h5,
        CSRRSI = 3'h6,
        CSRRCI = 3'h7
    } csr_op_t;
    
    typedef struct packed {
        logic [1:0]  rw;
        priv_lvl_t   priv_lvl;
        logic  [7:0] address;
    } csr_addr_t;
    typedef union packed {
        csr_reg_t   address;
        csr_addr_t  csr_decode;
    } csr_t;
    
    typedef struct packed {
        logic [31:15] reserved;  
        logic [6:0]   fprec;     
        logic [2:0]   frm;       
        logic [4:0]   fflags;    
    } fcsr_t;
    
    typedef enum logic [1:0] {
        OFF   = 2'b00,
        TOR   = 2'b01,
        NA4   = 2'b10,
        NAPOT = 2'b11
    } pmp_addr_mode_t;
    
    typedef enum logic [2:0] {
        ACCESS_NONE  = 3'b000,
        ACCESS_READ  = 3'b001,
        ACCESS_WRITE = 3'b010,
        ACCESS_EXEC  = 3'b100
    } pmp_access_t;
    typedef struct packed {
        logic           x;
        logic           w;
        logic           r;
    } pmpcfg_access_t;
    
    typedef struct packed {
        logic           locked;     
        logic [1:0]     reserved;
        pmp_addr_mode_t addr_mode;  
        pmpcfg_access_t access_type;
    } pmpcfg_t;
    
    
    
    typedef struct packed {
        logic [31:28]     xdebugver;
        logic [27:16]     zero2;
        logic             ebreakm;
        logic             zero1;
        logic             ebreaks;
        logic             ebreaku;
        logic             stepie;
        logic             stopcount;
        logic             stoptime;
        logic [8:6]       cause;
        logic             zero0;
        logic             mprven;
        logic             nmip;
        logic             step;
        priv_lvl_t        prv;
    } dcsr_t;
    
    function automatic logic [31:0] jal (logic[4:0] rd, logic [20:0] imm);
        
        return {imm[20], imm[10:1], imm[11], imm[19:12], rd, 7'h6f};
    endfunction
    function automatic logic [31:0] jalr (logic[4:0] rd, logic[4:0] rs1, logic [11:0] offset);
        
        return {offset[11:0], rs1, 3'b0, rd, 7'h67};
    endfunction
    function automatic logic [31:0] andi (logic[4:0] rd, logic[4:0] rs1, logic [11:0] imm);
        
        return {imm[11:0], rs1, 3'h7, rd, 7'h13};
    endfunction
    function automatic logic [31:0] slli (logic[4:0] rd, logic[4:0] rs1, logic [5:0] shamt);
        
        return {6'b0, shamt[5:0], rs1, 3'h1, rd, 7'h13};
    endfunction
    function automatic logic [31:0] srli (logic[4:0] rd, logic[4:0] rs1, logic [5:0] shamt);
        
        return {6'b0, shamt[5:0], rs1, 3'h5, rd, 7'h13};
    endfunction
    function automatic logic [31:0] load (logic [2:0] size, logic[4:0] dest, logic[4:0] base, logic [11:0] offset);
        
        return {offset[11:0], base, size, dest, 7'h03};
    endfunction
    function automatic logic [31:0] auipc (logic[4:0] rd, logic [20:0] imm);
        
        return {imm[20], imm[10:1], imm[11], imm[19:12], rd, 7'h17};
    endfunction
    function automatic logic [31:0] store (logic [2:0] size, logic[4:0] src, logic[4:0] base, logic [11:0] offset);
        
        return {offset[11:5], src, base, size, offset[4:0], 7'h23};
    endfunction
    function automatic logic [31:0] float_load (logic [2:0] size, logic[4:0] dest, logic[4:0] base, logic [11:0] offset);
        
        return {offset[11:0], base, size, dest, 7'b00_001_11};
    endfunction
    function automatic logic [31:0] float_store (logic [2:0] size, logic[4:0] src, logic[4:0] base, logic [11:0] offset);
        
        return {offset[11:5], src, base, size, offset[4:0], 7'b01_001_11};
    endfunction
    function automatic logic [31:0] csrw (csr_reg_t csr, logic[4:0] rs1);
                         
        return {csr, rs1, 3'h1, 5'h0, 7'h73};
    endfunction
    function automatic logic [31:0] csrr (csr_reg_t csr, logic [4:0] dest);
                  
        return {csr, 5'h0, 3'h2, dest, 7'h73};
    endfunction
    function automatic logic [31:0] branch(logic [4:0] src2, logic [4:0] src1, logic [2:0] funct3, logic [11:0] offset);
        
        return {offset[11], offset[9:4], src2, src1, funct3, offset[3:0], offset[10], 7'b11_000_11};
    endfunction
    function automatic logic [31:0] ebreak ();
        return 32'h00100073;
    endfunction
    function automatic logic [31:0] wfi ();
        return 32'h10500073;
    endfunction
    function automatic logic [31:0] nop ();
        return 32'h00000013;
    endfunction
    function automatic logic [31:0] illegal ();
        return 32'h00000000;
    endfunction
    
    
    function string spikeCommitLog(logic [63:0] pc, priv_lvl_t priv_lvl, logic [31:0] instr, logic [4:0] rd, logic [63:0] result, logic rd_fpr);
        string rd_s;
        string instr_word;
        automatic string rf_s = rd_fpr ? "f" : "x";
        if (instr[1:0] != 2'b11) begin
          instr_word = $sformatf("(0x%h)", instr[15:0]);
        end else begin
          instr_word = $sformatf("(0x%h)", instr);
        end
        if (rd < 10) rd_s = $sformatf("%s %0d", rf_s, rd);
        else rd_s = $sformatf("%s%0d", rf_s, rd);
        if (rd_fpr || rd != 0) begin
            
            return $sformatf("%d 0x%h %s %s 0x%h\n", priv_lvl, pc, instr_word, rd_s, result);
        end else begin
            
            return $sformatf("%d 0x%h %s\n", priv_lvl, pc, instr_word);
        end
    endfunction
    typedef struct {
        byte priv;
        longint unsigned pc;
        byte is_fp;
        byte rd;
        longint unsigned data;
        int unsigned instr;
        byte was_exception;
    } commit_log_t;
    
endpackage
package dm;
    localparam logic [3:0] DbgVersion013 = 4'h2;
    
    localparam logic [4:0] ProgBufSize   = 5'h8;
    
    localparam logic [3:0] DataCount     = 4'h2;
    
    localparam logic [63:0] HaltAddress = 64'h800;
    localparam logic [63:0] ResumeAddress = HaltAddress + 4;
    localparam logic [63:0] ExceptionAddress = HaltAddress + 8;
    
    
    localparam logic [11:0] DataAddr = 12'h380; 
    
    typedef enum logic [7:0] {
        Data0        = 8'h04,
        Data1        = 8'h05,
        Data2        = 8'h06,
        Data3        = 8'h07,
        Data4        = 8'h08,
        Data5        = 8'h09,
        Data6        = 8'h0A,
        Data7        = 8'h0B,
        Data8        = 8'h0C,
        Data9        = 8'h0D,
        Data10       = 8'h0E,
        Data11       = 8'h0F,
        DMControl    = 8'h10,
        DMStatus     = 8'h11, 
        Hartinfo     = 8'h12,
        HaltSum1     = 8'h13,
        HAWindowSel  = 8'h14,
        HAWindow     = 8'h15,
        AbstractCS   = 8'h16,
        Command      = 8'h17,
        AbstractAuto = 8'h18,
        DevTreeAddr0 = 8'h19,
        DevTreeAddr1 = 8'h1A,
        DevTreeAddr2 = 8'h1B,
        DevTreeAddr3 = 8'h1C,
        NextDM       = 8'h1D,
        ProgBuf0     = 8'h20,
        ProgBuf15    = 8'h2F,
        AuthData     = 8'h30,
        HaltSum2     = 8'h34,
        HaltSum3     = 8'h35,
        SBAddress3   = 8'h37,
        SBCS         = 8'h38,
        SBAddress0   = 8'h39,
        SBAddress1   = 8'h3A,
        SBAddress2   = 8'h3B,
        SBData0      = 8'h3C,
        SBData1      = 8'h3D,
        SBData2      = 8'h3E,
        SBData3      = 8'h3F,
        HaltSum0     = 8'h40
    } dm_csr_e;
    
    localparam logic [2:0] CauseBreakpoint = 3'h1;
    localparam logic [2:0] CauseTrigger    = 3'h2;
    localparam logic [2:0] CauseRequest    = 3'h3;
    localparam logic [2:0] CauseSingleStep = 3'h4;
    typedef struct packed {
        logic [31:23] zero1;
        logic         impebreak;
        logic [21:20] zero0;
        logic         allhavereset;
        logic         anyhavereset;
        logic         allresumeack;
        logic         anyresumeack;
        logic         allnonexistent;
        logic         anynonexistent;
        logic         allunavail;
        logic         anyunavail;
        logic         allrunning;
        logic         anyrunning;
        logic         allhalted;
        logic         anyhalted;
        logic         authenticated;
        logic         authbusy;
        logic         hasresethaltreq;
        logic         devtreevalid;
        logic [3:0]   version;
    } dmstatus_t;
    typedef struct packed {
        logic         haltreq;
        logic         resumereq;
        logic         hartreset;
        logic         ackhavereset;
        logic         zero1;
        logic         hasel;
        logic [25:16] hartsello;
        logic [15:6]  hartselhi;
        logic [5:4]   zero0;
        logic         setresethaltreq;
        logic         clrresethaltreq;
        logic         ndmreset;
        logic         dmactive;
    } dmcontrol_t;
    typedef struct packed {
        logic [31:24] zero1;
        logic [23:20] nscratch;
        logic [19:17] zero0;
        logic         dataaccess;
        logic [15:12] datasize;
        logic [11:0]  dataaddr;
    } hartinfo_t;
    typedef enum logic [2:0] {  CmdErrNone, CmdErrBusy, CmdErrNotSupported,
                                CmdErrorException, CmdErrorHaltResume,
                                CmdErrorBus, CmdErrorOther = 7
                             } cmderr_e;
    typedef struct packed {
        logic [31:29] zero3;
        logic [28:24] progbufsize;
        logic [23:13] zero2;
        logic         busy;
        logic         zero1;
        cmderr_e      cmderr;
        logic [7:4]   zero0;
        logic [3:0]   datacount;
    } abstractcs_t;
    typedef enum logic [7:0] {
                                 AccessRegister = 8'h0,
                                 QuickAccess    = 8'h1,
                                 AccessMemory   = 8'h2
                             } cmd_e;
    typedef struct packed {
        cmd_e        cmdtype;
        logic [23:0] control;
    } command_t;
    typedef struct packed {
        logic [31:16] autoexecprogbuf;
        logic [15:12] zero0;
        logic [11:0]  autoexecdata;
    } abstractauto_t;
    typedef struct packed {
        logic         zero1;
        logic [22:20] aarsize;
        logic         aarpostincrement;
        logic         postexec;
        logic         transfer;
        logic         write;
        logic [15:0]  regno;
    } ac_ar_cmd_t;
    
    typedef enum logic [1:0] {
        DTM_NOP   = 2'h0,
        DTM_READ  = 2'h1,
        DTM_WRITE = 2'h2
    } dtm_op_e;
    typedef struct packed {
        logic [31:29] sbversion;
        logic [28:23] zero0;
        logic         sbbusyerror;
        logic         sbbusy;
        logic         sbreadonaddr;
        logic [19:17] sbaccess;
        logic         sbautoincrement;
        logic         sbreadondata;
        logic [14:12] sberror;
        logic [11:5]  sbasize;
        logic         sbaccess128;
        logic         sbaccess64;
        logic         sbaccess32;
        logic         sbaccess16;
        logic         sbaccess8;
    } sbcs_t;
    localparam logic[1:0] DTM_SUCCESS = 2'h0;
    typedef struct packed {
        logic [6:0]  addr;
        dtm_op_e     op;
        logic [31:0] data;
    } dmi_req_t;
    typedef struct packed  {
        logic [31:0] data;
        logic [1:0]  resp;
    } dmi_resp_t;
    
    typedef enum logic[1:0] {
      PRIV_LVL_M = 2'b11,
      PRIV_LVL_S = 2'b01,
      PRIV_LVL_U = 2'b00
    } priv_lvl_t;
    
    typedef struct packed {
        logic [31:28]     xdebugver;
        logic [27:16]     zero2;
        logic             ebreakm;
        logic             zero1;
        logic             ebreaks;
        logic             ebreaku;
        logic             stepie;
        logic             stopcount;
        logic             stoptime;
        logic [8:6]       cause;
        logic             zero0;
        logic             mprven;
        logic             nmip;
        logic             step;
        priv_lvl_t        prv;
    } dcsr_t;
    
    typedef enum logic [11:0] {
        
        CSR_FFLAGS         = 12'h001,
        CSR_FRM            = 12'h002,
        CSR_FCSR           = 12'h003,
        CSR_FTRAN          = 12'h800,
        
        CSR_SSTATUS        = 12'h100,
        CSR_SIE            = 12'h104,
        CSR_STVEC          = 12'h105,
        CSR_SCOUNTEREN     = 12'h106,
        CSR_SSCRATCH       = 12'h140,
        CSR_SEPC           = 12'h141,
        CSR_SCAUSE         = 12'h142,
        CSR_STVAL          = 12'h143,
        CSR_SIP            = 12'h144,
        CSR_SATP           = 12'h180,
        
        CSR_MSTATUS        = 12'h300,
        CSR_MISA           = 12'h301,
        CSR_MEDELEG        = 12'h302,
        CSR_MIDELEG        = 12'h303,
        CSR_MIE            = 12'h304,
        CSR_MTVEC          = 12'h305,
        CSR_MCOUNTEREN     = 12'h306,
        CSR_MSCRATCH       = 12'h340,
        CSR_MEPC           = 12'h341,
        CSR_MCAUSE         = 12'h342,
        CSR_MTVAL          = 12'h343,
        CSR_MIP            = 12'h344,
        CSR_PMPCFG0        = 12'h3A0,
        CSR_PMPADDR0       = 12'h3B0,
        CSR_MVENDORID      = 12'hF11,
        CSR_MARCHID        = 12'hF12,
        CSR_MIMPID         = 12'hF13,
        CSR_MHARTID        = 12'hF14,
        CSR_MCYCLE         = 12'hB00,
        CSR_MINSTRET       = 12'hB02,
        CSR_DCACHE         = 12'h701,
        CSR_ICACHE         = 12'h700,
        CSR_TSELECT        = 12'h7A0,
        CSR_TDATA1         = 12'h7A1,
        CSR_TDATA2         = 12'h7A2,
        CSR_TDATA3         = 12'h7A3,
        CSR_TINFO          = 12'h7A4,
        
        CSR_DCSR           = 12'h7b0,
        CSR_DPC            = 12'h7b1,
        CSR_DSCRATCH0      = 12'h7b2, 
        CSR_DSCRATCH1      = 12'h7b3, 
        
        CSR_CYCLE          = 12'hC00,
        CSR_TIME           = 12'hC01,
        CSR_INSTRET        = 12'hC02
    } csr_reg_t;
    
    function automatic logic [31:0] jal (logic[4:0] rd, logic [20:0] imm);
        
        return {imm[20], imm[10:1], imm[11], imm[19:12], rd, 7'h6f};
    endfunction
    function automatic logic [31:0] jalr (logic[4:0] rd, logic[4:0] rs1, logic [11:0] offset);
        
        return {offset[11:0], rs1, 3'b0, rd, 7'h67};
    endfunction
    function automatic logic [31:0] andi (logic[4:0] rd, logic[4:0] rs1, logic [11:0] imm);
        
        return {imm[11:0], rs1, 3'h7, rd, 7'h13};
    endfunction
    function automatic logic [31:0] slli (logic[4:0] rd, logic[4:0] rs1, logic [5:0] shamt);
        
        return {6'b0, shamt[5:0], rs1, 3'h1, rd, 7'h13};
    endfunction
    function automatic logic [31:0] srli (logic[4:0] rd, logic[4:0] rs1, logic [5:0] shamt);
        
        return {6'b0, shamt[5:0], rs1, 3'h5, rd, 7'h13};
    endfunction
    function automatic logic [31:0] load (logic [2:0] size, logic[4:0] dest, logic[4:0] base, logic [11:0] offset);
        
        return {offset[11:0], base, size, dest, 7'h03};
    endfunction
    function automatic logic [31:0] auipc (logic[4:0] rd, logic [20:0] imm);
        
        return {imm[20], imm[10:1], imm[11], imm[19:12], rd, 7'h17};
    endfunction
    function automatic logic [31:0] store (logic [2:0] size, logic[4:0] src, logic[4:0] base, logic [11:0] offset);
        
        return {offset[11:5], src, base, size, offset[4:0], 7'h23};
    endfunction
    function automatic logic [31:0] float_load (logic [2:0] size, logic[4:0] dest, logic[4:0] base, logic [11:0] offset);
        
        return {offset[11:0], base, size, dest, 7'b00_001_11};
    endfunction
    function automatic logic [31:0] float_store (logic [2:0] size, logic[4:0] src, logic[4:0] base, logic [11:0] offset);
        
        return {offset[11:5], src, base, size, offset[4:0], 7'b01_001_11};
    endfunction
    function automatic logic [31:0] csrw (csr_reg_t csr, logic[4:0] rs1);
        
        return {csr, rs1, 3'h1, 5'h0, 7'h73};
    endfunction
    function automatic logic [31:0] csrr (csr_reg_t csr, logic [4:0] dest);
        
        return {csr, 5'h0, 3'h2, dest, 7'h73};
    endfunction
    function automatic logic [31:0] branch(logic [4:0] src2, logic [4:0] src1, logic [2:0] funct3, logic [11:0] offset);
        
        return {offset[11], offset[9:4], src2, src1, funct3, offset[3:0], offset[10], 7'b11_000_11};
    endfunction
    function automatic logic [31:0] ebreak ();
        return 32'h00100073;
    endfunction
    function automatic logic [31:0] wfi ();
        return 32'h10500073;
    endfunction
    function automatic logic [31:0] nop ();
        return 32'h00000013;
    endfunction
    function automatic logic [31:0] illegal ();
        return 32'h00000000;
    endfunction
endpackage
  
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
  
  
  
  
  
  
  
  
 
 
 
package ariane_pkg;
    
    
    
    
    
    
    localparam NrMaxRules = 16;
    typedef struct packed {
      int                               RASDepth;
      int                               BTBEntries;
      int                               BHTEntries;
      
      int unsigned                      NrNonIdempotentRules;  
      logic [NrMaxRules-1:0][63:0]      NonIdempotentAddrBase; 
      logic [NrMaxRules-1:0][63:0]      NonIdempotentLength;   
      int unsigned                      NrExecuteRegionRules;  
      logic [NrMaxRules-1:0][63:0]      ExecuteRegionAddrBase; 
      logic [NrMaxRules-1:0][63:0]      ExecuteRegionLength;   
      int unsigned                      NrCachedRegionRules;   
      logic [NrMaxRules-1:0][63:0]      CachedRegionAddrBase;  
      logic [NrMaxRules-1:0][63:0]      CachedRegionLength;    
      
      bit                               Axi64BitCompliant;     
      bit                               SwapEndianess;         
      
      logic [63:0]                      DmBaseAddress;         
      int unsigned                      NrPMPEntries;          
    } ariane_cfg_t;
    localparam ariane_cfg_t ArianeDefaultConfig = '{
      RASDepth: 2,
      BTBEntries: 32,
      BHTEntries: 128,
      
      NrNonIdempotentRules: 2,
      NonIdempotentAddrBase: {64'b0, 64'b0},
      NonIdempotentLength:   {64'b0, 64'b0},
      NrExecuteRegionRules: 3,
      
      ExecuteRegionAddrBase: {64'h8000_0000, 64'h1_0000, 64'h0},
      ExecuteRegionLength:   {64'h40000000,  64'h10000,  64'h1000},
      
      NrCachedRegionRules:    1,
      CachedRegionAddrBase:  {64'h8000_0000},
      CachedRegionLength:    {64'h40000000},
      
      Axi64BitCompliant:      1'b1,
      SwapEndianess:          1'b0,
      
      DmBaseAddress:          64'h0,
      NrPMPEntries:           8
    };
    
    function automatic void check_cfg (ariane_cfg_t Cfg);
      
      
      
      
    endfunction
    function automatic logic range_check(logic[63:0] base, logic[63:0] len, logic[63:0] address);
      
      return (address >= base) && (address < (base+len));
    endfunction : range_check
    function automatic logic is_inside_nonidempotent_regions (ariane_cfg_t Cfg, logic[63:0] address);
      logic[NrMaxRules-1:0] pass;
      pass = '0;
      for (int unsigned k = 0; k < Cfg.NrNonIdempotentRules; k++) begin
        pass[k] = range_check(Cfg.NonIdempotentAddrBase[k], Cfg.NonIdempotentLength[k], address);
      end
      return |pass;
    endfunction : is_inside_nonidempotent_regions
    function automatic logic is_inside_execute_regions (ariane_cfg_t Cfg, logic[63:0] address);
      
      logic[NrMaxRules-1:0] pass;
      pass = '0;
      for (int unsigned k = 0; k < Cfg.NrExecuteRegionRules; k++) begin
        pass[k] = range_check(Cfg.ExecuteRegionAddrBase[k], Cfg.ExecuteRegionLength[k], address);
      end
      return |pass;
    endfunction : is_inside_execute_regions
    function automatic logic is_inside_cacheable_regions (ariane_cfg_t Cfg, logic[63:0] address);
      automatic logic[NrMaxRules-1:0] pass;
      pass = '0;
      for (int unsigned k = 0; k < Cfg.NrCachedRegionRules; k++) begin
        pass[k] = range_check(Cfg.CachedRegionAddrBase[k], Cfg.CachedRegionLength[k], address);
      end
      return |pass;
    endfunction : is_inside_cacheable_regions
    
    localparam NR_SB_ENTRIES = 8; 
    localparam TRANS_ID_BITS = $clog2(NR_SB_ENTRIES); 
                                                      
    localparam ASID_WIDTH    = (riscv::XLEN == 64) ? 16 : 1;
    localparam BITS_SATURATION_COUNTER = 2;
    localparam NR_COMMIT_PORTS = 2;
    localparam ENABLE_RENAME = 1'b0;
    localparam ISSUE_WIDTH = 1;
    
    
    localparam int unsigned NR_LOAD_PIPE_REGS = 1;
    localparam int unsigned NR_STORE_PIPE_REGS = 0;
    
    localparam int unsigned DEPTH_SPEC   = 4;
    
    localparam int unsigned DEPTH_COMMIT = 8;
    
    localparam bit RVF = riscv::IS_XLEN64; 
    localparam bit RVD = riscv::IS_XLEN64; 
              
    localparam bit RVA = 1'b1; 
    
    localparam bit XF16    = 1'b0; 
    localparam bit XF16ALT = 1'b0; 
    localparam bit XF8     = 1'b0; 
    localparam bit XFVEC   = 1'b0; 
    
    localparam int unsigned LAT_COMP_FP32    = 'd2;
    localparam int unsigned LAT_COMP_FP64    = 'd3;
    localparam int unsigned LAT_COMP_FP16    = 'd1;
    localparam int unsigned LAT_COMP_FP16ALT = 'd1;
    localparam int unsigned LAT_COMP_FP8     = 'd1;
    localparam int unsigned LAT_DIVSQRT      = 'd2;
    localparam int unsigned LAT_NONCOMP      = 'd1;
    localparam int unsigned LAT_CONV         = 'd2;
    
    
    localparam bit FP_PRESENT = RVF | RVD | XF16 | XF16ALT | XF8;
    
    localparam FLEN    = RVD     ? 64 : 
                         RVF     ? 32 : 
                         XF16    ? 16 : 
                         XF16ALT ? 16 : 
                         XF8     ? 8 :  
                         1;             
    localparam bit NSX = XF16 | XF16ALT | XF8 | XFVEC; 
    localparam bit RVFVEC     = RVF     & XFVEC & FLEN>32; 
    localparam bit XF16VEC    = XF16    & XFVEC & FLEN>16; 
    localparam bit XF16ALTVEC = XF16ALT & XFVEC & FLEN>16; 
    localparam bit XF8VEC     = XF8     & XFVEC & FLEN>8;  
    
    
    localparam riscv::xlen_t ARIANE_MARCHID = {{riscv::XLEN-32{1'b0}}, 32'd3};
    localparam riscv::xlen_t ISA_CODE = (RVA <<  0)  
                                     | (1   <<  2)  
                                     | (RVD <<  3)  
                                     | (RVF <<  5)  
                                     | (1   <<  8)  
                                     | (1   << 12)  
                                     | (0   << 13)  
                                     | (1   << 18)  
                                     | (1   << 20)  
                                     | (NSX << 23)  
                                     | ((riscv::XLEN == 64 ? 2 : 1) << riscv::XLEN-2);  
    
    localparam REG_ADDR_SIZE = 6;
    localparam NR_WB_PORTS = 4;
    
    localparam dm::hartinfo_t DebugHartInfo = '{
                                                zero1:        '0,
                                                nscratch:      2, 
                                                zero0:        '0,
                                                dataaccess: 1'b1, 
                                                datasize: dm::DataCount,
                                                dataaddr: dm::DataAddr
                                              };
    
    localparam bit ENABLE_SPIKE_COMMIT_LOG = 1'b1;
    
    
    
    
    localparam logic INVALIDATE_ON_FLUSH = 1'b1;
    localparam bit ENABLE_CYCLE_COUNT = 1'b1;
    localparam bit ENABLE_WFI = 1'b1;
    localparam bit ZERO_TVAL = 1'b0;
    
    localparam logic [63:0] SMODE_STATUS_READ_MASK = riscv::SSTATUS_UIE
                                                   | riscv::SSTATUS_SIE
                                                   | riscv::SSTATUS_SPIE
                                                   | riscv::SSTATUS_SPP
                                                   | riscv::SSTATUS_FS
                                                   | riscv::SSTATUS_XS
                                                   | riscv::SSTATUS_SUM
                                                   | riscv::SSTATUS_MXR
                                                   | riscv::SSTATUS_UPIE
                                                   | riscv::SSTATUS_SPIE
                                                   | riscv::SSTATUS_UXL
                                                   | riscv::SSTATUS_SD;
    localparam logic [63:0] SMODE_STATUS_WRITE_MASK = riscv::SSTATUS_SIE
                                                    | riscv::SSTATUS_SPIE
                                                    | riscv::SSTATUS_SPP
                                                    | riscv::SSTATUS_FS
                                                    | riscv::SSTATUS_SUM
                                                    | riscv::SSTATUS_MXR;
    
    
    
    
    localparam int unsigned FETCH_FIFO_DEPTH  = 4;
    localparam int unsigned FETCH_WIDTH       = 32;
    
    localparam int unsigned INSTR_PER_FETCH = FETCH_WIDTH / 16;
    
    
    typedef struct packed {
         riscv::xlen_t       cause; 
         riscv::xlen_t       tval;  
                             
         logic        valid;
    } exception_t;
    typedef enum logic [2:0] {
      NoCF,   
      Branch, 
      Jump,   
      JumpR,  
      Return  
    } cf_t;
    
    
    
    
    typedef struct packed {
        logic                   valid;           
        logic [riscv::VLEN-1:0] pc;              
        logic [riscv::VLEN-1:0] target_address;  
        logic                   is_mispredict;   
        logic                   is_taken;        
        cf_t                    cf_type;         
    } bp_resolve_t;
    
    
    
    typedef struct packed {
        cf_t                    cf;              
        logic [riscv::VLEN-1:0] predict_address; 
    } branchpredict_sbe_t;
    typedef struct packed {
        logic                   valid;
        logic [riscv::VLEN-1:0] pc;             
        logic [riscv::VLEN-1:0] target_address;
    } btb_update_t;
    typedef struct packed {
        logic                   valid;
        logic [riscv::VLEN-1:0] target_address;
    } btb_prediction_t;
    typedef struct packed {
        logic                   valid;
        logic [riscv::VLEN-1:0] ra;
    } ras_t;
    typedef struct packed {
        logic                   valid;
        logic [riscv::VLEN-1:0] pc;          
        logic                   taken;
    } bht_update_t;
    typedef struct packed {
        logic       valid;
        logic       taken;
    } bht_prediction_t;
    typedef enum logic[3:0] {
        NONE,      
        LOAD,      
        STORE,     
        ALU,       
        CTRL_FLOW, 
        MULT,      
        CSR,       
        FPU,       
        FPU_VEC    
    } fu_t;
    localparam EXC_OFF_RST      = 8'h80;
    localparam SupervisorIrq = 1;
    localparam MachineIrq = 0;
    
    
    typedef struct packed {
      riscv::xlen_t       mie;
      riscv::xlen_t       mip;
      riscv::xlen_t       mideleg;
      logic        sie;
      logic        global_enable;
    } irq_ctrl_t;
    
    
    
    
    localparam int unsigned ICACHE_LINE_WIDTH  = 256;
    localparam int unsigned ICACHE_SET_ASSOC   = 4;
    localparam int unsigned ICACHE_INDEX_WIDTH = $clog2(16384 / ICACHE_SET_ASSOC);
    localparam int unsigned ICACHE_TAG_WIDTH   = riscv::PLEN - ICACHE_INDEX_WIDTH;
    
    localparam int unsigned DCACHE_LINE_WIDTH  = 128;
    localparam int unsigned DCACHE_SET_ASSOC   = 4;
    localparam int unsigned DCACHE_INDEX_WIDTH = $clog2(8192 / DCACHE_SET_ASSOC);
    localparam int unsigned DCACHE_TAG_WIDTH   = riscv::PLEN - DCACHE_INDEX_WIDTH;
 
    
    
    
    typedef enum logic [6:0] { 
                               ADD, SUB, ADDW, SUBW,
                               
                               XORL, ORL, ANDL,
                               
                               SRA, SRL, SLL, SRLW, SLLW, SRAW,
                               
                               LTS, LTU, GES, GEU, EQ, NE,
                               
                               JALR, BRANCH,
                               
                               SLTS, SLTU,
                               
                               MRET, SRET, DRET, ECALL, WFI, FENCE, FENCE_I, SFENCE_VMA, CSR_WRITE, CSR_READ, CSR_SET, CSR_CLEAR,
                               
                               LD, SD, LW, LWU, SW, LH, LHU, SH, LB, SB, LBU,
                               
                               AMO_LRW, AMO_LRD, AMO_SCW, AMO_SCD,
                               AMO_SWAPW, AMO_ADDW, AMO_ANDW, AMO_ORW, AMO_XORW, AMO_MAXW, AMO_MAXWU, AMO_MINW, AMO_MINWU,
                               AMO_SWAPD, AMO_ADDD, AMO_ANDD, AMO_ORD, AMO_XORD, AMO_MAXD, AMO_MAXDU, AMO_MIND, AMO_MINDU,
                               
                               MUL, MULH, MULHU, MULHSU, MULW,
                               
                               DIV, DIVU, DIVW, DIVUW, REM, REMU, REMW, REMUW,
                               
                               FLD, FLW, FLH, FLB, FSD, FSW, FSH, FSB,
                               
                               FADD, FSUB, FMUL, FDIV, FMIN_MAX, FSQRT, FMADD, FMSUB, FNMSUB, FNMADD,
                               
                               FCVT_F2I, FCVT_I2F, FCVT_F2F, FSGNJ, FMV_F2X, FMV_X2F,
                               
                               FCMP,
                               
                               FCLASS,
                               
                               VFMIN, VFMAX, VFSGNJ, VFSGNJN, VFSGNJX, VFEQ, VFNE, VFLT, VFGE, VFLE, VFGT, VFCPKAB_S, VFCPKCD_S, VFCPKAB_D, VFCPKCD_D
                             } fu_op;
    typedef struct packed {
        fu_t                      fu;
        fu_op                     operator;
        riscv::xlen_t             operand_a;
        riscv::xlen_t             operand_b;
        riscv::xlen_t             imm;
        logic [TRANS_ID_BITS-1:0] trans_id;
    } fu_data_t;
    function automatic logic op_is_branch (input fu_op op);
        unique case (op) inside
            EQ, NE, LTS, GES, LTU, GEU: return 1'b1;
            default                   : return 1'b0; 
        endcase
    endfunction
    
    
    
    function automatic logic is_rs1_fpr (input fu_op op);
        if (FP_PRESENT) begin 
            unique case (op) inside
                [FMUL:FNMADD],                   
                FCVT_F2I,                        
                FCVT_F2F,                        
                FSGNJ,                           
                FMV_F2X,                         
                FCMP,                            
                FCLASS,                          
                [VFMIN:VFCPKCD_D] : return 1'b1; 
                default           : return 1'b0; 
            endcase
        end else
            return 1'b0;
    endfunction
    function automatic logic is_rs2_fpr (input fu_op op);
        if (FP_PRESENT) begin 
            unique case (op) inside
                [FSD:FSB],                       
                [FADD:FMIN_MAX],                 
                [FMADD:FNMADD],                  
                FCVT_F2F,                        
                [FSGNJ:FMV_F2X],                 
                FCMP,                            
                [VFMIN:VFCPKCD_D] : return 1'b1; 
                default           : return 1'b0; 
            endcase
        end else
            return 1'b0;
    endfunction
    
    function automatic logic is_imm_fpr (input fu_op op);
        if (FP_PRESENT) begin 
            unique case (op) inside
                [FADD:FSUB],                         
                [FMADD:FNMADD],                      
                [VFCPKAB_S:VFCPKCD_D] : return 1'b1; 
                default               : return 1'b0; 
            endcase
        end else
            return 1'b0;
    endfunction
    function automatic logic is_rd_fpr (input fu_op op);
        if (FP_PRESENT) begin 
            unique case (op) inside
                [FLD:FLB],                           
                [FADD:FNMADD],                       
                FCVT_I2F,                            
                FCVT_F2F,                            
                FSGNJ,                               
                FMV_X2F,                             
                [VFMIN:VFSGNJX],                     
                [VFCPKAB_S:VFCPKCD_D] : return 1'b1; 
                default               : return 1'b0; 
            endcase
        end else
            return 1'b0;
    endfunction
    function automatic logic is_amo (fu_op op);
        case (op) inside
            [AMO_LRW:AMO_MINDU]: begin
                return 1'b1;
            end
            default: return 1'b0;
        endcase
    endfunction
    typedef struct packed {
        logic                     valid;
        logic [riscv::VLEN-1:0]   vaddr;
        logic                     overflow;
        logic [63:0]              data;
        logic [7:0]               be;
        fu_t                      fu;
        fu_op                     operator;
        logic [TRANS_ID_BITS-1:0] trans_id;
    } lsu_ctrl_t;
    
    
    
    
    typedef struct packed {
        logic [riscv::VLEN-1:0] address;        
        logic [31:0]            instruction;    
        branchpredict_sbe_t     branch_predict; 
        exception_t             ex;             
    } fetch_entry_t;
    
    
    
    typedef struct packed {
        logic [riscv::VLEN-1:0]   pc;            
        logic [TRANS_ID_BITS-1:0] trans_id;      
                                                 
        fu_t                      fu;            
        fu_op                     op;            
        logic [REG_ADDR_SIZE-1:0] rs1;           
        logic [REG_ADDR_SIZE-1:0] rs2;           
        logic [REG_ADDR_SIZE-1:0] rd;            
        riscv::xlen_t             result;        
                                                 
                                                 
                                                 
        logic                     valid;         
        logic                     use_imm;       
        logic                     use_zimm;      
        logic                     use_pc;        
        exception_t               ex;            
        branchpredict_sbe_t       bp;            
        logic                     is_compressed; 
                                                 
    } scoreboard_entry_t;
    
    
    
     localparam bit MMU_PRESENT = 1'b1;  
    
    
    
    typedef enum logic [3:0] {
        AMO_NONE =4'b0000,
        AMO_LR   =4'b0001,
        AMO_SC   =4'b0010,
        AMO_SWAP =4'b0011,
        AMO_ADD  =4'b0100,
        AMO_AND  =4'b0101,
        AMO_OR   =4'b0110,
        AMO_XOR  =4'b0111,
        AMO_MAX  =4'b1000,
        AMO_MAXU =4'b1001,
        AMO_MIN  =4'b1010,
        AMO_MINU =4'b1011,
        AMO_CAS1 =4'b1100, 
        AMO_CAS2 =4'b1101  
    } amo_t;
    typedef struct packed {
        logic                  valid;      
        logic                  is_2M;      
        logic                  is_1G;      
        logic [27-1:0]         vpn;        
        logic [ASID_WIDTH-1:0] asid;
        riscv::pte_t           content;
    } tlb_update_t;
    
    
    localparam PPN4K_WIDTH = 38;
    typedef struct packed {
        logic                  valid;      
        logic                  is_4M;      
        logic [20-1:0]         vpn;        
        logic [9-1:0]          asid;       
        riscv::pte_sv32_t      content;
    } tlb_update_sv32_t;
    typedef enum logic [1:0] {
      FE_NONE,
      FE_INSTR_ACCESS_FAULT,
      FE_INSTR_PAGE_FAULT
    } frontend_exception_t;
    
    
    
    
    typedef struct packed {
        logic                     fetch_valid;     
        logic [riscv::PLEN-1:0]   fetch_paddr;     
        exception_t               fetch_exception; 
    } icache_areq_i_t;
    typedef struct packed {
        logic                     fetch_req;       
        logic [riscv::VLEN-1:0]   fetch_vaddr;     
    } icache_areq_o_t;
    
    typedef struct packed {
        logic                     req;                    
        logic                     kill_s1;                
        logic                     kill_s2;                
        logic                     spec;                   
        logic [riscv::VLEN-1:0]   vaddr;                  
    } icache_dreq_i_t;
    typedef struct packed {
        logic                     ready;                  
        logic                     valid;                  
        logic [FETCH_WIDTH-1:0]   data;                   
        logic [riscv::VLEN-1:0]   vaddr;                  
        exception_t               ex;                     
    } icache_dreq_o_t;
    
    
    
    
    typedef struct packed {
        logic        req;       
        amo_t        amo_op;    
        logic [1:0]  size;      
        logic [63:0] operand_a; 
        logic [63:0] operand_b; 
    } amo_req_t;
    
    typedef struct packed {
        logic        ack;    
        logic [63:0] result; 
    } amo_resp_t;
    
    typedef struct packed {
        logic [DCACHE_INDEX_WIDTH-1:0] address_index;
        logic [DCACHE_TAG_WIDTH-1:0]   address_tag;
        logic [63:0]                   data_wdata;
        logic                          data_req;
        logic                          data_we;
        logic [7:0]                    data_be;
        logic [1:0]                    data_size;
        logic                          kill_req;
        logic                          tag_valid;
    } dcache_req_i_t;
    typedef struct packed {
        logic                          data_gnt;
        logic                          data_rvalid;
        logic [63:0]                   data_rdata;
    } dcache_req_o_t;
    
    
    
    function automatic riscv::xlen_t sext32 (logic [31:0] operand);
        return {{riscv::XLEN-32{operand[31]}}, operand[31:0]};
    endfunction
    
    
    
    function automatic logic [riscv::VLEN-1:0] uj_imm (logic [31:0] instruction_i);
        return { {44+riscv::VLEN-64 {instruction_i[31]}}, instruction_i[19:12], instruction_i[20], instruction_i[30:21], 1'b0 };
    endfunction
    function automatic logic [riscv::VLEN-1:0] i_imm (logic [31:0] instruction_i);
        return { {52+riscv::VLEN-64 {instruction_i[31]}}, instruction_i[31:20] };
    endfunction
    function automatic logic [riscv::VLEN-1:0] sb_imm (logic [31:0] instruction_i);
        return { {51+riscv::VLEN-64 {instruction_i[31]}}, instruction_i[31], instruction_i[7], instruction_i[30:25], instruction_i[11:8], 1'b0 };
    endfunction
    
    
    
    
    function automatic riscv::xlen_t data_align (logic [2:0] addr, logic [63:0] data);
        
        logic [2:0] addr_tmp = {(addr[2] && riscv::IS_XLEN64), addr[1:0]};
        logic [63:0] data_tmp = {64{1'b0}};
        case (addr_tmp)
            3'b000: data_tmp[riscv::XLEN-1:0] = {data[riscv::XLEN-1:0]};
            3'b001: data_tmp[riscv::XLEN-1:0] = {data[riscv::XLEN-9:0],  data[riscv::XLEN-1:riscv::XLEN-8]};
            3'b010: data_tmp[riscv::XLEN-1:0] = {data[riscv::XLEN-17:0], data[riscv::XLEN-1:riscv::XLEN-16]};
            3'b011: data_tmp[riscv::XLEN-1:0] = {data[riscv::XLEN-25:0], data[riscv::XLEN-1:riscv::XLEN-24]};
            3'b100: data_tmp = {data[31:0], data[63:32]};
            3'b101: data_tmp = {data[23:0], data[63:24]};
            3'b110: data_tmp = {data[15:0], data[63:16]};
            3'b111: data_tmp = {data[7:0],  data[63:8]};
        endcase
        return data_tmp[riscv::XLEN-1:0];
    endfunction
    
    function automatic logic [7:0] be_gen(logic [2:0] addr, logic [1:0] size);
        case (size)
            2'b11: begin
                return 8'b1111_1111;
            end
            2'b10: begin
                case (addr[2:0])
                    3'b000: return 8'b0000_1111;
                    3'b001: return 8'b0001_1110;
                    3'b010: return 8'b0011_1100;
                    3'b011: return 8'b0111_1000;
                    3'b100: return 8'b1111_0000;
                endcase
            end
            2'b01: begin
                case (addr[2:0])
                    3'b000: return 8'b0000_0011;
                    3'b001: return 8'b0000_0110;
                    3'b010: return 8'b0000_1100;
                    3'b011: return 8'b0001_1000;
                    3'b100: return 8'b0011_0000;
                    3'b101: return 8'b0110_0000;
                    3'b110: return 8'b1100_0000;
                endcase
            end
            2'b00: begin
                case (addr[2:0])
                    3'b000: return 8'b0000_0001;
                    3'b001: return 8'b0000_0010;
                    3'b010: return 8'b0000_0100;
                    3'b011: return 8'b0000_1000;
                    3'b100: return 8'b0001_0000;
                    3'b101: return 8'b0010_0000;
                    3'b110: return 8'b0100_0000;
                    3'b111: return 8'b1000_0000;
                endcase
            end
        endcase
        return 8'b0;
    endfunction
    
    
    
    function automatic logic [1:0] extract_transfer_size(fu_op op);
        case (op)
            LD, SD, FLD, FSD,
            AMO_LRD,   AMO_SCD,
            AMO_SWAPD, AMO_ADDD,
            AMO_ANDD,  AMO_ORD,
            AMO_XORD,  AMO_MAXD,
            AMO_MAXDU, AMO_MIND,
            AMO_MINDU: begin
                return 2'b11;
            end
            LW, LWU, SW, FLW, FSW,
            AMO_LRW,   AMO_SCW,
            AMO_SWAPW, AMO_ADDW,
            AMO_ANDW,  AMO_ORW,
            AMO_XORW,  AMO_MAXW,
            AMO_MAXWU, AMO_MINW,
            AMO_MINWU: begin
                return 2'b10;
            end
            LH, LHU, SH, FLH, FSH: return 2'b01;
            LB, LBU, SB, FLB, FSB: return 2'b00;
            default:     return 2'b11;
        endcase
    endfunction
endpackage
module rrarbiter #(
  parameter int unsigned NUM_REQ   = 64,
  parameter bit          LOCK_IN   = 1'b0
) (
  input logic                         clk_i,
  input logic                         rst_ni,
  input logic                         flush_i, 
  input logic                         en_i,    
  input logic [NUM_REQ-1:0]           req_i,   
  output logic [NUM_REQ-1:0]          ack_o,   
  output logic                        vld_o,   
  output logic [$clog2(NUM_REQ)-1:0]  idx_o    
);
  logic req;
  assign vld_o = (|req_i) & en_i;
  rr_arb_tree #(
    .NumIn     ( NUM_REQ ),
    .DataWidth ( 1       ),
    .LockIn    ( LOCK_IN ))
  i_rr_arb_tree (
    .clk_i   ( clk_i      ),
    .rst_ni  ( rst_ni     ),
    .flush_i ( flush_i    ),
    .rr_i    ( '0         ),
    .req_i   ( req_i      ),
    .gnt_o   ( ack_o      ),
    .data_i  ( '0         ),
    .gnt_i   ( en_i & req ),
    .req_o   ( req        ),
    .data_o  (            ),
    .idx_o   ( idx_o      )
  );
endmodule : rrarbiter
module fifo #(
    parameter bit          FALL_THROUGH = 1'b0, 
    parameter int unsigned DATA_WIDTH   = 32,   
    parameter int unsigned DEPTH        = 8,    
    parameter int unsigned THRESHOLD    = 1,    
    parameter type dtype                = logic [DATA_WIDTH-1:0]
)(
    input  logic  clk_i,            
    input  logic  rst_ni,           
    input  logic  flush_i,          
    input  logic  testmode_i,       
    
    output logic  full_o,           
    output logic  empty_o,          
    output logic  threshold_o,      
    
    input  dtype  data_i,           
    input  logic  push_i,           
    
    output dtype  data_o,           
    input  logic  pop_i             
);
    fifo_v2 #(
        .FALL_THROUGH ( FALL_THROUGH ),
        .DATA_WIDTH   ( DATA_WIDTH   ),
        .DEPTH        ( DEPTH        ),
        .ALM_FULL_TH  ( THRESHOLD    ),
        .dtype        ( dtype        )
    ) impl (
        .clk_i       ( clk_i       ),
        .rst_ni      ( rst_ni      ),
        .flush_i     ( flush_i     ),
        .testmode_i  ( testmode_i  ),
        .full_o      ( full_o      ),
        .empty_o     ( empty_o     ),
        .alm_full_o  ( threshold_o ),
        .alm_empty_o (             ),
        .data_i      ( data_i      ),
        .push_i      ( push_i      ),
        .data_o      ( data_o      ),
        .pop_i       ( pop_i       )
    );
endmodule
module fifo_v2 #(
    parameter bit          FALL_THROUGH = 1'b0, 
    parameter int unsigned DATA_WIDTH   = 32,   
    parameter int unsigned DEPTH        = 8,    
    parameter int unsigned ALM_EMPTY_TH = 1,    
    parameter int unsigned ALM_FULL_TH  = 1,    
    parameter type dtype                = logic [DATA_WIDTH-1:0],
    
    parameter int unsigned ADDR_DEPTH   = (DEPTH > 1) ? $clog2(DEPTH) : 1
)(
    input  logic  clk_i,            
    input  logic  rst_ni,           
    input  logic  flush_i,          
    input  logic  testmode_i,       
    
    output logic  full_o,           
    output logic  empty_o,          
    output logic  alm_full_o,       
    output logic  alm_empty_o,      
    
    input  dtype  data_i,           
    input  logic  push_i,           
    
    output dtype  data_o,           
    input  logic  pop_i             
);
    logic [ADDR_DEPTH-1:0] usage;
    
    if (DEPTH == 0) begin
        assign alm_full_o  = 1'b0; 
        assign alm_empty_o = 1'b0; 
    end else begin
        assign alm_full_o   = (usage >= ALM_FULL_TH[ADDR_DEPTH-1:0]);
        assign alm_empty_o  = (usage <= ALM_EMPTY_TH[ADDR_DEPTH-1:0]);
    end
    fifo_v3 #(
        .FALL_THROUGH ( FALL_THROUGH ),
        .DATA_WIDTH   ( DATA_WIDTH   ),
        .DEPTH        ( DEPTH        ),
        .dtype        ( dtype        )
    ) i_fifo_v3 (
        .clk_i,
        .rst_ni,
        .flush_i,
        .testmode_i,
        .full_o,
        .empty_o,
        .usage_o (usage),
        .data_i,
        .push_i,
        .data_o,
        .pop_i
    );
    
    
    
    
endmodule 
module fifo_v3 #(
    parameter bit          FALL_THROUGH = 1'b0, 
    parameter int unsigned DATA_WIDTH   = 32,   
    parameter int unsigned DEPTH        = 8,    
    parameter type dtype                = logic [DATA_WIDTH-1:0],
    
    parameter int unsigned ADDR_DEPTH   = (DEPTH > 1) ? $clog2(DEPTH) : 1
)(
    input  logic  clk_i,            
    input  logic  rst_ni,           
    input  logic  flush_i,          
    input  logic  testmode_i,       
    
    output logic  full_o,           
    output logic  empty_o,          
    output logic  [ADDR_DEPTH-1:0] usage_o,  
    
    input  dtype  data_i,           
    input  logic  push_i,           
    
    output dtype  data_o,           
    input  logic  pop_i             
);
    
    
    localparam int unsigned FIFO_DEPTH = (DEPTH > 0) ? DEPTH : 1;
    
    logic gate_clock;
    
    logic [ADDR_DEPTH - 1:0] read_pointer_n, read_pointer_q, write_pointer_n, write_pointer_q;
    
    logic [ADDR_DEPTH:0] status_cnt_n, status_cnt_q; 
    
    dtype [FIFO_DEPTH - 1:0] mem_n, mem_q;
    assign usage_o = status_cnt_q[ADDR_DEPTH-1:0];
    if (DEPTH == 0) begin
        assign empty_o     = ~push_i;
        assign full_o      = ~pop_i;
    end else begin
        assign full_o       = (status_cnt_q == FIFO_DEPTH[ADDR_DEPTH:0]);
        assign empty_o      = (status_cnt_q == 0) & ~(FALL_THROUGH & push_i);
    end
    
    
    always_comb begin : read_write_comb
        
        read_pointer_n  = read_pointer_q;
        write_pointer_n = write_pointer_q;
        status_cnt_n    = status_cnt_q;
        data_o          = (DEPTH == 0) ? data_i : mem_q[read_pointer_q];
        mem_n           = mem_q;
        gate_clock      = 1'b1;
        
        if (push_i && ~full_o) begin
            
            mem_n[write_pointer_q] = data_i;
            
            gate_clock = 1'b0;
            
            if (write_pointer_q == FIFO_DEPTH[ADDR_DEPTH-1:0] - 1)
                write_pointer_n = '0;
            else
                write_pointer_n = write_pointer_q + 1;
            
            status_cnt_n    = status_cnt_q + 1;
        end
        if (pop_i && ~empty_o) begin
            
            
            if (read_pointer_n == FIFO_DEPTH[ADDR_DEPTH-1:0] - 1)
                read_pointer_n = '0;
            else
                read_pointer_n = read_pointer_q + 1;
            
            status_cnt_n   = status_cnt_q - 1;
        end
        
        if (push_i && pop_i &&  ~full_o && ~empty_o)
            status_cnt_n   = status_cnt_q;
        
        if (FALL_THROUGH && (status_cnt_q == 0) && push_i) begin
            data_o = data_i;
            if (pop_i) begin
                status_cnt_n = status_cnt_q;
                read_pointer_n = read_pointer_q;
                write_pointer_n = write_pointer_q;
            end
        end
    end
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if(~rst_ni) begin
            read_pointer_q  <= '0;
            write_pointer_q <= '0;
            status_cnt_q    <= '0;
        end else begin
            if (flush_i) begin
                read_pointer_q  <= '0;
                write_pointer_q <= '0;
                status_cnt_q    <= '0;
             end else begin
                read_pointer_q  <= read_pointer_n;
                write_pointer_q <= write_pointer_n;
                status_cnt_q    <= status_cnt_n;
            end
        end
    end
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if(~rst_ni) begin
            mem_q <= '0;
        end else if (!gate_clock) begin
            mem_q <= mem_n;
        end
    end
endmodule 
module lfsr_8bit #(
    parameter logic [7:0]  SEED  = 8'b0,
    parameter int unsigned WIDTH = 8
)(
    input  logic                      clk_i,
    input  logic                      rst_ni,
    input  logic                      en_i,
    output logic [WIDTH-1:0]          refill_way_oh,
    output logic [$clog2(WIDTH)-1:0]  refill_way_bin
);
    localparam int unsigned LOG_WIDTH = $clog2(WIDTH);
    logic [7:0] shift_d, shift_q;
    always_comb begin
        automatic logic shift_in;
        shift_in = !(shift_q[7] ^ shift_q[3] ^ shift_q[2] ^ shift_q[1]);
        shift_d = shift_q;
        if (en_i)
            shift_d = {shift_q[6:0], shift_in};
        
        refill_way_oh = 'b0;
        refill_way_oh[shift_q[LOG_WIDTH-1:0]] = 1'b1;
        refill_way_bin = shift_q;
    end
    always_ff @(posedge clk_i or negedge rst_ni) begin : proc_
        if(~rst_ni) begin
            shift_q <= SEED;
        end else begin
            shift_q <= shift_d;
        end
    end
    
    initial begin
        assert (WIDTH <= 8) else $fatal(1, "WIDTH needs to be less than 8 because of the 8-bit LFSR");
    end
    
endmodule
module lzc #(
  
  parameter int unsigned WIDTH = 2,
  parameter bit          MODE  = 1'b0, 
  
  parameter int unsigned CNT_WIDTH = WIDTH == 1 ? 1 : $clog2(WIDTH)
) (
  input  logic [WIDTH-1:0]     in_i,
  output logic [CNT_WIDTH-1:0] cnt_o,
  output logic                 empty_o 
);
  if (WIDTH == 1) begin: gen_degenerate_lzc
    assign cnt_o[0] = !in_i[0];
    assign empty_o  = !in_i[0];
  end else begin: gen_lzc
    localparam int unsigned NUM_LEVELS = $clog2(WIDTH);
    
    initial begin
      assert(WIDTH > 0) else $fatal(1, "input must be at least one bit wide");
    end
    
    logic [WIDTH-1:0][NUM_LEVELS-1:0]          index_lut;
    logic [2**NUM_LEVELS-1:0]                  sel_nodes;
    logic [2**NUM_LEVELS-1:0][NUM_LEVELS-1:0]  index_nodes;
    logic [WIDTH-1:0] in_tmp;
    
    always_comb begin : flip_vector
      for (int unsigned i = 0; i < WIDTH; i++) begin
        in_tmp[i] = (MODE) ? in_i[WIDTH-1-i] : in_i[i];
      end
    end
    for (genvar j = 0; unsigned'(j) < WIDTH; j++) begin : g_index_lut
      assign index_lut[j] = (NUM_LEVELS)'(unsigned'(j));
    end
    for (genvar level = 0; unsigned'(level) < NUM_LEVELS; level++) begin : g_levels
      if (unsigned'(level) == NUM_LEVELS-1) begin : g_last_level
        for (genvar k = 0; k < 2**level; k++) begin : g_level
          
          if (unsigned'(k) * 2 < WIDTH-1) begin
            assign sel_nodes[2**level-1+k]   = in_tmp[k*2] | in_tmp[k*2+1];
            assign index_nodes[2**level-1+k] = (in_tmp[k*2] == 1'b1) ? index_lut[k*2] :
                                                                       index_lut[k*2+1];
          end
          
          if (unsigned'(k) * 2 == WIDTH-1) begin
            assign sel_nodes[2**level-1+k]   = in_tmp[k*2];
            assign index_nodes[2**level-1+k] = index_lut[k*2];
          end
          
          if (unsigned'(k) * 2 > WIDTH-1) begin
            assign sel_nodes[2**level-1+k]   = 1'b0;
            assign index_nodes[2**level-1+k] = '0;
          end
        end
      end else begin
        for (genvar l = 0; l < 2**level; l++) begin : g_level
          assign sel_nodes[2**level-1+l]   = sel_nodes[2**(level+1)-1+l*2] | sel_nodes[2**(level+1)-1+l*2+1];
          assign index_nodes[2**level-1+l] = (sel_nodes[2**(level+1)-1+l*2] == 1'b1) ? index_nodes[2**(level+1)-1+l*2] :
                                                                                       index_nodes[2**(level+1)-1+l*2+1];
        end
      end
    end
    assign cnt_o   = NUM_LEVELS > unsigned'(0) ? index_nodes[0] : {($clog2(WIDTH)){1'b0}};
    assign empty_o = NUM_LEVELS > unsigned'(0) ? ~sel_nodes[0]  : ~(|in_i);
  end : gen_lzc
endmodule : lzc
module rr_arb_tree #(
  parameter int unsigned NumIn      = 64,
  parameter int unsigned DataWidth  = 32,
  parameter type         DataType   = logic [DataWidth-1:0],
  parameter bit          ExtPrio    = 1'b0, 
  parameter bit          AxiVldRdy  = 1'b0, 
  parameter bit          LockIn     = 1'b0  
) (
  input  logic                             clk_i,
  input  logic                             rst_ni,
  input  logic                             flush_i, 
  input  logic [$clog2(NumIn)-1:0]         rr_i,    
  
  input  logic [NumIn-1:0]                 req_i,
  
  output logic [NumIn-1:0]                 gnt_o,
  
  input  DataType [NumIn-1:0]              data_i,
  
  input  logic                             gnt_i,
  output logic                             req_o,
  output DataType                          data_o,
  output logic [$clog2(NumIn)-1:0]         idx_o
);
  
  
  
  
  
  if (NumIn == unsigned'(1)) begin
    assign req_o    = req_i[0];
    assign gnt_o[0] = gnt_i;
    assign data_o   = data_i[0];
    assign idx_o    = '0;
  
  end else begin
    localparam int unsigned NumLevels = $clog2(NumIn);
    
    logic [2**NumLevels-2:0][NumLevels-1:0]  index_nodes; 
    DataType [2**NumLevels-2:0]              data_nodes;  
    logic [2**NumLevels-2:0]                 gnt_nodes;   
    logic [2**NumLevels-2:0]                 req_nodes;   
    
    logic [NumLevels-1:0]                    rr_q;
    logic [NumIn-1:0]                        req_d;
    
    assign req_o        = req_nodes[0];
    assign data_o       = data_nodes[0];
    assign idx_o        = index_nodes[0];
    if (ExtPrio) begin : gen_ext_rr
      assign rr_q       = rr_i;
      assign req_d      = req_i;
    end else begin : gen_int_rr
      logic [NumLevels-1:0] rr_d;
      
      if (LockIn) begin : gen_lock
        logic  lock_d, lock_q;
        logic [NumIn-1:0]     req_q;
        assign lock_d     = req_o & ~gnt_i;
        assign req_d      = (lock_q) ? req_q : req_i;
        always_ff @(posedge clk_i or negedge rst_ni) begin : p_lock_reg
          if (!rst_ni) begin
            lock_q <= '0;
          end else begin
            if (flush_i) begin
              lock_q <= '0;
            end else begin
              lock_q <= lock_d;
            end
          end
        end
        
        
        
        
        always_ff @(posedge clk_i or negedge rst_ni) begin : p_req_regs
          if (!rst_ni) begin
            req_q  <= '0;
          end else begin
            if (flush_i) begin
              req_q  <= '0;
            end else begin
              req_q  <= req_d;
            end
          end
        end
      end else begin : gen_no_lock
        assign req_d = req_i;
      end
      assign rr_d       = (gnt_i && req_o) ? ((rr_q == NumLevels'(NumIn-1)) ? '0 : rr_q + 1'b1) : rr_q;
      always_ff @(posedge clk_i or negedge rst_ni) begin : p_rr_regs
        if (!rst_ni) begin
          rr_q   <= '0;
        end else begin
          if (flush_i) begin
            rr_q   <= '0;
          end else begin
            rr_q   <= rr_d;
          end
        end
      end
    end
    assign gnt_nodes[0] = gnt_i;
    
    for (genvar level = 0; unsigned'(level) < NumLevels; level++) begin : gen_levels
      for (genvar l = 0; l < 2**level; l++) begin : gen_level
        
        logic sel;
        
        localparam int unsigned idx0 = 2**level-1+l;
        localparam int unsigned idx1 = 2**(level+1)-1+l*2;
        
        
        if (unsigned'(level) == NumLevels-1) begin : gen_first_level
          
          if (unsigned'(l) * 2 < NumIn-1) begin
            assign req_nodes[idx0]   = req_d[l*2] | req_d[l*2+1];
            
            assign sel =  ~req_d[l*2] | req_d[l*2+1] & rr_q[NumLevels-1-level];
            assign index_nodes[idx0] = NumLevels'(sel);
            assign data_nodes[idx0]  = (sel) ? data_i[l*2+1] : data_i[l*2];
            assign gnt_o[l*2]        = gnt_nodes[idx0] & (AxiVldRdy | req_d[l*2])   & ~sel;
            assign gnt_o[l*2+1]      = gnt_nodes[idx0] & (AxiVldRdy | req_d[l*2+1]) & sel;
          end
          
          if (unsigned'(l) * 2 == NumIn-1) begin
            assign req_nodes[idx0]   = req_d[l*2];
            assign index_nodes[idx0] = '0;
            assign data_nodes[idx0]  = data_i[l*2];
            assign gnt_o[l*2]        = gnt_nodes[idx0] & (AxiVldRdy | req_d[l*2]);
          end
          
          if (unsigned'(l) * 2 > NumIn-1) begin
            assign req_nodes[idx0]   = 1'b0;
            assign index_nodes[idx0] = DataType'('0);
            assign data_nodes[idx0]  = DataType'('0);
          end
        
        
        end else begin : gen_other_levels
          assign req_nodes[idx0]   = req_nodes[idx1] | req_nodes[idx1+1];
          
          assign sel =  ~req_nodes[idx1] | req_nodes[idx1+1] & rr_q[NumLevels-1-level];
          assign index_nodes[idx0] = (sel) ? NumLevels'({1'b1, index_nodes[idx1+1][NumLevels-unsigned'(level)-2:0]}) :
                                             NumLevels'({1'b0, index_nodes[idx1][NumLevels-unsigned'(level)-2:0]});
          assign data_nodes[idx0]  = (sel) ? data_nodes[idx1+1] : data_nodes[idx1];
          assign gnt_nodes[idx1]   = gnt_nodes[idx0] & ~sel;
          assign gnt_nodes[idx1+1] = gnt_nodes[idx0] & sel;
        end
        
      end
    end
    
    
    
    
  end
endmodule : rr_arb_tree
module rstgen_bypass #(
    parameter NumRegs = 4
) (
    input  logic clk_i,
    input  logic rst_ni,
    input  logic rst_test_mode_ni,
    input  logic test_mode_i,
    output logic rst_no,
    output logic init_no
);
    
    logic rst_n;
    logic [NumRegs-1:0] synch_regs_q;
    
    always_comb begin
        if (test_mode_i == 1'b0) begin
            rst_n   = rst_ni;
            rst_no  = synch_regs_q[NumRegs-1];
            init_no = synch_regs_q[NumRegs-1];
        end else begin
            rst_n   = rst_test_mode_ni;
            rst_no  = rst_test_mode_ni;
            init_no = 1'b1;
        end
    end
    always @(posedge clk_i or negedge rst_n) begin
        if (~rst_n) begin
            synch_regs_q <= 0;
        end else begin
            synch_regs_q <= {synch_regs_q[NumRegs-2:0], 1'b1};
        end
    end
    initial begin : p_assertions
        if (NumRegs < 1) $fatal(1, "At least one register is required.");
    end
endmodule
module cdc_2phase #(
  parameter type T = logic
)(
  input  logic src_rst_ni,
  input  logic src_clk_i,
  input  T     src_data_i,
  input  logic src_valid_i,
  output logic src_ready_o,
  input  logic dst_rst_ni,
  input  logic dst_clk_i,
  output T     dst_data_o,
  output logic dst_valid_o,
  input  logic dst_ready_i
);
  
  (* dont_touch = "true" *) logic async_req;
  (* dont_touch = "true" *) logic async_ack;
  (* dont_touch = "true" *) T async_data;
  
  cdc_2phase_src #(.T(T)) i_src (
    .rst_ni       ( src_rst_ni  ),
    .clk_i        ( src_clk_i   ),
    .data_i       ( src_data_i  ),
    .valid_i      ( src_valid_i ),
    .ready_o      ( src_ready_o ),
    .async_req_o  ( async_req   ),
    .async_ack_i  ( async_ack   ),
    .async_data_o ( async_data  )
  );
  
  cdc_2phase_dst #(.T(T)) i_dst (
    .rst_ni       ( dst_rst_ni  ),
    .clk_i        ( dst_clk_i   ),
    .data_o       ( dst_data_o  ),
    .valid_o      ( dst_valid_o ),
    .ready_i      ( dst_ready_i ),
    .async_req_i  ( async_req   ),
    .async_ack_o  ( async_ack   ),
    .async_data_i ( async_data  )
  );
endmodule
module cdc_2phase_src #(
  parameter type T = logic
)(
  input  logic rst_ni,
  input  logic clk_i,
  input  T     data_i,
  input  logic valid_i,
  output logic ready_o,
  output logic async_req_o,
  input  logic async_ack_i,
  output T     async_data_o
);
  (* dont_touch = "true" *)
  logic req_src_q, ack_src_q, ack_q;
  (* dont_touch = "true" *)
  T data_src_q;
  
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      req_src_q  <= 0;
      data_src_q <= '0;
    end else if (valid_i && ready_o) begin
      req_src_q  <= ~req_src_q;
      data_src_q <= data_i;
    end
  end
  
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      ack_src_q <= 0;
      ack_q     <= 0;
    end else begin
      ack_src_q <= async_ack_i;
      ack_q     <= ack_src_q;
    end
  end
  
  assign ready_o = (req_src_q == ack_q);
  assign async_req_o = req_src_q;
  assign async_data_o = data_src_q;
endmodule
module cdc_2phase_dst #(
  parameter type T = logic
)(
  input  logic rst_ni,
  input  logic clk_i,
  output T     data_o,
  output logic valid_o,
  input  logic ready_i,
  input  logic async_req_i,
  output logic async_ack_o,
  input  T     async_data_i
);
  (* dont_touch = "true" *)
  (* async_reg = "true" *)
  logic req_dst_q, req_q0, req_q1, ack_dst_q;
  (* dont_touch = "true" *)
  T data_dst_q;
  
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      ack_dst_q  <= 0;
    end else if (valid_o && ready_i) begin
      ack_dst_q  <= ~ack_dst_q;
    end
  end
  
  
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      data_dst_q <= '0;
    end else if (req_q0 != req_q1 && !valid_o) begin
      data_dst_q <= async_data_i;
    end
  end
  
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      req_dst_q <= 0;
      req_q0    <= 0;
      req_q1    <= 0;
    end else begin
      req_dst_q <= async_req_i;
      req_q0    <= req_dst_q;
      req_q1    <= req_q0;
    end
  end
  
  assign valid_o = (ack_dst_q != req_q1);
  assign data_o = data_dst_q;
  assign async_ack_o = ack_dst_q;
endmodule
module shift_reg #(
    parameter type dtype         = logic,
    parameter int unsigned Depth = 1
)(
    input  logic clk_i,    
    input  logic rst_ni,   
    input  dtype d_i,
    output dtype d_o
);
    
    if (Depth == 0) begin
        assign d_o = d_i;
    
    end else if (Depth == 1) begin
        always_ff @(posedge clk_i or negedge rst_ni) begin
            if (~rst_ni) begin
                d_o <= '0;
            end else begin
                d_o <= d_i;
            end
        end
    
    end else if (Depth > 1) begin
        dtype [Depth-1:0] reg_d, reg_q;
        assign d_o = reg_q[Depth-1];
        assign reg_d = {reg_q[Depth-2:0], d_i};
        always_ff @(posedge clk_i or negedge rst_ni) begin
            if (~rst_ni) begin
                reg_q <= '0;
            end else begin
                reg_q <= reg_d;
            end
        end
    end
endmodule
module unread (
    input logic d_i
);
endmodule
module popcount #(
    parameter int unsigned INPUT_WIDTH = 256,
    localparam POPCOUNT_WIDTH          = $clog2(INPUT_WIDTH)+1
) (
    input logic [INPUT_WIDTH-1:0]     data_i,
    output logic [POPCOUNT_WIDTH-1:0] popcount_o
);
   localparam int unsigned PADDED_WIDTH = 1 << $clog2(INPUT_WIDTH);
   logic [PADDED_WIDTH-1:0]           padded_input;
   logic [POPCOUNT_WIDTH-2:0]         left_child_result, right_child_result;
   
   always_comb begin
     padded_input = '0;
     padded_input[INPUT_WIDTH-1:0] = data_i;
   end
   
   if (INPUT_WIDTH == 1) begin : single_node
     assign left_child_result  = 1'b0;
     assign right_child_result = padded_input[0];
   end else if (INPUT_WIDTH == 2) begin : leaf_node
     assign left_child_result  = padded_input[1];
     assign right_child_result = padded_input[0];
   end else begin : non_leaf_node
     popcount #(.INPUT_WIDTH(PADDED_WIDTH / 2))
         left_child(
                    .data_i(padded_input[PADDED_WIDTH-1:PADDED_WIDTH/2]),
                    .popcount_o(left_child_result));
     popcount #(.INPUT_WIDTH(PADDED_WIDTH / 2))
         right_child(
                     .data_i(padded_input[PADDED_WIDTH/2-1:0]),
                     .popcount_o(right_child_result));
   end
   
   assign popcount_o = left_child_result + right_child_result;
endmodule : popcount
module exp_backoff #(
  parameter int unsigned Seed   = 'hffff, 
  parameter int unsigned MaxExp = 16      
) (
  input  logic clk_i,
  input  logic rst_ni,
  
  input  logic set_i,     
  input  logic clr_i,     
  output logic is_zero_o  
);
  
  localparam WIDTH = 16;
  logic [WIDTH-1:0] lfsr_d, lfsr_q, cnt_d, cnt_q, mask_d, mask_q;
  logic lfsr;
  
  
  
  
  assign lfsr = lfsr_q[15-15] ^
                lfsr_q[15-13] ^
                lfsr_q[15-12] ^
                lfsr_q[15-10];
  assign lfsr_d = (set_i) ? {lfsr, lfsr_q[$high(lfsr_q):1]} :
                            lfsr_q;
  
  assign mask_d = (clr_i) ? '0                                :
                  (set_i) ? {{(WIDTH-MaxExp){1'b0}},mask_q[MaxExp-2:0], 1'b1} :
                            mask_q;
  assign cnt_d =  (clr_i)      ? '0                :
                  (set_i)      ? (mask_q & lfsr_q) :
                  (!is_zero_o) ? cnt_q - 1'b1      : '0;
  assign is_zero_o = (cnt_q=='0);
  always_ff @(posedge clk_i or negedge rst_ni) begin : p_regs
    if (!rst_ni) begin
      lfsr_q <= WIDTH'(Seed);
      mask_q <= '0;
      cnt_q  <= '0;
    end else begin
      lfsr_q <= lfsr_d;
      mask_q <= mask_d;
      cnt_q  <= cnt_d;
    end
  end
endmodule 
module apb_to_reg (
  input  logic          clk_i,
  input  logic          rst_ni,
  input  logic          penable_i,
  input  logic          pwrite_i,
  input  logic [31:0]   paddr_i,
  input  logic          psel_i,
  input  logic [31:0]   pwdata_i,
  output logic [31:0]   prdata_o,
  output logic          pready_o,
  output logic          pslverr_o,
  REG_BUS.out  reg_o
);
  always_comb begin
    reg_o.addr = paddr_i;
    reg_o.write = pwrite_i;
    reg_o.wdata = pwdata_i;
    reg_o.wstrb = '1;
    reg_o.valid = psel_i & penable_i;
    pready_o = reg_o.ready;
    pslverr_o = reg_o.error;
    prdata_o = reg_o.rdata;
  end
endmodule
package reg_intf;
    
    typedef struct packed {
        logic [31:0] addr;
        logic        write;
        logic [31:0] wdata;
        logic [3:0]  wstrb;
        logic        valid;
    } reg_intf_req_a32_d32;
    
    typedef struct packed {
        logic [31:0] addr;
        logic        write;
        logic [63:0] wdata;
        logic [7:0]  wstrb;
        logic        valid;
    } reg_intf_req_a32_d64;
    
    typedef struct packed {
        logic [31:0] rdata;
        logic        error;
        logic        ready;
    } reg_intf_resp_d32;
    
    typedef struct packed {
        logic [63:0] rdata;
        logic        error;
        logic        ready;
    } reg_intf_resp_d64;
endpackage
interface REG_BUS #(
  
  parameter int ADDR_WIDTH = -1,
  
  parameter int DATA_WIDTH = -1
)(
  input logic clk_i
);
  logic [ADDR_WIDTH-1:0]   addr;
  logic                    write; 
  logic [DATA_WIDTH-1:0]   rdata;
  logic [DATA_WIDTH-1:0]   wdata;
  logic [DATA_WIDTH/8-1:0] wstrb; 
  logic                    error; 
  logic                    valid;
  logic                    ready;
  modport in  (input  addr, write, wdata, wstrb, valid, output rdata, error, ready);
  modport out (output addr, write, wdata, wstrb, valid, input  rdata, error, ready);
endinterface
package fpnew_pkg;
  
  
  
  
  
  
  
  
  
  
  
  
  typedef struct packed {
    int unsigned exp_bits;
    int unsigned man_bits;
  } fp_encoding_t;
  localparam int unsigned NUM_FP_FORMATS = 5; 
  localparam int unsigned FP_FORMAT_BITS = $clog2(NUM_FP_FORMATS);
  
  typedef enum logic [FP_FORMAT_BITS-1:0] {
    FP32    = 'd0,
    FP64    = 'd1,
    FP16    = 'd2,
    FP8     = 'd3,
    FP16ALT = 'd4
    
  } fp_format_e;
  
  localparam fp_encoding_t [0:NUM_FP_FORMATS-1] FP_ENCODINGS  = '{
    '{8,  23}, 
    '{11, 52}, 
    '{5,  10}, 
    '{5,  2},  
    '{8,  7}   
    
  };
  typedef logic [0:NUM_FP_FORMATS-1]       fmt_logic_t;    
  typedef logic [0:NUM_FP_FORMATS-1][31:0] fmt_unsigned_t; 
  localparam fmt_logic_t CPK_FORMATS = 5'b11000; 
  
  
  
  
  
  
  
  
  
  
  localparam int unsigned NUM_INT_FORMATS = 4; 
  localparam int unsigned INT_FORMAT_BITS = $clog2(NUM_INT_FORMATS);
  
  typedef enum logic [INT_FORMAT_BITS-1:0] {
    INT8,
    INT16,
    INT32,
    INT64
    
  } int_format_e;
  
  function automatic int unsigned int_width(int_format_e ifmt);
    unique case (ifmt)
      INT8:  return 8;
      INT16: return 16;
      INT32: return 32;
      INT64: return 64;
    endcase
  endfunction
  typedef logic [0:NUM_INT_FORMATS-1] ifmt_logic_t; 
  
  
  
  localparam int unsigned NUM_OPGROUPS = 4;
  
  typedef enum logic [1:0] {
    ADDMUL, DIVSQRT, NONCOMP, CONV
  } opgroup_e;
  localparam int unsigned OP_BITS = 4;
  typedef enum logic [OP_BITS-1:0] {
    FMADD, FNMSUB, ADD, MUL,     
    DIV, SQRT,                   
    SGNJ, MINMAX, CMP, CLASSIFY, 
    F2F, F2I, I2F, CPKAB, CPKCD  
  } operation_e;
  
  
  
  
  typedef enum logic [2:0] {
    RNE = 3'b000,
    RTZ = 3'b001,
    RDN = 3'b010,
    RUP = 3'b011,
    RMM = 3'b100,
    DYN = 3'b111
  } roundmode_e;
  
  typedef struct packed {
    logic NV; 
    logic DZ; 
    logic OF; 
    logic UF; 
    logic NX; 
  } status_t;
  
  typedef struct packed {
    logic is_normal;     
    logic is_subnormal;  
    logic is_zero;       
    logic is_inf;        
    logic is_nan;        
    logic is_signalling; 
    logic is_quiet;      
    logic is_boxed;      
  } fp_info_t;
  
  typedef enum logic [9:0] {
    NEGINF     = 10'b00_0000_0001,
    NEGNORM    = 10'b00_0000_0010,
    NEGSUBNORM = 10'b00_0000_0100,
    NEGZERO    = 10'b00_0000_1000,
    POSZERO    = 10'b00_0001_0000,
    POSSUBNORM = 10'b00_0010_0000,
    POSNORM    = 10'b00_0100_0000,
    POSINF     = 10'b00_1000_0000,
    SNAN       = 10'b01_0000_0000,
    QNAN       = 10'b10_0000_0000
  } classmask_e;
  
  
  
  
  typedef enum logic [1:0] {
    BEFORE,     
    AFTER,      
    INSIDE,     
    DISTRIBUTED 
  } pipe_config_t;
  
  typedef enum logic [1:0] {
    DISABLED, 
    PARALLEL, 
    MERGED    
  } unit_type_t;
  
  typedef unit_type_t [0:NUM_FP_FORMATS-1] fmt_unit_types_t;
  
  typedef fmt_unit_types_t [0:NUM_OPGROUPS-1] opgrp_fmt_unit_types_t;
  
  typedef fmt_unsigned_t [0:NUM_OPGROUPS-1] opgrp_fmt_unsigned_t;
  
  typedef struct packed {
    int unsigned Width;
    logic        EnableVectors;
    logic        EnableNanBox;
    fmt_logic_t  FpFmtMask;
    ifmt_logic_t IntFmtMask;
  } fpu_features_t;
  localparam fpu_features_t RV64D = '{
    Width:         64,
    EnableVectors: 1'b0,
    EnableNanBox:  1'b1,
    FpFmtMask:     5'b11000,
    IntFmtMask:    4'b0011
  };
  localparam fpu_features_t RV32D = '{
    Width:         64,
    EnableVectors: 1'b1,
    EnableNanBox:  1'b1,
    FpFmtMask:     5'b11000,
    IntFmtMask:    4'b0010
  };
  localparam fpu_features_t RV32F = '{
    Width:         32,
    EnableVectors: 1'b0,
    EnableNanBox:  1'b1,
    FpFmtMask:     5'b10000,
    IntFmtMask:    4'b0010
  };
  localparam fpu_features_t RV64D_Xsflt = '{
    Width:         64,
    EnableVectors: 1'b1,
    EnableNanBox:  1'b1,
    FpFmtMask:     5'b11111,
    IntFmtMask:    4'b1111
  };
  localparam fpu_features_t RV32F_Xsflt = '{
    Width:         32,
    EnableVectors: 1'b1,
    EnableNanBox:  1'b1,
    FpFmtMask:     5'b10111,
    IntFmtMask:    4'b1110
  };
  localparam fpu_features_t RV32F_Xf16alt_Xfvec = '{
    Width:         32,
    EnableVectors: 1'b1,
    EnableNanBox:  1'b1,
    FpFmtMask:     5'b10001,
    IntFmtMask:    4'b0110
  };
  
  typedef struct packed {
    opgrp_fmt_unsigned_t   PipeRegs;
    opgrp_fmt_unit_types_t UnitTypes;
    pipe_config_t          PipeConfig;
  } fpu_implementation_t;
  localparam fpu_implementation_t DEFAULT_NOREGS = '{
    PipeRegs:   '{default: 0},
    UnitTypes:  '{'{default: PARALLEL}, 
                  '{default: MERGED},   
                  '{default: PARALLEL}, 
                  '{default: MERGED}},  
    PipeConfig: BEFORE
  };
  localparam fpu_implementation_t DEFAULT_SNITCH = '{
    PipeRegs:   '{default: 1},
    UnitTypes:  '{'{default: PARALLEL}, 
                  '{default: DISABLED}, 
                  '{default: PARALLEL}, 
                  '{default: MERGED}},  
    PipeConfig: BEFORE
  };
  
  
  
  localparam logic DONT_CARE = 1'b1; 
  
  
  
  function automatic int minimum(int a, int b);
    return (a < b) ? a : b;
  endfunction
  function automatic int maximum(int a, int b);
    return (a > b) ? a : b;
  endfunction
  
  
  
  
  function automatic int unsigned fp_width(fp_format_e fmt);
    return FP_ENCODINGS[fmt].exp_bits + FP_ENCODINGS[fmt].man_bits + 1;
  endfunction
  
  function automatic int unsigned max_fp_width(fmt_logic_t cfg);
    automatic int unsigned res = 0;
    for (int unsigned i = 0; i < NUM_FP_FORMATS; i++)
      if (cfg[i])
        res = unsigned'(maximum(res, fp_width(fp_format_e'(i))));
    return res;
  endfunction
  
  function automatic int unsigned min_fp_width(fmt_logic_t cfg);
    automatic int unsigned res = max_fp_width(cfg);
    for (int unsigned i = 0; i < NUM_FP_FORMATS; i++)
      if (cfg[i])
        res = unsigned'(minimum(res, fp_width(fp_format_e'(i))));
    return res;
  endfunction
  
  function automatic int unsigned exp_bits(fp_format_e fmt);
    return FP_ENCODINGS[fmt].exp_bits;
  endfunction
  
  function automatic int unsigned man_bits(fp_format_e fmt);
    return FP_ENCODINGS[fmt].man_bits;
  endfunction
  
  function automatic int unsigned bias(fp_format_e fmt);
    return unsigned'(2**(FP_ENCODINGS[fmt].exp_bits-1)-1); 
  endfunction
  function automatic fp_encoding_t super_format(fmt_logic_t cfg);
    automatic fp_encoding_t res;
    res = '0;
    for (int unsigned fmt = 0; fmt < NUM_FP_FORMATS; fmt++)
      if (cfg[fmt]) begin 
        res.exp_bits = unsigned'(maximum(res.exp_bits, exp_bits(fp_format_e'(fmt))));
        res.man_bits = unsigned'(maximum(res.man_bits, man_bits(fp_format_e'(fmt))));
      end
    return res;
  endfunction
  
  
  
  
  function automatic int unsigned max_int_width(ifmt_logic_t cfg);
    automatic int unsigned res = 0;
    for (int ifmt = 0; ifmt < NUM_INT_FORMATS; ifmt++) begin
      if (cfg[ifmt]) res = maximum(res, int_width(int_format_e'(ifmt)));
    end
    return res;
  endfunction
  
  
  
  
  function automatic opgroup_e get_opgroup(operation_e op);
    unique case (op)
      FMADD, FNMSUB, ADD, MUL:     return ADDMUL;
      DIV, SQRT:                   return DIVSQRT;
      SGNJ, MINMAX, CMP, CLASSIFY: return NONCOMP;
      F2F, F2I, I2F, CPKAB, CPKCD: return CONV;
      default:                     return NONCOMP;
    endcase
  endfunction
  
  function automatic int unsigned num_operands(opgroup_e grp);
    unique case (grp)
      ADDMUL:  return 3;
      DIVSQRT: return 2;
      NONCOMP: return 2;
      CONV:    return 3; 
      default: return 0;
    endcase
  endfunction
  
  function automatic int unsigned num_lanes(int unsigned width, fp_format_e fmt, logic vec);
    return vec ? width / fp_width(fmt) : 1; 
  endfunction
  
  function automatic int unsigned max_num_lanes(int unsigned width, fmt_logic_t cfg, logic vec);
    return vec ? width / min_fp_width(cfg) : 1; 
  endfunction
  
  function automatic fmt_logic_t get_lane_formats(int unsigned width,
                                                  fmt_logic_t cfg,
                                                  int unsigned lane_no);
    automatic fmt_logic_t res;
    for (int unsigned fmt = 0; fmt < NUM_FP_FORMATS; fmt++)
      
      res[fmt] = cfg[fmt] & (width / fp_width(fp_format_e'(fmt)) > lane_no);
    return res;
  endfunction
  
  function automatic ifmt_logic_t get_lane_int_formats(int unsigned width,
                                                       fmt_logic_t cfg,
                                                       ifmt_logic_t icfg,
                                                       int unsigned lane_no);
    automatic ifmt_logic_t res;
    automatic fmt_logic_t lanefmts;
    res = '0;
    lanefmts = get_lane_formats(width, cfg, lane_no);
    for (int unsigned ifmt = 0; ifmt < NUM_INT_FORMATS; ifmt++)
      for (int unsigned fmt = 0; fmt < NUM_FP_FORMATS; fmt++)
        
        if ((fp_width(fp_format_e'(fmt)) == int_width(int_format_e'(ifmt))))
          res[ifmt] |= icfg[ifmt] && lanefmts[fmt];
    return res;
  endfunction
  
  function automatic fmt_logic_t get_conv_lane_formats(int unsigned width,
                                                       fmt_logic_t cfg,
                                                       int unsigned lane_no);
    automatic fmt_logic_t res;
    for (int unsigned fmt = 0; fmt < NUM_FP_FORMATS; fmt++)
      
      res[fmt] = cfg[fmt] && ((width / fp_width(fp_format_e'(fmt)) > lane_no) ||
                             (CPK_FORMATS[fmt] && (lane_no < 2)));
    return res;
  endfunction
  
  function automatic ifmt_logic_t get_conv_lane_int_formats(int unsigned width,
                                                            fmt_logic_t cfg,
                                                            ifmt_logic_t icfg,
                                                            int unsigned lane_no);
    automatic ifmt_logic_t res;
    automatic fmt_logic_t lanefmts;
    res = '0;
    lanefmts = get_conv_lane_formats(width, cfg, lane_no);
    for (int unsigned ifmt = 0; ifmt < NUM_INT_FORMATS; ifmt++)
      for (int unsigned fmt = 0; fmt < NUM_FP_FORMATS; fmt++)
        
        res[ifmt] |= icfg[ifmt] && lanefmts[fmt] &&
                     (fp_width(fp_format_e'(fmt)) == int_width(int_format_e'(ifmt)));
    return res;
  endfunction
  
  function automatic logic any_enabled_multi(fmt_unit_types_t types, fmt_logic_t cfg);
    for (int unsigned i = 0; i < NUM_FP_FORMATS; i++)
      if (cfg[i] && types[i] == MERGED)
        return 1'b1;
      return 1'b0;
  endfunction
  
  function automatic logic is_first_enabled_multi(fp_format_e fmt,
                                                  fmt_unit_types_t types,
                                                  fmt_logic_t cfg);
    for (int unsigned i = 0; i < NUM_FP_FORMATS; i++) begin
      if (cfg[i] && types[i] == MERGED) return (fp_format_e'(i) == fmt);
    end
    return 1'b0;
  endfunction
  
  function automatic fp_format_e get_first_enabled_multi(fmt_unit_types_t types, fmt_logic_t cfg);
    for (int unsigned i = 0; i < NUM_FP_FORMATS; i++)
      if (cfg[i] && types[i] == MERGED)
        return fp_format_e'(i);
      return fp_format_e'(0);
  endfunction
  
  function automatic int unsigned get_num_regs_multi(fmt_unsigned_t regs,
                                                     fmt_unit_types_t types,
                                                     fmt_logic_t cfg);
    automatic int unsigned res = 0;
    for (int unsigned i = 0; i < NUM_FP_FORMATS; i++) begin
      if (cfg[i] && types[i] == MERGED) res = maximum(res, regs[i]);
    end
    return res;
  endfunction
endpackage
package defs_div_sqrt_mvp;
   
   localparam C_RM                  = 3;
   localparam C_RM_NEAREST          = 3'h0;
   localparam C_RM_TRUNC            = 3'h1;
   localparam C_RM_PLUSINF          = 3'h2;
   localparam C_RM_MINUSINF         = 3'h3;
   localparam C_PC                  = 6; 
   localparam C_FS                  = 2; 
   localparam C_IUNC                = 2; 
   localparam Iteration_unit_num_S  = 2'b10;
   
   localparam C_OP_FP64             = 64;
   localparam C_MANT_FP64           = 52;
   localparam C_EXP_FP64            = 11;
   localparam C_BIAS_FP64           = 1023;
   localparam C_BIAS_AONE_FP64      = 11'h400;
   localparam C_HALF_BIAS_FP64      = 511;
   localparam C_EXP_ZERO_FP64       = 11'h000;
   localparam C_EXP_ONE_FP64        = 13'h001; 
   localparam C_EXP_INF_FP64        = 11'h7FF;
   localparam C_MANT_ZERO_FP64      = 52'h0;
   localparam C_MANT_NAN_FP64       = 52'h8_0000_0000_0000;
   localparam C_PZERO_FP64          = 64'h0000_0000_0000_0000;
   localparam C_MZERO_FP64          = 64'h8000_0000_0000_0000;
   localparam C_QNAN_FP64           = 64'h7FF8_0000_0000_0000;
   
   localparam C_OP_FP32             = 32;
   localparam C_MANT_FP32           = 23;
   localparam C_EXP_FP32            = 8;
   localparam C_BIAS_FP32           = 127;
   localparam C_BIAS_AONE_FP32      = 8'h80;
   localparam C_HALF_BIAS_FP32      = 63;
   localparam C_EXP_ZERO_FP32       = 8'h00;
   localparam C_EXP_INF_FP32        = 8'hFF;
   localparam C_MANT_ZERO_FP32      = 23'h0;
   localparam C_PZERO_FP32          = 32'h0000_0000;
   localparam C_MZERO_FP32          = 32'h8000_0000;
   localparam C_QNAN_FP32           = 32'h7FC0_0000;
   
   localparam C_OP_FP16             = 16;
   localparam C_MANT_FP16           = 10;
   localparam C_EXP_FP16            = 5;
   localparam C_BIAS_FP16           = 15;
   localparam C_BIAS_AONE_FP16      = 5'h10;
   localparam C_HALF_BIAS_FP16      = 7;
   localparam C_EXP_ZERO_FP16       = 5'h00;
   localparam C_EXP_INF_FP16        = 5'h1F;
   localparam C_MANT_ZERO_FP16      = 10'h0;
   localparam C_PZERO_FP16          = 16'h0000;
   localparam C_MZERO_FP16          = 16'h8000;
   localparam C_QNAN_FP16           = 16'h7E00;
   
   localparam C_OP_FP16ALT           = 16;
   localparam C_MANT_FP16ALT         = 7;
   localparam C_EXP_FP16ALT          = 8;
   localparam C_BIAS_FP16ALT         = 127;
   localparam C_BIAS_AONE_FP16ALT    = 8'h80;
   localparam C_HALF_BIAS_FP16ALT    = 63;
   localparam C_EXP_ZERO_FP16ALT     = 8'h00;
   localparam C_EXP_INF_FP16ALT      = 8'hFF;
   localparam C_MANT_ZERO_FP16ALT    = 7'h0;
   localparam C_QNAN_FP16ALT         = 16'h7FC0;
endpackage : defs_div_sqrt_mvp
import defs_div_sqrt_mvp::*;
module control_mvp
  (
   input logic                                        Clk_CI,
   input logic                                        Rst_RBI,
   input logic                                        Div_start_SI ,
   input logic                                        Sqrt_start_SI,
   input logic                                        Start_SI,
   input logic                                        Kill_SI,
   input logic                                        Special_case_SBI,
   input logic                                        Special_case_dly_SBI,
   input logic [C_PC-1:0]                             Precision_ctl_SI,
   input logic [1:0]                                  Format_sel_SI,
   input logic [C_MANT_FP64:0]                        Numerator_DI,
   input logic [C_EXP_FP64:0]                         Exp_num_DI,
   input logic [C_MANT_FP64:0]                        Denominator_DI,
   input logic [C_EXP_FP64:0]                         Exp_den_DI,
   output logic                                       Div_start_dly_SO ,
   output logic                                       Sqrt_start_dly_SO,
   output logic                                       Div_enable_SO,
   output logic                                       Sqrt_enable_SO,
   
   output logic                                       Full_precision_SO,
   output logic                                       FP32_SO,
   output logic                                       FP64_SO,
   output logic                                       FP16_SO,
   output logic                                       FP16ALT_SO,
   output logic                                       Ready_SO,
   output logic                                       Done_SO,
   output logic [C_MANT_FP64+4:0]                     Mant_result_prenorm_DO,
 
   output logic [C_EXP_FP64+1:0]                      Exp_result_prenorm_DO
 );
   logic  [C_MANT_FP64+1+4:0]                         Partial_remainder_DN,Partial_remainder_DP; 
   logic  [C_MANT_FP64+4:0]                           Quotient_DP; 
   
   
   
   logic [C_MANT_FP64+1:0]                            Numerator_se_D;  
   logic [C_MANT_FP64+1:0]                            Denominator_se_D; 
   logic [C_MANT_FP64+1:0]                            Denominator_se_DB;  
   assign  Numerator_se_D={1'b0,Numerator_DI};
   assign  Denominator_se_D={1'b0,Denominator_DI};
  always_comb
   begin
     if(FP32_SO)
       begin
         Denominator_se_DB={~Denominator_se_D[C_MANT_FP64+1:C_MANT_FP64-C_MANT_FP32], {(C_MANT_FP64-C_MANT_FP32){1'b0}} };
       end
     else if(FP64_SO) begin
         Denominator_se_DB=~Denominator_se_D;
     end
     else if(FP16_SO) begin
         Denominator_se_DB={~Denominator_se_D[C_MANT_FP64+1:C_MANT_FP64-C_MANT_FP16], {(C_MANT_FP64-C_MANT_FP16){1'b0}} };
     end
     else begin
         Denominator_se_DB={~Denominator_se_D[C_MANT_FP64+1:C_MANT_FP64-C_MANT_FP16ALT], {(C_MANT_FP64-C_MANT_FP16ALT){1'b0}} };
     end
   end
   logic [C_MANT_FP64+1:0]                            Mant_D_sqrt_Norm;
   assign Mant_D_sqrt_Norm=Exp_num_DI[0]?{1'b0,Numerator_DI}:{Numerator_DI,1'b0}; 
   
   
   
   logic [1:0]                                      Format_sel_S;
   always_ff @(posedge Clk_CI, negedge Rst_RBI)
     begin
        if(~Rst_RBI)
          begin
            Format_sel_S<='b0;
          end
        else if(Start_SI&&Ready_SO)
          begin
            Format_sel_S<=Format_sel_SI;
          end
        else
          begin
            Format_sel_S<=Format_sel_S;
          end
    end
   assign FP32_SO = (Format_sel_S==2'b00);
   assign FP64_SO = (Format_sel_S==2'b01);
   assign FP16_SO = (Format_sel_S==2'b10);
   assign FP16ALT_SO = (Format_sel_S==2'b11);
   
   
   
   logic [C_PC-1:0]                                   Precision_ctl_S;
   always_ff @(posedge Clk_CI, negedge Rst_RBI)
     begin
        if(~Rst_RBI)
          begin
            Precision_ctl_S<='b0;
          end
        else if(Start_SI&&Ready_SO)
          begin
            Precision_ctl_S<=Precision_ctl_SI;
          end
        else
          begin
            Precision_ctl_S<=Precision_ctl_S;
          end
    end
  assign Full_precision_SO = (Precision_ctl_S==6'h00);
     logic [5:0]                                     State_ctl_S;
     logic [5:0]                                     State_Two_iteration_unit_S;
     logic [5:0]                                     State_Four_iteration_unit_S;
    assign State_Two_iteration_unit_S = Precision_ctl_S[C_PC-1:1];  
    assign State_Four_iteration_unit_S = Precision_ctl_S[C_PC-1:2];  
     always_comb
       begin
         case(Iteration_unit_num_S)
           2'b00:  
             begin
               case(Format_sel_S)
                 2'b00: 
                   begin
                     if(Full_precision_SO)
                       begin
                         State_ctl_S = 6'h1b;  
                       end
                     else
                       begin
                         State_ctl_S = Precision_ctl_S;
                       end
                   end
                 2'b01: 
                   begin
                     if(Full_precision_SO)
                       begin
                         State_ctl_S = 6'h38;  
                       end
                     else
                       begin
                         State_ctl_S = Precision_ctl_S;
                       end
                   end
                 2'b10: 
                   begin
                     if(Full_precision_SO)
                       begin
                         State_ctl_S = 6'h0e;  
                       end
                     else
                       begin
                         State_ctl_S = Precision_ctl_S;
                       end
                   end
                 2'b11: 
                   begin
                     if(Full_precision_SO)
                       begin
                         State_ctl_S = 6'h0b;  
                       end
                     else
                       begin
                         State_ctl_S = Precision_ctl_S;
                       end
                  end
                endcase
              end
           2'b01:  
             begin
               case(Format_sel_S)
                 2'b00: 
                   begin
                     if(Full_precision_SO)
                       begin
                         State_ctl_S = 6'h0d;  
                       end
                     else
                       begin
                         State_ctl_S = State_Two_iteration_unit_S;
                       end
                   end
                 2'b01: 
                   begin
                     if(Full_precision_SO)
                       begin
                         State_ctl_S = 6'h1b;  
                       end
                     else
                       begin
                         State_ctl_S = State_Two_iteration_unit_S;
                       end
                   end
                 2'b10: 
                   begin
                     if(Full_precision_SO)
                       begin
                         State_ctl_S = 6'h06;  
                       end
                     else
                       begin
                         State_ctl_S = State_Two_iteration_unit_S;
                       end
                   end
                 2'b11: 
                   begin
                     if(Full_precision_SO)
                       begin
                         State_ctl_S = 6'h05;  
                       end
                     else
                       begin
                         State_ctl_S = State_Two_iteration_unit_S;
                       end
                  end
                endcase
              end
           2'b10:  
             begin
               case(Format_sel_S)
                 2'b00: 
                   begin
                     case(Precision_ctl_S)
                       6'h00:
                         begin
                           State_ctl_S = 6'h08;  
                         end
                       6'h06,6'h07,6'h08:
                         begin
                           State_ctl_S = 6'h02;
                         end
                       6'h09,6'h0a,6'h0b:
                         begin
                           State_ctl_S = 6'h03;
                         end
                       6'h0c,6'h0d,6'h0e:
                         begin
                           State_ctl_S = 6'h04;
                         end
                       6'h0f,6'h10,6'h11:
                         begin
                           State_ctl_S = 6'h05;
                         end
                       6'h12,6'h13,6'h14:
                         begin
                           State_ctl_S = 6'h06;
                         end
                       6'h15,6'h16,6'h17:
                         begin
                           State_ctl_S = 6'h07;
                         end
                       default:
                         begin
                           State_ctl_S = 6'h08;  
                         end
                     endcase
                   end
                 2'b01: 
                   begin
                     case(Precision_ctl_S)
                       6'h00:
                         begin
                           State_ctl_S = 6'h12;  
                         end
                       6'h06,6'h07,6'h08:
                         begin
                           State_ctl_S = 6'h02;
                         end
                       6'h09,6'h0a,6'h0b:
                         begin
                           State_ctl_S = 6'h03;
                         end
                       6'h0c,6'h0d,6'h0e:
                         begin
                           State_ctl_S = 6'h04;
                         end
                       6'h0f,6'h10,6'h11:
                         begin
                           State_ctl_S = 6'h05;
                         end
                       6'h12,6'h13,6'h14:
                         begin
                           State_ctl_S = 6'h06;
                         end
                       6'h15,6'h16,6'h17:
                         begin
                           State_ctl_S = 6'h07;
                         end
                       6'h18,6'h19,6'h1a:
                         begin
                           State_ctl_S = 6'h08;
                         end
                       6'h1b,6'h1c,6'h1d:
                         begin
                           State_ctl_S = 6'h09;
                         end
                       6'h1e,6'h1f,6'h20:
                         begin
                           State_ctl_S = 6'h0a;
                         end
                       6'h21,6'h22,6'h23:
                         begin
                           State_ctl_S = 6'h0b;
                         end
                       6'h24,6'h25,6'h26:
                         begin
                           State_ctl_S = 6'h0c;
                         end
                       6'h27,6'h28,6'h29:
                         begin
                           State_ctl_S = 6'h0d;
                         end
                       6'h2a,6'h2b,6'h2c:
                         begin
                           State_ctl_S = 6'h0e;
                         end
                       6'h2d,6'h2e,6'h2f:
                         begin
                           State_ctl_S = 6'h0f;
                         end
                       6'h30,6'h31,6'h32:
                         begin
                           State_ctl_S = 6'h10;
                         end
                       6'h33,6'h34,6'h35:
                         begin
                           State_ctl_S = 6'h11;
                         end
                       default:
                         begin
                           State_ctl_S = 6'h12;  
                         end
                     endcase
                   end
                 2'b10: 
                   begin
                     case(Precision_ctl_S)
                       6'h00:
                         begin
                           State_ctl_S = 6'h04;  
                         end
                       6'h06,6'h07,6'h08:
                         begin
                           State_ctl_S = 6'h02;
                         end
                       6'h09,6'h0a,6'h0b:
                         begin
                           State_ctl_S = 6'h03;
                         end
                       default:
                         begin
                           State_ctl_S = 6'h04;  
                         end
                     endcase
                   end
                 2'b11: 
                   begin
                     case(Precision_ctl_S)
                       6'h00:
                         begin
                           State_ctl_S = 6'h03;  
                         end
                       6'h06,6'h07,6'h08:
                         begin
                           State_ctl_S = 6'h02;
                         end
                       default:
                         begin
                           State_ctl_S = 6'h03;  
                         end
                     endcase
                  end
                endcase
              end
           2'b11:  
             begin
               case(Format_sel_S)
                 2'b00: 
                   begin
                     if(Full_precision_SO)
                       begin
                         State_ctl_S = 6'h06;  
                       end
                     else
                       begin
                         State_ctl_S = State_Four_iteration_unit_S;
                       end
                   end
                 2'b01: 
                   begin
                     if(Full_precision_SO)
                       begin
                         State_ctl_S = 6'h0d;  
                       end
                     else
                       begin
                         State_ctl_S = State_Four_iteration_unit_S;
                       end
                   end
                 2'b10: 
                   begin
                     if(Full_precision_SO)
                       begin
                         State_ctl_S = 6'h03;  
                       end
                     else
                       begin
                         State_ctl_S = State_Four_iteration_unit_S;
                       end
                   end
                 2'b11: 
                   begin
                     if(Full_precision_SO)
                       begin
                         State_ctl_S = 6'h02;  
                       end
                     else
                       begin
                         State_ctl_S = State_Four_iteration_unit_S;
                       end
                  end
                endcase
              end
           endcase
        end
   
   
   
   logic                                               Div_start_dly_S;
   always_ff @(posedge Clk_CI, negedge Rst_RBI)   
     begin
        if(~Rst_RBI)
          begin
            Div_start_dly_S<=1'b0;
          end
        else if(Div_start_SI&&Ready_SO)
         begin
           Div_start_dly_S<=1'b1;
         end
        else
          begin
            Div_start_dly_S<=1'b0;
          end
    end
   assign Div_start_dly_SO=Div_start_dly_S;
  always_ff @(posedge Clk_CI, negedge Rst_RBI) begin  
    if(~Rst_RBI)
      Div_enable_SO<=1'b0;
    
    else if (Kill_SI)
      Div_enable_SO <= 1'b0;
    else if(Div_start_SI&&Ready_SO)
      Div_enable_SO<=1'b1;
    else if(Done_SO)
      Div_enable_SO<=1'b0;
    else
      Div_enable_SO<=Div_enable_SO;
  end
   logic                                                Sqrt_start_dly_S;
   always_ff @(posedge Clk_CI, negedge Rst_RBI)   
     begin
        if(~Rst_RBI)
          begin
            Sqrt_start_dly_S<=1'b0;
          end
        else if(Sqrt_start_SI&&Ready_SO)
         begin
           Sqrt_start_dly_S<=1'b1;
         end
        else
          begin
            Sqrt_start_dly_S<=1'b0;
          end
      end
    assign Sqrt_start_dly_SO=Sqrt_start_dly_S;
   always_ff @(posedge Clk_CI, negedge Rst_RBI) begin   
    if(~Rst_RBI)
      Sqrt_enable_SO<=1'b0;
    else if (Kill_SI)
      Sqrt_enable_SO <= 1'b0;
    else if(Sqrt_start_SI&&Ready_SO)
      Sqrt_enable_SO<=1'b1;
    else if(Done_SO)
      Sqrt_enable_SO<=1'b0;
    else
      Sqrt_enable_SO<=Sqrt_enable_SO;
  end
   logic [5:0]                                                  Crtl_cnt_S;
   logic                                                        Start_dly_S;
   assign   Start_dly_S=Div_start_dly_S |Sqrt_start_dly_S;
   logic       Fsm_enable_S;
   assign      Fsm_enable_S=( (Start_dly_S | (| Crtl_cnt_S)) && (~Kill_SI) && Special_case_dly_SBI);
   logic                                                        Final_state_S;
   assign     Final_state_S= (Crtl_cnt_S==State_ctl_S);
   always_ff @(posedge Clk_CI, negedge Rst_RBI) 
     begin
        if (~Rst_RBI)
          begin
             Crtl_cnt_S    <= '0;
          end
          else if (Final_state_S | Kill_SI)
            begin
              Crtl_cnt_S    <= '0;
            end
          else if(Fsm_enable_S) 
            begin
              Crtl_cnt_S    <= Crtl_cnt_S+1;
            end
          else
            begin
              Crtl_cnt_S    <= '0;
            end
     end 
    always_ff @(posedge Clk_CI, negedge Rst_RBI) 
      begin
        if(~Rst_RBI)
          begin
            Done_SO<=1'b0;
          end
        else if(Start_SI&&Ready_SO)
          begin
            if(~Special_case_SBI)
              begin
                Done_SO<=1'b1;
              end
            else
              begin
                Done_SO<=1'b0;
              end
          end
        else if(Final_state_S)
          begin
            Done_SO<=1'b1;
          end
        else
          begin
            Done_SO<=1'b0;
          end
       end
   always_ff @(posedge Clk_CI, negedge Rst_RBI) 
     begin
       if(~Rst_RBI)
         begin
           Ready_SO<=1'b1;
         end
       else if(Start_SI&&Ready_SO)
         begin
            if(~Special_case_SBI)
              begin
                Ready_SO<=1'b1;
              end
            else
              begin
                Ready_SO<=1'b0;
              end
         end
       else if(Final_state_S | Kill_SI)
         begin
           Ready_SO<=1'b1;
         end
       else
         begin
           Ready_SO<=Ready_SO;
         end
     end
  
   
   
  logic                                    Qcnt_one_0;
  logic                                    Qcnt_one_1;
  logic [1:0]                              Qcnt_one_2;
  logic [2:0]                              Qcnt_one_3;
  logic [3:0]                              Qcnt_one_4;
  logic [4:0]                              Qcnt_one_5;
  logic [5:0]                              Qcnt_one_6;
  logic [6:0]                              Qcnt_one_7;
  logic [7:0]                              Qcnt_one_8;
  logic [8:0]                              Qcnt_one_9;
  logic [9:0]                              Qcnt_one_10;
  logic [10:0]                             Qcnt_one_11;
  logic [11:0]                             Qcnt_one_12;
  logic [12:0]                             Qcnt_one_13;
  logic [13:0]                             Qcnt_one_14;
  logic [14:0]                             Qcnt_one_15;
  logic [15:0]                             Qcnt_one_16;
  logic [16:0]                             Qcnt_one_17;
  logic [17:0]                             Qcnt_one_18;
  logic [18:0]                             Qcnt_one_19;
  logic [19:0]                             Qcnt_one_20;
  logic [20:0]                             Qcnt_one_21;
  logic [21:0]                             Qcnt_one_22;
  logic [22:0]                             Qcnt_one_23;
  logic [23:0]                             Qcnt_one_24;
  logic [24:0]                             Qcnt_one_25;
  logic [25:0]                             Qcnt_one_26;
  logic [26:0]                             Qcnt_one_27;
  logic [27:0]                             Qcnt_one_28;
  logic [28:0]                             Qcnt_one_29;
  logic [29:0]                             Qcnt_one_30;
  logic [30:0]                             Qcnt_one_31;
  logic [31:0]                             Qcnt_one_32;
  logic [32:0]                             Qcnt_one_33;
  logic [33:0]                             Qcnt_one_34;
  logic [34:0]                             Qcnt_one_35;
  logic [35:0]                             Qcnt_one_36;
  logic [36:0]                             Qcnt_one_37;
  logic [37:0]                             Qcnt_one_38;
  logic [38:0]                             Qcnt_one_39;
  logic [39:0]                             Qcnt_one_40;
  logic [40:0]                             Qcnt_one_41;
  logic [41:0]                             Qcnt_one_42;
  logic [42:0]                             Qcnt_one_43;
  logic [43:0]                             Qcnt_one_44;
  logic [44:0]                             Qcnt_one_45;
  logic [45:0]                             Qcnt_one_46;
  logic [46:0]                             Qcnt_one_47;
  logic [47:0]                             Qcnt_one_48;
  logic [48:0]                             Qcnt_one_49;
  logic [49:0]                             Qcnt_one_50;
  logic [50:0]                             Qcnt_one_51;
  logic [51:0]                             Qcnt_one_52;
  logic [52:0]                             Qcnt_one_53;
  logic [53:0]                             Qcnt_one_54;
  logic [54:0]                             Qcnt_one_55;
  logic [55:0]                             Qcnt_one_56;
  logic [56:0]                             Qcnt_one_57;
  logic [57:0]                             Qcnt_one_58;
  logic [58:0]                             Qcnt_one_59;
  logic [59:0]                             Qcnt_one_60;
  
   
   
  
   
   
  logic [1:0]                              Qcnt_two_0;
  logic [2:0]                              Qcnt_two_1;
  logic [4:0]                              Qcnt_two_2;
  logic [6:0]                              Qcnt_two_3;
  logic [8:0]                              Qcnt_two_4;
  logic [10:0]                             Qcnt_two_5;
  logic [12:0]                             Qcnt_two_6;
  logic [14:0]                             Qcnt_two_7;
  logic [16:0]                             Qcnt_two_8;
  logic [18:0]                             Qcnt_two_9;
  logic [20:0]                             Qcnt_two_10;
  logic [22:0]                             Qcnt_two_11;
  logic [24:0]                             Qcnt_two_12;
  logic [26:0]                             Qcnt_two_13;
  logic [28:0]                             Qcnt_two_14;
  logic [30:0]                             Qcnt_two_15;
  logic [32:0]                             Qcnt_two_16;
  logic [34:0]                             Qcnt_two_17;
  logic [36:0]                             Qcnt_two_18;
  logic [38:0]                             Qcnt_two_19;
  logic [40:0]                             Qcnt_two_20;
  logic [42:0]                             Qcnt_two_21;
  logic [44:0]                             Qcnt_two_22;
  logic [46:0]                             Qcnt_two_23;
  logic [48:0]                             Qcnt_two_24;
  logic [50:0]                             Qcnt_two_25;
  logic [52:0]                             Qcnt_two_26;
  logic [54:0]                             Qcnt_two_27;
  logic [56:0]                             Qcnt_two_28;
  
   
   
  
   
   
  logic [2:0]                              Qcnt_three_0;
  logic [4:0]                              Qcnt_three_1;
  logic [7:0]                              Qcnt_three_2;
  logic [10:0]                             Qcnt_three_3;
  logic [13:0]                             Qcnt_three_4;
  logic [16:0]                             Qcnt_three_5;
  logic [19:0]                             Qcnt_three_6;
  logic [22:0]                             Qcnt_three_7;
  logic [25:0]                             Qcnt_three_8;
  logic [28:0]                             Qcnt_three_9;
  logic [31:0]                             Qcnt_three_10;
  logic [34:0]                             Qcnt_three_11;
  logic [37:0]                             Qcnt_three_12;
  logic [40:0]                             Qcnt_three_13;
  logic [43:0]                             Qcnt_three_14;
  logic [46:0]                             Qcnt_three_15;
  logic [49:0]                             Qcnt_three_16;
  logic [52:0]                             Qcnt_three_17;
  logic [55:0]                             Qcnt_three_18;
  logic [58:0]                             Qcnt_three_19;
  logic [61:0]                             Qcnt_three_20;
  
   
   
  
   
   
  logic [3:0]                              Qcnt_four_0;
  logic [6:0]                              Qcnt_four_1;
  logic [10:0]                             Qcnt_four_2;
  logic [14:0]                             Qcnt_four_3;
  logic [18:0]                             Qcnt_four_4;
  logic [22:0]                             Qcnt_four_5;
  logic [26:0]                             Qcnt_four_6;
  logic [30:0]                             Qcnt_four_7;
  logic [34:0]                             Qcnt_four_8;
  logic [38:0]                             Qcnt_four_9;
  logic [42:0]                             Qcnt_four_10;
  logic [46:0]                             Qcnt_four_11;
  logic [50:0]                             Qcnt_four_12;
  logic [54:0]                             Qcnt_four_13;
  logic [58:0]                             Qcnt_four_14;
  
   
   
   logic [C_MANT_FP64+1+4:0]                                      Sqrt_R0,Sqrt_Q0,Q_sqrt0,Q_sqrt_com_0;
   logic [C_MANT_FP64+1+4:0]                                      Sqrt_R1,Sqrt_Q1,Q_sqrt1,Q_sqrt_com_1;
   logic [C_MANT_FP64+1+4:0]                                      Sqrt_R2,Sqrt_Q2,Q_sqrt2,Q_sqrt_com_2;
   logic [C_MANT_FP64+1+4:0]                                      Sqrt_R3,Sqrt_Q3,Q_sqrt3,Q_sqrt_com_3,Sqrt_R4; 
   logic [1:0]                                                    Sqrt_DI  [3:0];
   logic [1:0]                                                    Sqrt_DO  [3:0];
   logic                                                          Sqrt_carry_DO;
  logic  [C_MANT_FP64+1+4:0]                                      Iteration_cell_a_D [3:0];
  logic  [C_MANT_FP64+1+4:0]                                      Iteration_cell_b_D [3:0];
  logic  [C_MANT_FP64+1+4:0]                                      Iteration_cell_a_BMASK_D [3:0];
  logic  [C_MANT_FP64+1+4:0]                                      Iteration_cell_b_BMASK_D [3:0];
  logic                                                           Iteration_cell_carry_D [3:0];
  logic  [C_MANT_FP64+1+4:0]                                      Iteration_cell_sum_D [3:0];
  logic  [C_MANT_FP64+1+4:0]                                      Iteration_cell_sum_AMASK_D [3:0];
  logic [3:0]                                                     Sqrt_quotinent_S;
   always_comb
    begin  
      case (Format_sel_S)
        2'b00:
          begin
            Sqrt_quotinent_S = {(~Iteration_cell_sum_AMASK_D[0][C_MANT_FP32+5]),(~Iteration_cell_sum_AMASK_D[1][C_MANT_FP32+5]),(~Iteration_cell_sum_AMASK_D[2][C_MANT_FP32+5]),(~Iteration_cell_sum_AMASK_D[3][C_MANT_FP32+5])};
            Q_sqrt_com_0 ={ {(C_MANT_FP64-C_MANT_FP32){1'b0}},~Q_sqrt0[C_MANT_FP32+5:0] };
            Q_sqrt_com_1 ={ {(C_MANT_FP64-C_MANT_FP32){1'b0}},~Q_sqrt1[C_MANT_FP32+5:0] };
            Q_sqrt_com_2 ={ {(C_MANT_FP64-C_MANT_FP32){1'b0}},~Q_sqrt2[C_MANT_FP32+5:0] };
            Q_sqrt_com_3 ={ {(C_MANT_FP64-C_MANT_FP32){1'b0}},~Q_sqrt3[C_MANT_FP32+5:0] };
          end
        2'b01:
          begin
            Sqrt_quotinent_S = {Iteration_cell_carry_D[0],Iteration_cell_carry_D[1],Iteration_cell_carry_D[2],Iteration_cell_carry_D[3]};
            Q_sqrt_com_0=~Q_sqrt0;
            Q_sqrt_com_1=~Q_sqrt1;
            Q_sqrt_com_2=~Q_sqrt2;
            Q_sqrt_com_3=~Q_sqrt3;
          end
        2'b10:
          begin
            Sqrt_quotinent_S = {(~Iteration_cell_sum_AMASK_D[0][C_MANT_FP16+5]),(~Iteration_cell_sum_AMASK_D[1][C_MANT_FP16+5]),(~Iteration_cell_sum_AMASK_D[2][C_MANT_FP16+5]),(~Iteration_cell_sum_AMASK_D[3][C_MANT_FP16+5])};
            Q_sqrt_com_0 ={ {(C_MANT_FP64-C_MANT_FP16){1'b0}},~Q_sqrt0[C_MANT_FP16+5:0] };
            Q_sqrt_com_1 ={ {(C_MANT_FP64-C_MANT_FP16){1'b0}},~Q_sqrt1[C_MANT_FP16+5:0] };
            Q_sqrt_com_2 ={ {(C_MANT_FP64-C_MANT_FP16){1'b0}},~Q_sqrt2[C_MANT_FP16+5:0] };
            Q_sqrt_com_3 ={ {(C_MANT_FP64-C_MANT_FP16){1'b0}},~Q_sqrt3[C_MANT_FP16+5:0] };
          end
        2'b11:
          begin
            Sqrt_quotinent_S = {(~Iteration_cell_sum_AMASK_D[0][C_MANT_FP16ALT+5]),(~Iteration_cell_sum_AMASK_D[1][C_MANT_FP16ALT+5]),(~Iteration_cell_sum_AMASK_D[2][C_MANT_FP16ALT+5]),(~Iteration_cell_sum_AMASK_D[3][C_MANT_FP16ALT+5])};
            Q_sqrt_com_0 ={ {(C_MANT_FP64-C_MANT_FP16ALT){1'b0}},~Q_sqrt0[C_MANT_FP16ALT+5:0] };
            Q_sqrt_com_1 ={ {(C_MANT_FP64-C_MANT_FP16ALT){1'b0}},~Q_sqrt1[C_MANT_FP16ALT+5:0] };
            Q_sqrt_com_2 ={ {(C_MANT_FP64-C_MANT_FP16ALT){1'b0}},~Q_sqrt2[C_MANT_FP16ALT+5:0] };
            Q_sqrt_com_3 ={ {(C_MANT_FP64-C_MANT_FP16ALT){1'b0}},~Q_sqrt3[C_MANT_FP16ALT+5:0] };
          end
        endcase
    end
  assign  Qcnt_one_0=    {1'b0};  
  assign  Qcnt_one_1=    {Quotient_DP[0]};
  assign  Qcnt_one_2=    {Quotient_DP[1:0]};
  assign  Qcnt_one_3=    {Quotient_DP[2:0]};
  assign  Qcnt_one_4=    {Quotient_DP[3:0]};
  assign  Qcnt_one_5=    {Quotient_DP[4:0]};
  assign  Qcnt_one_6=    {Quotient_DP[5:0]};
  assign  Qcnt_one_7=    {Quotient_DP[6:0]};
  assign  Qcnt_one_8=    {Quotient_DP[7:0]};
  assign  Qcnt_one_9=    {Quotient_DP[8:0]};
  assign  Qcnt_one_10=    {Quotient_DP[9:0]};
  assign  Qcnt_one_11=    {Quotient_DP[10:0]};
  assign  Qcnt_one_12=    {Quotient_DP[11:0]};
  assign  Qcnt_one_13=    {Quotient_DP[12:0]};
  assign  Qcnt_one_14=    {Quotient_DP[13:0]};
  assign  Qcnt_one_15=    {Quotient_DP[14:0]};
  assign  Qcnt_one_16=    {Quotient_DP[15:0]};
  assign  Qcnt_one_17=    {Quotient_DP[16:0]};
  assign  Qcnt_one_18=    {Quotient_DP[17:0]};
  assign  Qcnt_one_19=    {Quotient_DP[18:0]};
  assign  Qcnt_one_20=    {Quotient_DP[19:0]};
  assign  Qcnt_one_21=    {Quotient_DP[20:0]};
  assign  Qcnt_one_22=    {Quotient_DP[21:0]};
  assign  Qcnt_one_23=    {Quotient_DP[22:0]};
  assign  Qcnt_one_24=    {Quotient_DP[23:0]};
  assign  Qcnt_one_25=    {Quotient_DP[24:0]};
  assign  Qcnt_one_26=    {Quotient_DP[25:0]};
  assign  Qcnt_one_27=    {Quotient_DP[26:0]};
  assign  Qcnt_one_28=    {Quotient_DP[27:0]};
  assign  Qcnt_one_29=    {Quotient_DP[28:0]};
  assign  Qcnt_one_30=    {Quotient_DP[29:0]};
  assign  Qcnt_one_31=    {Quotient_DP[30:0]};
  assign  Qcnt_one_32=    {Quotient_DP[31:0]};
  assign  Qcnt_one_33=    {Quotient_DP[32:0]};
  assign  Qcnt_one_34=    {Quotient_DP[33:0]};
  assign  Qcnt_one_35=    {Quotient_DP[34:0]};
  assign  Qcnt_one_36=    {Quotient_DP[35:0]};
  assign  Qcnt_one_37=    {Quotient_DP[36:0]};
  assign  Qcnt_one_38=    {Quotient_DP[37:0]};
  assign  Qcnt_one_39=    {Quotient_DP[38:0]};
  assign  Qcnt_one_40=    {Quotient_DP[39:0]};
  assign  Qcnt_one_41=    {Quotient_DP[40:0]};
  assign  Qcnt_one_42=    {Quotient_DP[41:0]};
  assign  Qcnt_one_43=    {Quotient_DP[42:0]};
  assign  Qcnt_one_44=    {Quotient_DP[43:0]};
  assign  Qcnt_one_45=    {Quotient_DP[44:0]};
  assign  Qcnt_one_46=    {Quotient_DP[45:0]};
  assign  Qcnt_one_47=    {Quotient_DP[46:0]};
  assign  Qcnt_one_48=    {Quotient_DP[47:0]};
  assign  Qcnt_one_49=    {Quotient_DP[48:0]};
  assign  Qcnt_one_50=    {Quotient_DP[49:0]};
  assign  Qcnt_one_51=    {Quotient_DP[50:0]};
  assign  Qcnt_one_52=    {Quotient_DP[51:0]};
  assign  Qcnt_one_53=    {Quotient_DP[52:0]};
  assign  Qcnt_one_54=    {Quotient_DP[53:0]};
  assign  Qcnt_one_55=    {Quotient_DP[54:0]};
  assign  Qcnt_one_56=    {Quotient_DP[55:0]};
  assign  Qcnt_one_57=    {Quotient_DP[56:0]};
  assign  Qcnt_two_0 =    {1'b0,            Sqrt_quotinent_S[3]};  
  assign  Qcnt_two_1 =    {Quotient_DP[1:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_2 =    {Quotient_DP[3:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_3 =    {Quotient_DP[5:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_4 =    {Quotient_DP[7:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_5 =    {Quotient_DP[9:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_6 =    {Quotient_DP[11:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_7 =    {Quotient_DP[13:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_8 =    {Quotient_DP[15:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_9 =    {Quotient_DP[17:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_10 =    {Quotient_DP[19:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_11 =    {Quotient_DP[21:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_12 =    {Quotient_DP[23:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_13 =    {Quotient_DP[25:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_14 =    {Quotient_DP[27:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_15 =    {Quotient_DP[29:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_16 =    {Quotient_DP[31:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_17 =    {Quotient_DP[33:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_18 =    {Quotient_DP[35:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_19 =    {Quotient_DP[37:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_20 =    {Quotient_DP[39:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_21 =    {Quotient_DP[41:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_22 =    {Quotient_DP[43:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_23 =    {Quotient_DP[45:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_24 =    {Quotient_DP[47:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_25 =    {Quotient_DP[49:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_26 =    {Quotient_DP[51:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_27 =    {Quotient_DP[53:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_two_28 =    {Quotient_DP[55:0],Sqrt_quotinent_S[3]};
  assign  Qcnt_three_0 =    {1'b0,            Sqrt_quotinent_S[3],Sqrt_quotinent_S[2]};  
  assign  Qcnt_three_1 =    {Quotient_DP[2:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2]};
  assign  Qcnt_three_2 =    {Quotient_DP[5:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2]};
  assign  Qcnt_three_3 =    {Quotient_DP[8:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2]};
  assign  Qcnt_three_4 =    {Quotient_DP[11:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2]};
  assign  Qcnt_three_5 =    {Quotient_DP[14:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2]};
  assign  Qcnt_three_6 =    {Quotient_DP[17:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2]};
  assign  Qcnt_three_7 =    {Quotient_DP[20:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2]};
  assign  Qcnt_three_8 =    {Quotient_DP[23:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2]};
  assign  Qcnt_three_9 =    {Quotient_DP[26:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2]};
  assign  Qcnt_three_10 =    {Quotient_DP[29:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2]};
  assign  Qcnt_three_11 =    {Quotient_DP[32:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2]};
  assign  Qcnt_three_12 =    {Quotient_DP[35:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2]};
  assign  Qcnt_three_13 =    {Quotient_DP[38:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2]};
  assign  Qcnt_three_14 =    {Quotient_DP[41:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2]};
  assign  Qcnt_three_15 =    {Quotient_DP[44:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2]};
  assign  Qcnt_three_16 =    {Quotient_DP[47:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2]};
  assign  Qcnt_three_17 =    {Quotient_DP[50:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2]};
  assign  Qcnt_three_18 =    {Quotient_DP[53:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2]};
  assign  Qcnt_three_19 =    {Quotient_DP[56:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2]};
  assign      Qcnt_four_0 =    {1'b0,            Sqrt_quotinent_S[3],Sqrt_quotinent_S[2],Sqrt_quotinent_S[1]};
  assign      Qcnt_four_1 =    {Quotient_DP[3:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2],Sqrt_quotinent_S[1]};
  assign      Qcnt_four_2 =    {Quotient_DP[7:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2],Sqrt_quotinent_S[1]};
  assign      Qcnt_four_3 =    {Quotient_DP[11:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2],Sqrt_quotinent_S[1]};
  assign      Qcnt_four_4 =    {Quotient_DP[15:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2],Sqrt_quotinent_S[1]};
  assign      Qcnt_four_5 =    {Quotient_DP[19:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2],Sqrt_quotinent_S[1]};
  assign      Qcnt_four_6 =    {Quotient_DP[23:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2],Sqrt_quotinent_S[1]};
  assign      Qcnt_four_7 =    {Quotient_DP[27:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2],Sqrt_quotinent_S[1]};
  assign      Qcnt_four_8 =    {Quotient_DP[31:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2],Sqrt_quotinent_S[1]};
  assign      Qcnt_four_9 =    {Quotient_DP[35:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2],Sqrt_quotinent_S[1]};
  assign      Qcnt_four_10 =    {Quotient_DP[39:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2],Sqrt_quotinent_S[1]};
  assign      Qcnt_four_11 =    {Quotient_DP[43:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2],Sqrt_quotinent_S[1]};
  assign      Qcnt_four_12 =    {Quotient_DP[47:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2],Sqrt_quotinent_S[1]};
  assign      Qcnt_four_13 =    {Quotient_DP[51:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2],Sqrt_quotinent_S[1]};
  assign      Qcnt_four_14 =    {Quotient_DP[55:0],Sqrt_quotinent_S[3],Sqrt_quotinent_S[2],Sqrt_quotinent_S[1]};
  always_comb begin  
  case(Iteration_unit_num_S)
    2'b00:
      begin
  
   
   
        case(Crtl_cnt_S)
          6'b000000:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64+1:C_MANT_FP64];
              Q_sqrt0={{(C_MANT_FP64+5){1'b0}},Qcnt_one_0};
              Sqrt_Q0=Q_sqrt_com_0;
            end
          6'b000001:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-1:C_MANT_FP64-2];
              Q_sqrt0={{(C_MANT_FP64+5){1'b0}},Qcnt_one_1};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b000010:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-3:C_MANT_FP64-4];
              Q_sqrt0={{(C_MANT_FP64+4){1'b0}},Qcnt_one_2};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b000011:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-5:C_MANT_FP64-6];
              Q_sqrt0={{(C_MANT_FP64+3){1'b0}},Qcnt_one_3};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b000100:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-7:C_MANT_FP64-8];
              Q_sqrt0={{(C_MANT_FP64+2){1'b0}},Qcnt_one_4};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b000101:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-9:C_MANT_FP64-10];
              Q_sqrt0={{(C_MANT_FP64+1){1'b0}},Qcnt_one_5};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b000110:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-11:C_MANT_FP64-12];
              Q_sqrt0={{(C_MANT_FP64){1'b0}},Qcnt_one_6};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b000111:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-13:C_MANT_FP64-14];
              Q_sqrt0={{(C_MANT_FP64-1){1'b0}},Qcnt_one_7};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b001000:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-15:C_MANT_FP64-16];
              Q_sqrt0={{(C_MANT_FP64-2){1'b0}},Qcnt_one_8};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b001001:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-17:C_MANT_FP64-18];
              Q_sqrt0={{(C_MANT_FP64-3){1'b0}},Qcnt_one_9};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b001010:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-19:C_MANT_FP64-20];
              Q_sqrt0={{(C_MANT_FP64-4){1'b0}},Qcnt_one_10};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b001011:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-21:C_MANT_FP64-22];
              Q_sqrt0={{(C_MANT_FP64-5){1'b0}},Qcnt_one_11};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b001100:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-23:C_MANT_FP64-24];
              Q_sqrt0={{(C_MANT_FP64-6){1'b0}},Qcnt_one_12};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b001101:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-25:C_MANT_FP64-26];
              Q_sqrt0={{(C_MANT_FP64-7){1'b0}},Qcnt_one_13};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b001110:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-27:C_MANT_FP64-28];
              Q_sqrt0={{(C_MANT_FP64-8){1'b0}},Qcnt_one_14};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b001111:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-29:C_MANT_FP64-30];
              Q_sqrt0={{(C_MANT_FP64-9){1'b0}},Qcnt_one_15};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b010000:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-31:C_MANT_FP64-32];
              Q_sqrt0={{(C_MANT_FP64-10){1'b0}},Qcnt_one_16};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b010001:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-33:C_MANT_FP64-34];
              Q_sqrt0={{(C_MANT_FP64-11){1'b0}},Qcnt_one_17};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b010010:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-35:C_MANT_FP64-36];
              Q_sqrt0={{(C_MANT_FP64-12){1'b0}},Qcnt_one_18};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b010011:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-37:C_MANT_FP64-38];
              Q_sqrt0={{(C_MANT_FP64-13){1'b0}},Qcnt_one_19};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b010100:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-39:C_MANT_FP64-40];
              Q_sqrt0={{(C_MANT_FP64-14){1'b0}},Qcnt_one_20};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b010101:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-41:C_MANT_FP64-42];
              Q_sqrt0={{(C_MANT_FP64-15){1'b0}},Qcnt_one_21};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b010110:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-43:C_MANT_FP64-44];
              Q_sqrt0={{(C_MANT_FP64-16){1'b0}},Qcnt_one_22};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b010111:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-45:C_MANT_FP64-46];
              Q_sqrt0={{(C_MANT_FP64-17){1'b0}},Qcnt_one_23};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b011000:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-47:C_MANT_FP64-48];
              Q_sqrt0={{(C_MANT_FP64-18){1'b0}},Qcnt_one_24};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b011001:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-49:C_MANT_FP64-50];
              Q_sqrt0={{(C_MANT_FP64-19){1'b0}},Qcnt_one_25};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b011010:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-51:C_MANT_FP64-52];
              Q_sqrt0={{(C_MANT_FP64-20){1'b0}},Qcnt_one_26};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b011011:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-21){1'b0}},Qcnt_one_27};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b011100:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-22){1'b0}},Qcnt_one_28};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b011101:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-23){1'b0}},Qcnt_one_29};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b011110:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-24){1'b0}},Qcnt_one_30};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b011111:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-25){1'b0}},Qcnt_one_31};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b100000:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-26){1'b0}},Qcnt_one_32};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b100001:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-27){1'b0}},Qcnt_one_33};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b100010:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-28){1'b0}},Qcnt_one_34};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b100011:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-29){1'b0}},Qcnt_one_35};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b100100:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-30){1'b0}},Qcnt_one_36};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b100101:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-31){1'b0}},Qcnt_one_37};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b100110:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-32){1'b0}},Qcnt_one_38};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b100111:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-33){1'b0}},Qcnt_one_39};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b101000:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-34){1'b0}},Qcnt_one_40};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b101001:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-35){1'b0}},Qcnt_one_41};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b101010:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-36){1'b0}},Qcnt_one_42};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b101011:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-37){1'b0}},Qcnt_one_43};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b101100:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-38){1'b0}},Qcnt_one_44};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b101101:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-39){1'b0}},Qcnt_one_45};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b101110:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-40){1'b0}},Qcnt_one_46};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b101111:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-41){1'b0}},Qcnt_one_47};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b110000:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-42){1'b0}},Qcnt_one_48};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b110001:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-43){1'b0}},Qcnt_one_49};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b110010:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-44){1'b0}},Qcnt_one_50};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b110011:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-45){1'b0}},Qcnt_one_51};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b110100:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-46){1'b0}},Qcnt_one_52};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b110101:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-47){1'b0}},Qcnt_one_53};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b110110:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-48){1'b0}},Qcnt_one_54};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b110111:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-49){1'b0}},Qcnt_one_55};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          6'b111000:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-50){1'b0}},Qcnt_one_56};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
            end
          default:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0='0;
              Sqrt_Q0='0;
            end
        endcase
      end
   
   
   
    2'b01:
      begin
   
   
   
        case(Crtl_cnt_S)
          6'b000000:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64+1:C_MANT_FP64];
              Q_sqrt0={{(C_MANT_FP64+5){1'b0}},Qcnt_two_0[1]};
              Sqrt_Q0=Q_sqrt_com_0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-1:C_MANT_FP64-2];
              Q_sqrt1={{(C_MANT_FP64+4){1'b0}},Qcnt_two_0[1:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b000001:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-3:C_MANT_FP64-4];
              Q_sqrt0={{(C_MANT_FP64+4){1'b0}},Qcnt_two_1[2:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-5:C_MANT_FP64-6];
              Q_sqrt1={{(C_MANT_FP64+3){1'b0}},Qcnt_two_1[2:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b000010:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-7:C_MANT_FP64-8];
              Q_sqrt0={{(C_MANT_FP64+2){1'b0}},Qcnt_two_2[4:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-9:C_MANT_FP64-10];
              Q_sqrt1={{(C_MANT_FP64+1){1'b0}},Qcnt_two_2[4:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b000011:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-11:C_MANT_FP64-12];
              Q_sqrt0={{(C_MANT_FP64){1'b0}},Qcnt_two_3[6:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-13:C_MANT_FP64-14];
              Q_sqrt1={{(C_MANT_FP64-1){1'b0}},Qcnt_two_3[6:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b000100:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-15:C_MANT_FP64-16];
              Q_sqrt0={{(C_MANT_FP64-2){1'b0}},Qcnt_two_4[8:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-17:C_MANT_FP64-18];
              Q_sqrt1={{(C_MANT_FP64-3){1'b0}},Qcnt_two_4[8:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
            6'b000101:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-19:C_MANT_FP64-20];
              Q_sqrt0={{(C_MANT_FP64-4){1'b0}},Qcnt_two_5[10:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-21:C_MANT_FP64-22];
              Q_sqrt1={{(C_MANT_FP64-5){1'b0}},Qcnt_two_5[10:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b000110:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-23:C_MANT_FP64-24];
              Q_sqrt0={{(C_MANT_FP64-6){1'b0}},Qcnt_two_6[12:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-25:C_MANT_FP64-26];
              Q_sqrt1={{(C_MANT_FP64-7){1'b0}},Qcnt_two_6[12:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b000111:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-27:C_MANT_FP64-28];
              Q_sqrt0={{(C_MANT_FP64-8){1'b0}},Qcnt_two_7[14:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-29:C_MANT_FP64-30];
              Q_sqrt1={{(C_MANT_FP64-9){1'b0}},Qcnt_two_7[14:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b001000:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-31:C_MANT_FP64-32];
              Q_sqrt0={{(C_MANT_FP64-10){1'b0}},Qcnt_two_8[16:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-33:C_MANT_FP64-34];
              Q_sqrt1={{(C_MANT_FP64-11){1'b0}},Qcnt_two_8[16:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b001001:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-35:C_MANT_FP64-36];
              Q_sqrt0={{(C_MANT_FP64-12){1'b0}},Qcnt_two_9[18:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-37:C_MANT_FP64-38];
              Q_sqrt1={{(C_MANT_FP64-13){1'b0}},Qcnt_two_9[18:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b001010:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-39:C_MANT_FP64-40];
              Q_sqrt0={{(C_MANT_FP64-14){1'b0}},Qcnt_two_10[20:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-41:C_MANT_FP64-42];
              Q_sqrt1={{(C_MANT_FP64-15){1'b0}},Qcnt_two_10[20:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b001011:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-43:C_MANT_FP64-44];
              Q_sqrt0={{(C_MANT_FP64-16){1'b0}},Qcnt_two_11[22:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-45:C_MANT_FP64-46];
              Q_sqrt1={{(C_MANT_FP64-17){1'b0}},Qcnt_two_11[22:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b001100:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-47:C_MANT_FP64-48];
              Q_sqrt0={{(C_MANT_FP64-18){1'b0}},Qcnt_two_12[24:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-49:C_MANT_FP64-50];
              Q_sqrt1={{(C_MANT_FP64-19){1'b0}},Qcnt_two_12[24:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b001101:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-51:C_MANT_FP64-52];
              Q_sqrt0={{(C_MANT_FP64-20){1'b0}},Qcnt_two_13[26:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-21){1'b0}},Qcnt_two_13[26:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b001110:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-22){1'b0}},Qcnt_two_14[28:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-23){1'b0}},Qcnt_two_14[28:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b001111:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-24){1'b0}},Qcnt_two_15[30:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-25){1'b0}},Qcnt_two_15[30:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b010000:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-26){1'b0}},Qcnt_two_16[32:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-27){1'b0}},Qcnt_two_16[32:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b010001:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-28){1'b0}},Qcnt_two_17[34:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-29){1'b0}},Qcnt_two_17[34:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b010010:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-30){1'b0}},Qcnt_two_18[36:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-31){1'b0}},Qcnt_two_18[36:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b010011:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-32){1'b0}},Qcnt_two_19[38:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-33){1'b0}},Qcnt_two_19[38:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b010100:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-34){1'b0}},Qcnt_two_20[40:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-35){1'b0}},Qcnt_two_20[40:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b010101:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-36){1'b0}},Qcnt_two_21[42:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-37){1'b0}},Qcnt_two_21[42:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b010110:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-38){1'b0}},Qcnt_two_22[44:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-39){1'b0}},Qcnt_two_22[44:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b010111:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-40){1'b0}},Qcnt_two_23[46:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-41){1'b0}},Qcnt_two_23[46:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b011000:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-42){1'b0}},Qcnt_two_24[48:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-43){1'b0}},Qcnt_two_24[48:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b011001:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-44){1'b0}},Qcnt_two_25[50:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-45){1'b0}},Qcnt_two_25[50:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b011010:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-46){1'b0}},Qcnt_two_26[52:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-47){1'b0}},Qcnt_two_26[52:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b011011:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-48){1'b0}},Qcnt_two_27[54:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-49){1'b0}},Qcnt_two_27[54:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          6'b011100:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-50){1'b0}},Qcnt_two_28[56:1]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-51){1'b0}},Qcnt_two_28[56:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
          default:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64+1:C_MANT_FP64];
              Q_sqrt0={{(C_MANT_FP64+5){1'b0}},Qcnt_two_0[1]};
              Sqrt_Q0=Q_sqrt_com_0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-1:C_MANT_FP64-2];
              Q_sqrt1={{(C_MANT_FP64+4){1'b0}},Qcnt_two_0[1:0]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
            end
        endcase
      end
   
   
   
    2'b10:
      begin
   
   
   
        case(Crtl_cnt_S)
          6'b000000:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64+1:C_MANT_FP64];
              Q_sqrt0={{(C_MANT_FP64+5){1'b0}},Qcnt_three_0[2]};
              Sqrt_Q0=Q_sqrt_com_0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-1:C_MANT_FP64-2];
              Q_sqrt1={{(C_MANT_FP64+4){1'b0}},Qcnt_three_0[2:1]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
              Sqrt_DI[2]=Mant_D_sqrt_Norm[C_MANT_FP64-3:C_MANT_FP64-4];
              Q_sqrt2={{(C_MANT_FP64+3){1'b0}},Qcnt_three_0[2:0]};
              Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
            end
          6'b000001:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-5:C_MANT_FP64-6];
              Q_sqrt0={{(C_MANT_FP64+2){1'b0}},Qcnt_three_1[4:2]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-7:C_MANT_FP64-8];
              Q_sqrt1={{(C_MANT_FP64+1){1'b0}},Qcnt_three_1[4:1]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
              Sqrt_DI[2]=Mant_D_sqrt_Norm[C_MANT_FP64-9:C_MANT_FP64-10];
              Q_sqrt2={{(C_MANT_FP64){1'b0}},Qcnt_three_1[4:0]};
              Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
            end
          6'b000010:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-11:C_MANT_FP64-12];
              Q_sqrt0={{(C_MANT_FP64-1){1'b0}},Qcnt_three_2[7:2]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-13:C_MANT_FP64-14];
              Q_sqrt1={{(C_MANT_FP64-2){1'b0}},Qcnt_three_2[7:1]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
              Sqrt_DI[2]=Mant_D_sqrt_Norm[C_MANT_FP64-15:C_MANT_FP64-16];
              Q_sqrt2={{(C_MANT_FP64-3){1'b0}},Qcnt_three_2[7:0]};
              Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
            end
          6'b000011:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-17:C_MANT_FP64-18];
              Q_sqrt0={{(C_MANT_FP64-4){1'b0}},Qcnt_three_3[10:2]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-19:C_MANT_FP64-20];
              Q_sqrt1={{(C_MANT_FP64-5){1'b0}},Qcnt_three_3[10:1]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
              Sqrt_DI[2]=Mant_D_sqrt_Norm[C_MANT_FP64-21:C_MANT_FP64-22];
              Q_sqrt2={{(C_MANT_FP64-6){1'b0}},Qcnt_three_3[10:0]};
              Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
            end
          6'b000100:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-23:C_MANT_FP64-24];
              Q_sqrt0={{(C_MANT_FP64-7){1'b0}},Qcnt_three_4[13:2]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-25:C_MANT_FP64-26];
              Q_sqrt1={{(C_MANT_FP64-8){1'b0}},Qcnt_three_4[13:1]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
              Sqrt_DI[2]=Mant_D_sqrt_Norm[C_MANT_FP64-27:C_MANT_FP64-28];
              Q_sqrt2={{(C_MANT_FP64-9){1'b0}},Qcnt_three_4[13:0]};
              Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
            end
          6'b000101:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-29:C_MANT_FP64-30];
              Q_sqrt0={{(C_MANT_FP64-10){1'b0}},Qcnt_three_5[16:2]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-31:C_MANT_FP64-32];
              Q_sqrt1={{(C_MANT_FP64-11){1'b0}},Qcnt_three_5[16:1]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
              Sqrt_DI[2]=Mant_D_sqrt_Norm[C_MANT_FP64-33:C_MANT_FP64-34];
              Q_sqrt2={{(C_MANT_FP64-12){1'b0}},Qcnt_three_5[16:0]};
              Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
            end
          6'b000110:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-35:C_MANT_FP64-36];
              Q_sqrt0={{(C_MANT_FP64-13){1'b0}},Qcnt_three_6[19:2]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-37:C_MANT_FP64-38];
              Q_sqrt1={{(C_MANT_FP64-14){1'b0}},Qcnt_three_6[19:1]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
              Sqrt_DI[2]=Mant_D_sqrt_Norm[C_MANT_FP64-39:C_MANT_FP64-40];
              Q_sqrt2={{(C_MANT_FP64-15){1'b0}},Qcnt_three_6[19:0]};
              Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
            end
          6'b000111:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-41:C_MANT_FP64-42];
              Q_sqrt0={{(C_MANT_FP64-16){1'b0}},Qcnt_three_7[22:2]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-43:C_MANT_FP64-44];
              Q_sqrt1={{(C_MANT_FP64-17){1'b0}},Qcnt_three_7[22:1]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
              Sqrt_DI[2]=Mant_D_sqrt_Norm[C_MANT_FP64-45:C_MANT_FP64-46];
              Q_sqrt2={{(C_MANT_FP64-18){1'b0}},Qcnt_three_7[22:0]};
              Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
            end
          6'b001000:
            begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-47:C_MANT_FP64-48];
              Q_sqrt0={{(C_MANT_FP64-19){1'b0}},Qcnt_three_8[25:2]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-49:C_MANT_FP64-50];
              Q_sqrt1={{(C_MANT_FP64-20){1'b0}},Qcnt_three_8[25:1]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
              Sqrt_DI[2]=Mant_D_sqrt_Norm[C_MANT_FP64-51:C_MANT_FP64-52];
              Q_sqrt2={{(C_MANT_FP64-21){1'b0}},Qcnt_three_8[25:0]};
              Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
            end
          6'b001001:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-22){1'b0}},Qcnt_three_9[28:2]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-23){1'b0}},Qcnt_three_9[28:1]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
              Sqrt_DI[2]=2'b00;
              Q_sqrt2={{(C_MANT_FP64-24){1'b0}},Qcnt_three_9[28:0]};
              Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
            end
          6'b001010:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-25){1'b0}},Qcnt_three_10[31:2]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-26){1'b0}},Qcnt_three_10[31:1]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
              Sqrt_DI[2]=2'b00;
              Q_sqrt2={{(C_MANT_FP64-27){1'b0}},Qcnt_three_10[31:0]};
              Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
            end
          6'b001011:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-28){1'b0}},Qcnt_three_11[34:2]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-29){1'b0}},Qcnt_three_11[34:1]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
              Sqrt_DI[2]=2'b00;
              Q_sqrt2={{(C_MANT_FP64-30){1'b0}},Qcnt_three_11[34:0]};
              Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
            end
          6'b001100:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-31){1'b0}},Qcnt_three_12[37:2]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-32){1'b0}},Qcnt_three_12[37:1]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
              Sqrt_DI[2]=2'b00;
              Q_sqrt2={{(C_MANT_FP64-33){1'b0}},Qcnt_three_12[37:0]};
              Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
            end
          6'b001101:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-34){1'b0}},Qcnt_three_13[40:2]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-35){1'b0}},Qcnt_three_13[40:1]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
              Sqrt_DI[2]=2'b00;
              Q_sqrt2={{(C_MANT_FP64-36){1'b0}},Qcnt_three_13[40:0]};
              Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
            end
          6'b001110:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-37){1'b0}},Qcnt_three_14[43:2]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-38){1'b0}},Qcnt_three_14[43:1]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
              Sqrt_DI[2]=2'b00;
              Q_sqrt2={{(C_MANT_FP64-39){1'b0}},Qcnt_three_14[43:0]};
              Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
            end
          6'b001111:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-40){1'b0}},Qcnt_three_15[46:2]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-41){1'b0}},Qcnt_three_15[46:1]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
              Sqrt_DI[2]=2'b00;
              Q_sqrt2={{(C_MANT_FP64-42){1'b0}},Qcnt_three_15[46:0]};
              Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
            end
          6'b010000:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-43){1'b0}},Qcnt_three_16[49:2]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-44){1'b0}},Qcnt_three_16[49:1]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
              Sqrt_DI[2]=2'b00;
              Q_sqrt2={{(C_MANT_FP64-45){1'b0}},Qcnt_three_16[49:0]};
              Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
            end
          6'b010001:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-46){1'b0}},Qcnt_three_17[52:2]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-47){1'b0}},Qcnt_three_17[52:1]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
              Sqrt_DI[2]=2'b00;
              Q_sqrt2={{(C_MANT_FP64-48){1'b0}},Qcnt_three_17[52:0]};
              Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
            end
          6'b010010:
            begin
              Sqrt_DI[0]=2'b00;
              Q_sqrt0={{(C_MANT_FP64-49){1'b0}},Qcnt_three_18[55:2]};
              Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
              Sqrt_DI[1]=2'b00;
              Q_sqrt1={{(C_MANT_FP64-50){1'b0}},Qcnt_three_18[55:1]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
              Sqrt_DI[2]=2'b00;
              Q_sqrt2={{(C_MANT_FP64-51){1'b0}},Qcnt_three_18[55:0]};
              Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
            end
          default :
              begin
              Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64+1:C_MANT_FP64];
              Q_sqrt0={{(C_MANT_FP64+5){1'b0}},Qcnt_three_0[2]};
              Sqrt_Q0=Q_sqrt_com_0;
              Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-1:C_MANT_FP64-2];
              Q_sqrt1={{(C_MANT_FP64+4){1'b0}},Qcnt_three_0[2:1]};
              Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
              Sqrt_DI[2]=Mant_D_sqrt_Norm[C_MANT_FP64-3:C_MANT_FP64-4];
              Q_sqrt2={{(C_MANT_FP64+3){1'b0}},Qcnt_three_0[2:0]};
              Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
            end
        endcase
      end
   
   
   
    2'b11:
      begin
   
   
   
              case(Crtl_cnt_S)
                6'b000000:
                  begin
                    Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64+1:C_MANT_FP64];
                    Q_sqrt0={{(C_MANT_FP64+5){1'b0}},Qcnt_four_0[3]};
                    Sqrt_Q0=Q_sqrt_com_0;
                    Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-1:C_MANT_FP64-2];
                    Q_sqrt1={{(C_MANT_FP64+4){1'b0}},Qcnt_four_0[3:2]};
                    Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
                    Sqrt_DI[2]=Mant_D_sqrt_Norm[C_MANT_FP64-3:C_MANT_FP64-4];
                    Q_sqrt2={{(C_MANT_FP64+3){1'b0}},Qcnt_four_0[3:1]};
                    Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
                    Sqrt_DI[3]=Mant_D_sqrt_Norm[C_MANT_FP64-5:C_MANT_FP64-6];
                    Q_sqrt3={{(C_MANT_FP64+2){1'b0}},Qcnt_four_0[3:0]};
                    Sqrt_Q3=Sqrt_quotinent_S[1]?Q_sqrt_com_3:Q_sqrt3;
                  end
                6'b000001:
                  begin
                    Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-7:C_MANT_FP64-8];
                    Q_sqrt0={{(C_MANT_FP64+1){1'b0}},Qcnt_four_1[6:3]};
                    Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
                    Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-9:C_MANT_FP64-10];
                    Q_sqrt1={{(C_MANT_FP64){1'b0}},Qcnt_four_1[6:2]};
                    Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
                    Sqrt_DI[2]=Mant_D_sqrt_Norm[C_MANT_FP64-11:C_MANT_FP64-12];
                    Q_sqrt2={{(C_MANT_FP64-1){1'b0}},Qcnt_four_1[6:1]};
                    Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
                    Sqrt_DI[3]=Mant_D_sqrt_Norm[C_MANT_FP64-13:C_MANT_FP64-14];
                    Q_sqrt3={{(C_MANT_FP64-2){1'b0}},Qcnt_four_1[6:0]};
                    Sqrt_Q3=Sqrt_quotinent_S[1]?Q_sqrt_com_3:Q_sqrt3;
                  end
                6'b000010:
                  begin
                    Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-15:C_MANT_FP64-16];
                    Q_sqrt0={{(C_MANT_FP64-3){1'b0}},Qcnt_four_2[10:3]};
                    Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
                    Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-17:C_MANT_FP64-18];
                    Q_sqrt1={{(C_MANT_FP64-4){1'b0}},Qcnt_four_2[10:2]};
                    Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
                    Sqrt_DI[2]=Mant_D_sqrt_Norm[C_MANT_FP64-19:C_MANT_FP64-20];
                    Q_sqrt2={{(C_MANT_FP64-5){1'b0}},Qcnt_four_2[10:1]};
                    Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
                    Sqrt_DI[3]=Mant_D_sqrt_Norm[C_MANT_FP64-21:C_MANT_FP64-22];
                    Q_sqrt3={{(C_MANT_FP64-6){1'b0}},Qcnt_four_2[10:0]};
                    Sqrt_Q3=Sqrt_quotinent_S[1]?Q_sqrt_com_3:Q_sqrt3;
                  end
                6'b000011:
                  begin
                    Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-23:C_MANT_FP64-24];
                    Q_sqrt0={{(C_MANT_FP64-7){1'b0}},Qcnt_four_3[14:3]};
                    Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
                    Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-25:C_MANT_FP64-26];
                    Q_sqrt1={{(C_MANT_FP64-8){1'b0}},Qcnt_four_3[14:2]};
                    Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
                    Sqrt_DI[2]=Mant_D_sqrt_Norm[C_MANT_FP64-27:C_MANT_FP64-28];
                    Q_sqrt2={{(C_MANT_FP64-9){1'b0}},Qcnt_four_3[14:1]};
                    Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
                    Sqrt_DI[3]=Mant_D_sqrt_Norm[C_MANT_FP64-29:C_MANT_FP64-30];
                    Q_sqrt3={{(C_MANT_FP64-10){1'b0}},Qcnt_four_3[14:0]};
                    Sqrt_Q3=Sqrt_quotinent_S[1]?Q_sqrt_com_3:Q_sqrt3;
                  end
                6'b000100:
                  begin
                    Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-31:C_MANT_FP64-32];
                    Q_sqrt0={{(C_MANT_FP64-11){1'b0}},Qcnt_four_4[18:3]};
                    Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
                    Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-33:C_MANT_FP64-34];
                    Q_sqrt1={{(C_MANT_FP64-12){1'b0}},Qcnt_four_4[18:2]};
                    Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
                    Sqrt_DI[2]=Mant_D_sqrt_Norm[C_MANT_FP64-35:C_MANT_FP64-36];
                    Q_sqrt2={{(C_MANT_FP64-13){1'b0}},Qcnt_four_4[18:1]};
                    Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
                    Sqrt_DI[3]=Mant_D_sqrt_Norm[C_MANT_FP64-37:C_MANT_FP64-38];
                    Q_sqrt3={{(C_MANT_FP64-14){1'b0}},Qcnt_four_4[18:0]};
                    Sqrt_Q3=Sqrt_quotinent_S[1]?Q_sqrt_com_3:Q_sqrt3;
                  end
                6'b000101:
                  begin
                    Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-39:C_MANT_FP64-40];
                    Q_sqrt0={{(C_MANT_FP64-15){1'b0}},Qcnt_four_5[22:3]};
                    Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
                    Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-41:C_MANT_FP64-42];
                    Q_sqrt1={{(C_MANT_FP64-16){1'b0}},Qcnt_four_5[22:2]};
                    Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
                    Sqrt_DI[2]=Mant_D_sqrt_Norm[C_MANT_FP64-43:C_MANT_FP64-44];
                    Q_sqrt2={{(C_MANT_FP64-17){1'b0}},Qcnt_four_5[22:1]};
                    Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
                    Sqrt_DI[3]=Mant_D_sqrt_Norm[C_MANT_FP64-45:C_MANT_FP64-46];
                    Q_sqrt3={{(C_MANT_FP64-18){1'b0}},Qcnt_four_5[22:0]};
                    Sqrt_Q3=Sqrt_quotinent_S[1]?Q_sqrt_com_3:Q_sqrt3;
                  end
                6'b000110:
                  begin
                    Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64-47:C_MANT_FP64-48];
                    Q_sqrt0={{(C_MANT_FP64-19){1'b0}},Qcnt_four_6[26:3]};
                    Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
                    Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-49:C_MANT_FP64-50];
                    Q_sqrt1={{(C_MANT_FP64-20){1'b0}},Qcnt_four_6[26:2]};
                    Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
                    Sqrt_DI[2]=Mant_D_sqrt_Norm[C_MANT_FP64-51:C_MANT_FP64-52];
                    Q_sqrt2={{(C_MANT_FP64-21){1'b0}},Qcnt_four_6[26:1]};
                    Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
                    Sqrt_DI[3]=2'b00;
                    Q_sqrt3={{(C_MANT_FP64-22){1'b0}},Qcnt_four_6[26:0]};
                    Sqrt_Q3=Sqrt_quotinent_S[1]?Q_sqrt_com_3:Q_sqrt3;
                  end
                6'b000111:
                  begin
                    Sqrt_DI[0]=2'b00;
                    Q_sqrt0={{(C_MANT_FP64-23){1'b0}},Qcnt_four_7[30:3]};
                    Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
                    Sqrt_DI[1]=2'b00;
                    Q_sqrt1={{(C_MANT_FP64-24){1'b0}},Qcnt_four_7[30:2]};
                    Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
                    Sqrt_DI[2]=2'b00;
                    Q_sqrt2={{(C_MANT_FP64-25){1'b0}},Qcnt_four_7[30:1]};
                    Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
                    Sqrt_DI[3]=2'b00;
                    Q_sqrt3={{(C_MANT_FP64-26){1'b0}},Qcnt_four_7[30:0]};
                    Sqrt_Q3=Sqrt_quotinent_S[1]?Q_sqrt_com_3:Q_sqrt3;
                  end
                6'b001000:
                  begin
                    Sqrt_DI[0]=2'b00;
                    Q_sqrt0={{(C_MANT_FP64-27){1'b0}},Qcnt_four_8[34:3]};
                    Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
                    Sqrt_DI[1]=2'b00;
                    Q_sqrt1={{(C_MANT_FP64-28){1'b0}},Qcnt_four_8[34:2]};
                    Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
                    Sqrt_DI[2]=2'b00;
                    Q_sqrt2={{(C_MANT_FP64-29){1'b0}},Qcnt_four_8[34:1]};
                    Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
                    Sqrt_DI[3]=2'b00;
                    Q_sqrt3={{(C_MANT_FP64-30){1'b0}},Qcnt_four_8[34:0]};
                    Sqrt_Q3=Sqrt_quotinent_S[1]?Q_sqrt_com_3:Q_sqrt3;
                  end
                6'b001001:
                  begin
                    Sqrt_DI[0]=2'b00;
                    Q_sqrt0={{(C_MANT_FP64-31){1'b0}},Qcnt_four_9[38:3]};
                    Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
                    Sqrt_DI[1]=2'b00;
                    Q_sqrt1={{(C_MANT_FP64-32){1'b0}},Qcnt_four_9[38:2]};
                    Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
                    Sqrt_DI[2]=2'b00;
                    Q_sqrt2={{(C_MANT_FP64-33){1'b0}},Qcnt_four_9[38:1]};
                    Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
                    Sqrt_DI[3]=2'b00;
                    Q_sqrt3={{(C_MANT_FP64-34){1'b0}},Qcnt_four_9[38:0]};
                    Sqrt_Q3=Sqrt_quotinent_S[1]?Q_sqrt_com_3:Q_sqrt3;
                  end
                6'b001010:
                  begin
                    Sqrt_DI[0]=2'b00;
                    Q_sqrt0={{(C_MANT_FP64-35){1'b0}},Qcnt_four_10[42:3]};
                    Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
                    Sqrt_DI[1]=2'b00;
                    Q_sqrt1={{(C_MANT_FP64-36){1'b0}},Qcnt_four_10[42:2]};
                    Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
                    Sqrt_DI[2]=2'b00;
                    Q_sqrt2={{(C_MANT_FP64-37){1'b0}},Qcnt_four_10[42:1]};
                    Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
                    Sqrt_DI[3]=2'b00;
                    Q_sqrt3={{(C_MANT_FP64-38){1'b0}},Qcnt_four_10[42:0]};
                    Sqrt_Q3=Sqrt_quotinent_S[1]?Q_sqrt_com_3:Q_sqrt3;
                  end
                6'b001011:
                  begin
                    Sqrt_DI[0]=2'b00;
                    Q_sqrt0={{(C_MANT_FP64-39){1'b0}},Qcnt_four_11[46:3]};
                    Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
                    Sqrt_DI[1]=2'b00;
                    Q_sqrt1={{(C_MANT_FP64-40){1'b0}},Qcnt_four_11[46:2]};
                    Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
                    Sqrt_DI[2]=2'b00;
                    Q_sqrt2={{(C_MANT_FP64-41){1'b0}},Qcnt_four_11[46:1]};
                    Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
                    Sqrt_DI[3]=2'b00;
                    Q_sqrt3={{(C_MANT_FP64-42){1'b0}},Qcnt_four_11[46:0]};
                    Sqrt_Q3=Sqrt_quotinent_S[1]?Q_sqrt_com_3:Q_sqrt3;
                  end
                6'b001100:
                  begin
                    Sqrt_DI[0]=2'b00;
                    Q_sqrt0={{(C_MANT_FP64-43){1'b0}},Qcnt_four_12[50:3]};
                    Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
                    Sqrt_DI[1]=2'b00;
                    Q_sqrt1={{(C_MANT_FP64-44){1'b0}},Qcnt_four_12[50:2]};
                    Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
                    Sqrt_DI[2]=2'b00;
                    Q_sqrt2={{(C_MANT_FP64-45){1'b0}},Qcnt_four_12[50:1]};
                    Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
                    Sqrt_DI[3]=2'b00;
                    Q_sqrt3={{(C_MANT_FP64-46){1'b0}},Qcnt_four_12[50:0]};
                    Sqrt_Q3=Sqrt_quotinent_S[1]?Q_sqrt_com_3:Q_sqrt3;
                  end
                6'b001101:
                  begin
                    Sqrt_DI[0]=2'b00;
                    Q_sqrt0={{(C_MANT_FP64-47){1'b0}},Qcnt_four_13[54:3]};
                    Sqrt_Q0=Quotient_DP[0]?Q_sqrt_com_0:Q_sqrt0;
                    Sqrt_DI[1]=2'b00;
                    Q_sqrt1={{(C_MANT_FP64-48){1'b0}},Qcnt_four_13[54:2]};
                    Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
                    Sqrt_DI[2]=2'b00;
                    Q_sqrt2={{(C_MANT_FP64-49){1'b0}},Qcnt_four_13[54:1]};
                    Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
                    Sqrt_DI[3]=2'b00;
                    Q_sqrt3={{(C_MANT_FP64-50){1'b0}},Qcnt_four_13[54:0]};
                    Sqrt_Q3=Sqrt_quotinent_S[1]?Q_sqrt_com_3:Q_sqrt3;
                  end
                default:
                  begin
                    Sqrt_DI[0]=Mant_D_sqrt_Norm[C_MANT_FP64+1:C_MANT_FP64];
                    Q_sqrt0={{(C_MANT_FP64+5){1'b0}},Qcnt_four_0[3]};
                    Sqrt_Q0=Q_sqrt_com_0;
                    Sqrt_DI[1]=Mant_D_sqrt_Norm[C_MANT_FP64-1:C_MANT_FP64-2];
                    Q_sqrt1={{(C_MANT_FP64+4){1'b0}},Qcnt_four_0[3:2]};
                    Sqrt_Q1=Sqrt_quotinent_S[3]?Q_sqrt_com_1:Q_sqrt1;
                    Sqrt_DI[2]=Mant_D_sqrt_Norm[C_MANT_FP64-3:C_MANT_FP64-4];
                    Q_sqrt2={{(C_MANT_FP64+3){1'b0}},Qcnt_four_0[3:1]};
                    Sqrt_Q2=Sqrt_quotinent_S[2]?Q_sqrt_com_2:Q_sqrt2;
                    Sqrt_DI[3]=Mant_D_sqrt_Norm[C_MANT_FP64-5:C_MANT_FP64-6];
                    Q_sqrt3={{(C_MANT_FP64+2){1'b0}},Qcnt_four_0[3:0]};
                    Sqrt_Q3=Sqrt_quotinent_S[1]?Q_sqrt_com_3:Q_sqrt3;
                  end
              endcase
            end
      endcase
   
   
   
 end
  assign Sqrt_R0= ((Sqrt_start_dly_S)?'0:{Partial_remainder_DP[C_MANT_FP64+5:0]});
  assign Sqrt_R1= {Iteration_cell_sum_AMASK_D[0][C_MANT_FP64+5],Iteration_cell_sum_AMASK_D[0][C_MANT_FP64+2:0],Sqrt_DO[0]} ;
  assign Sqrt_R2= {Iteration_cell_sum_AMASK_D[1][C_MANT_FP64+5],Iteration_cell_sum_AMASK_D[1][C_MANT_FP64+2:0],Sqrt_DO[1]};
  assign Sqrt_R3= {Iteration_cell_sum_AMASK_D[2][C_MANT_FP64+5],Iteration_cell_sum_AMASK_D[2][C_MANT_FP64+2:0],Sqrt_DO[2]};
  assign Sqrt_R4= {Iteration_cell_sum_AMASK_D[3][C_MANT_FP64+5],Iteration_cell_sum_AMASK_D[3][C_MANT_FP64+2:0],Sqrt_DO[3]};
  logic [C_MANT_FP64+5:0]                               Denominator_se_format_DB;  
  assign Denominator_se_format_DB={Denominator_se_DB[C_MANT_FP64+1:C_MANT_FP64-C_MANT_FP16ALT],{FP16ALT_SO?FP16ALT_SO:Denominator_se_DB[C_MANT_FP64-C_MANT_FP16ALT-1]},
                                                         Denominator_se_DB[C_MANT_FP64-C_MANT_FP16ALT-2:C_MANT_FP64-C_MANT_FP16],{FP16_SO?FP16_SO:Denominator_se_DB[C_MANT_FP64-C_MANT_FP16-1]},
                                                         Denominator_se_DB[C_MANT_FP64-C_MANT_FP16-2:C_MANT_FP64-C_MANT_FP32],{FP32_SO?FP32_SO:Denominator_se_DB[C_MANT_FP64-C_MANT_FP32-1]},
                                                         Denominator_se_DB[C_MANT_FP64-C_MANT_FP32-2:C_MANT_FP64-C_MANT_FP64],FP64_SO,3'b0} ;
  
  logic [C_MANT_FP64+5:0]                           First_iteration_cell_div_a_D,First_iteration_cell_div_b_D;
  logic                                             Sel_b_for_first_S;
  assign First_iteration_cell_div_a_D=(Div_start_dly_S)?{Numerator_se_D[C_MANT_FP64+1:C_MANT_FP64-C_MANT_FP16ALT],{FP16ALT_SO?FP16ALT_SO:Numerator_se_D[C_MANT_FP64-C_MANT_FP16ALT-1]},
                                                         Numerator_se_D[C_MANT_FP64-C_MANT_FP16ALT-2:C_MANT_FP64-C_MANT_FP16],{FP16_SO?FP16_SO:Numerator_se_D[C_MANT_FP64-C_MANT_FP16-1]},
                                                         Numerator_se_D[C_MANT_FP64-C_MANT_FP16-2:C_MANT_FP64-C_MANT_FP32],{FP32_SO?FP32_SO:Numerator_se_D[C_MANT_FP64-C_MANT_FP32-1]},
                                                         Numerator_se_D[C_MANT_FP64-C_MANT_FP32-2:C_MANT_FP64-C_MANT_FP64],FP64_SO,3'b0}
                                                        :{Partial_remainder_DP[C_MANT_FP64+4:C_MANT_FP64-C_MANT_FP16ALT+3],{FP16ALT_SO?Quotient_DP[0]:Partial_remainder_DP[C_MANT_FP64-C_MANT_FP16ALT+2]},
                                                         Partial_remainder_DP[C_MANT_FP64-C_MANT_FP16ALT+1:C_MANT_FP64-C_MANT_FP16+3],{FP16_SO?Quotient_DP[0]:Partial_remainder_DP[C_MANT_FP64-C_MANT_FP16+2]},
                                                         Partial_remainder_DP[C_MANT_FP64-C_MANT_FP16+1:C_MANT_FP64-C_MANT_FP32+3],{FP32_SO?Quotient_DP[0]:Partial_remainder_DP[C_MANT_FP64-C_MANT_FP32+2]},
                                                         Partial_remainder_DP[C_MANT_FP64-C_MANT_FP32+1:C_MANT_FP64-C_MANT_FP64+3],FP64_SO&&Quotient_DP[0],3'b0};
  assign Sel_b_for_first_S=(Div_start_dly_S)?1:Quotient_DP[0];
  assign First_iteration_cell_div_b_D=Sel_b_for_first_S?Denominator_se_format_DB:{Denominator_se_D,4'b0};
  assign Iteration_cell_a_BMASK_D[0]=Sqrt_enable_SO?Sqrt_R0:{First_iteration_cell_div_a_D};
  assign Iteration_cell_b_BMASK_D[0]=Sqrt_enable_SO?Sqrt_Q0:{First_iteration_cell_div_b_D};
  
  logic [C_MANT_FP64+5:0]                          Sec_iteration_cell_div_a_D,Sec_iteration_cell_div_b_D;
  logic                                            Sel_b_for_sec_S;
  generate
    if(|Iteration_unit_num_S)
      begin
        assign Sel_b_for_sec_S=~Iteration_cell_sum_AMASK_D[0][C_MANT_FP64+5];
        assign Sec_iteration_cell_div_a_D={Iteration_cell_sum_AMASK_D[0][C_MANT_FP64+4:C_MANT_FP64-C_MANT_FP16ALT+3],{FP16ALT_SO?Sel_b_for_sec_S:Iteration_cell_sum_AMASK_D[0][C_MANT_FP64-C_MANT_FP16ALT+2]},
                                           Iteration_cell_sum_AMASK_D[0][C_MANT_FP64-C_MANT_FP16ALT+1:C_MANT_FP64-C_MANT_FP16+3],{FP16_SO?Sel_b_for_sec_S:Iteration_cell_sum_AMASK_D[0][C_MANT_FP64-C_MANT_FP16+2]},
                                           Iteration_cell_sum_AMASK_D[0][C_MANT_FP64-C_MANT_FP16+1:C_MANT_FP64-C_MANT_FP32+3],{FP32_SO?Sel_b_for_sec_S:Iteration_cell_sum_AMASK_D[0][C_MANT_FP64-C_MANT_FP32+2]},
                                           Iteration_cell_sum_AMASK_D[0][C_MANT_FP64-C_MANT_FP32+1:C_MANT_FP64-C_MANT_FP64+3],FP64_SO&&Sel_b_for_sec_S,3'b0};
        assign Sec_iteration_cell_div_b_D=Sel_b_for_sec_S?Denominator_se_format_DB:{Denominator_se_D,4'b0};
        assign Iteration_cell_a_BMASK_D[1]=Sqrt_enable_SO?Sqrt_R1:{Sec_iteration_cell_div_a_D};
        assign Iteration_cell_b_BMASK_D[1]=Sqrt_enable_SO?Sqrt_Q1:{Sec_iteration_cell_div_b_D};
      end
    endgenerate
  
  logic [C_MANT_FP64+5:0]                          Thi_iteration_cell_div_a_D,Thi_iteration_cell_div_b_D;
  logic                                            Sel_b_for_thi_S;
  generate
    if((Iteration_unit_num_S==2'b10) | (Iteration_unit_num_S==2'b11))
      begin
        assign Sel_b_for_thi_S=~Iteration_cell_sum_AMASK_D[1][C_MANT_FP64+5];
        assign Thi_iteration_cell_div_a_D={Iteration_cell_sum_AMASK_D[1][C_MANT_FP64+4:C_MANT_FP64-C_MANT_FP16ALT+3],{FP16ALT_SO?Sel_b_for_thi_S:Iteration_cell_sum_AMASK_D[1][C_MANT_FP64-C_MANT_FP16ALT+2]},
                                           Iteration_cell_sum_AMASK_D[1][C_MANT_FP64-C_MANT_FP16ALT+1:C_MANT_FP64-C_MANT_FP16+3],{FP16_SO?Sel_b_for_thi_S:Iteration_cell_sum_AMASK_D[1][C_MANT_FP64-C_MANT_FP16+2]},
                                           Iteration_cell_sum_AMASK_D[1][C_MANT_FP64-C_MANT_FP16+1:C_MANT_FP64-C_MANT_FP32+3],{FP32_SO?Sel_b_for_thi_S:Iteration_cell_sum_AMASK_D[1][C_MANT_FP64-C_MANT_FP32+2]},
                                           Iteration_cell_sum_AMASK_D[1][C_MANT_FP64-C_MANT_FP32+1:C_MANT_FP64-C_MANT_FP64+3],FP64_SO&&Sel_b_for_thi_S,3'b0};
        assign Thi_iteration_cell_div_b_D=Sel_b_for_thi_S?Denominator_se_format_DB:{Denominator_se_D,4'b0};
        assign Iteration_cell_a_BMASK_D[2]=Sqrt_enable_SO?Sqrt_R2:{Thi_iteration_cell_div_a_D};
        assign Iteration_cell_b_BMASK_D[2]=Sqrt_enable_SO?Sqrt_Q2:{Thi_iteration_cell_div_b_D};
      end
  endgenerate
  
  logic [C_MANT_FP64+5:0]                          Fou_iteration_cell_div_a_D,Fou_iteration_cell_div_b_D;
  logic                                            Sel_b_for_fou_S;
  generate
    if(Iteration_unit_num_S==2'b11)
      begin
        assign Sel_b_for_fou_S=~Iteration_cell_sum_AMASK_D[2][C_MANT_FP64+5];
        assign Fou_iteration_cell_div_a_D={Iteration_cell_sum_AMASK_D[2][C_MANT_FP64+4:C_MANT_FP64-C_MANT_FP16ALT+3],{FP16ALT_SO?Sel_b_for_fou_S:Iteration_cell_sum_AMASK_D[2][C_MANT_FP64-C_MANT_FP16ALT+2]},
                                           Iteration_cell_sum_AMASK_D[2][C_MANT_FP64-C_MANT_FP16ALT+1:C_MANT_FP64-C_MANT_FP16+3],{FP16_SO?Sel_b_for_fou_S:Iteration_cell_sum_AMASK_D[2][C_MANT_FP64-C_MANT_FP16+2]},
                                           Iteration_cell_sum_AMASK_D[2][C_MANT_FP64-C_MANT_FP16+1:C_MANT_FP64-C_MANT_FP32+3],{FP32_SO?Sel_b_for_fou_S:Iteration_cell_sum_AMASK_D[2][C_MANT_FP64-C_MANT_FP32+2]},
                                           Iteration_cell_sum_AMASK_D[2][C_MANT_FP64-C_MANT_FP32+1:C_MANT_FP64-C_MANT_FP64+3],FP64_SO&&Sel_b_for_fou_S,3'b0};
        assign Fou_iteration_cell_div_b_D=Sel_b_for_fou_S?Denominator_se_format_DB:{Denominator_se_D,4'b0};
        assign Iteration_cell_a_BMASK_D[3]=Sqrt_enable_SO?Sqrt_R3:{Fou_iteration_cell_div_a_D};
        assign Iteration_cell_b_BMASK_D[3]=Sqrt_enable_SO?Sqrt_Q3:{Fou_iteration_cell_div_b_D};
      end
  endgenerate
   
   
   
  logic [C_MANT_FP64+1+4:0]                          Mask_bits_ctl_S;  
  assign Mask_bits_ctl_S =58'h3ff_ffff_ffff_ffff;   
   
   
   
  logic                                             Div_enable_SI   [3:0];
  logic                                             Div_start_dly_SI   [3:0];
  logic                                             Sqrt_enable_SI   [3:0];
  generate
    genvar i,j;
      for (i=0; i <= Iteration_unit_num_S ; i++)
        begin
          for (j = 0; j <= C_MANT_FP64+5; j++) begin
              assign Iteration_cell_a_D[i][j] = Mask_bits_ctl_S[j] && Iteration_cell_a_BMASK_D[i][j];
              assign Iteration_cell_b_D[i][j] = Mask_bits_ctl_S[j] && Iteration_cell_b_BMASK_D[i][j];
              assign Iteration_cell_sum_AMASK_D[i][j] = Mask_bits_ctl_S[j] && Iteration_cell_sum_D[i][j];
          end
          assign  Div_enable_SI[i] = Div_enable_SO;
          assign  Div_start_dly_SI[i] = Div_start_dly_S;
          assign  Sqrt_enable_SI[i] = Sqrt_enable_SO;
          iteration_div_sqrt_mvp #(C_MANT_FP64+6) iteration_div_sqrt
          (
          .A_DI                                    (Iteration_cell_a_D[i]            ),
          .B_DI                                    (Iteration_cell_b_D[i]            ),
          .Div_enable_SI                           (Div_enable_SI[i]                 ),
          .Div_start_dly_SI                        (Div_start_dly_SI[i]              ),
          .Sqrt_enable_SI                          (Sqrt_enable_SI[i]                ),
          .D_DI                                    (Sqrt_DI[i]                       ),
          .D_DO                                    (Sqrt_DO[i]                       ),
          .Sum_DO                                  (Iteration_cell_sum_D[i]          ),
          .Carry_out_DO                            (Iteration_cell_carry_D[i]        )
         );
        end
  endgenerate
  always_comb
    begin
      case (Iteration_unit_num_S)
        2'b00:
          begin
            if(Fsm_enable_S)
               Partial_remainder_DN = Sqrt_enable_SO?Sqrt_R1:Iteration_cell_sum_AMASK_D[0];
            else
               Partial_remainder_DN = Partial_remainder_DP;
          end
        2'b01:
          begin
            if(Fsm_enable_S)
               Partial_remainder_DN = Sqrt_enable_SO?Sqrt_R2:Iteration_cell_sum_AMASK_D[1];
            else
               Partial_remainder_DN = Partial_remainder_DP;
          end
        2'b10:
          begin
            if(Fsm_enable_S)
               Partial_remainder_DN = Sqrt_enable_SO?Sqrt_R3:Iteration_cell_sum_AMASK_D[2];
            else
               Partial_remainder_DN = Partial_remainder_DP;
          end
        2'b11:
          begin
            if(Fsm_enable_S)
               Partial_remainder_DN = Sqrt_enable_SO?Sqrt_R4:Iteration_cell_sum_AMASK_D[3];
            else
               Partial_remainder_DN = Partial_remainder_DP;
          end
        endcase
     end
   always_ff @(posedge Clk_CI, negedge Rst_RBI)   
     begin
        if(~Rst_RBI)
          begin
             Partial_remainder_DP <= '0;
          end
        else
          begin
             Partial_remainder_DP <= Partial_remainder_DN;
          end
    end
   logic [C_MANT_FP64+4:0] Quotient_DN;
  always_comb                                                      
    begin
      case (Iteration_unit_num_S)
        2'b00:
          begin
            if(Fsm_enable_S)
               Quotient_DN= Sqrt_enable_SO ? {Quotient_DP[C_MANT_FP64+3:0],Sqrt_quotinent_S[3]} :{Quotient_DP[C_MANT_FP64+3:0],Iteration_cell_carry_D[0]};
            else
               Quotient_DN= Quotient_DP;
          end
        2'b01:
          begin
            if(Fsm_enable_S)
               Quotient_DN= Sqrt_enable_SO ? {Quotient_DP[C_MANT_FP64+2:0],Sqrt_quotinent_S[3:2]} :{Quotient_DP[C_MANT_FP64+2:0],Iteration_cell_carry_D[0],Iteration_cell_carry_D[1]};
            else
               Quotient_DN= Quotient_DP;
          end
        2'b10:
          begin
            if(Fsm_enable_S)
               Quotient_DN= Sqrt_enable_SO ? {Quotient_DP[C_MANT_FP64+1:0],Sqrt_quotinent_S[3:1]} : {Quotient_DP[C_MANT_FP64+1:0],Iteration_cell_carry_D[0],Iteration_cell_carry_D[1],Iteration_cell_carry_D[2]};
            else
               Quotient_DN= Quotient_DP;
          end
        2'b11:
          begin
            if(Fsm_enable_S)
               Quotient_DN= Sqrt_enable_SO ? {Quotient_DP[C_MANT_FP64:0],Sqrt_quotinent_S } : {Quotient_DP[C_MANT_FP64:0],Iteration_cell_carry_D[0],Iteration_cell_carry_D[1],Iteration_cell_carry_D[2],Iteration_cell_carry_D[3]};
            else
               Quotient_DN= Quotient_DP;
          end
        endcase
     end
   always_ff @(posedge Clk_CI, negedge Rst_RBI)   
     begin
        if(~Rst_RBI)
          begin
          Quotient_DP <= '0;
          end
        else
          Quotient_DP <= Quotient_DN;
    end
   
   
   
   generate
     if(Iteration_unit_num_S==2'b00)
       begin
        always_comb
          begin
            case (Format_sel_S)
              2'b00:
                begin
                  case (Precision_ctl_S)
                    6'h00:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32+4:0],{(C_MANT_FP64-C_MANT_FP32){1'b0}}}; 
                      end
                    6'h17:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32:0],{(C_MANT_FP64-C_MANT_FP32+4){1'b0}}}; 
                      end
                    6'h16:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-1:0],{(C_MANT_FP64-C_MANT_FP32+4+1){1'b0}}}; 
                      end
                    6'h15:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-2:0],{(C_MANT_FP64-C_MANT_FP32+4+2){1'b0}}}; 
                      end
                    6'h14:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-3:0],{(C_MANT_FP64-C_MANT_FP32+4+3){1'b0}}}; 
                      end
                    6'h13:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-4:0],{(C_MANT_FP64-C_MANT_FP32+4+4){1'b0}}}; 
                      end
                    6'h12:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-5:0],{(C_MANT_FP64-C_MANT_FP32+4+5){1'b0}}}; 
                      end
                    6'h11:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-6:0],{(C_MANT_FP64-C_MANT_FP32+4+6){1'b0}}}; 
                      end
                    6'h10:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-7:0],{(C_MANT_FP64-C_MANT_FP32+4+7){1'b0}}}; 
                      end
                    6'h0f:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-8:0],{(C_MANT_FP64-C_MANT_FP32+4+8){1'b0}}}; 
                      end
                    6'h0e:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-9:0],{(C_MANT_FP64-C_MANT_FP32+4+9){1'b0}}}; 
                      end
                    6'h0d:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-10:0],{(C_MANT_FP64-C_MANT_FP32+4+10){1'b0}}}; 
                      end
                    6'h0c:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-11:0],{(C_MANT_FP64-C_MANT_FP32+4+11){1'b0}}}; 
                      end
                    6'h0b:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-12:0],{(C_MANT_FP64-C_MANT_FP32+4+12){1'b0}}}; 
                      end
                    6'h0a:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-13:0],{(C_MANT_FP64-C_MANT_FP32+4+13){1'b0}}}; 
                      end
                    6'h09:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-14:0],{(C_MANT_FP64-C_MANT_FP32+4+14){1'b0}}}; 
                      end
                    6'h08:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-15:0],{(C_MANT_FP64-C_MANT_FP32+4+15){1'b0}}}; 
                      end
                    6'h07:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-16:0],{(C_MANT_FP64-C_MANT_FP32+4+16){1'b0}}}; 
                      end
                    default :
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32+4:0],{(C_MANT_FP64-C_MANT_FP32){1'b0}}}; 
                      end
                  endcase
                end
              2'b01:
                begin
                  case (Precision_ctl_S)
                    6'h00:
                      begin
                        Mant_result_prenorm_DO = Quotient_DP[C_MANT_FP64+4:0]; 
                      end
                    6'h34:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64:0],{(4){1'b0}}}; 
                      end
                    6'h33:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-1:0],{(4+1){1'b0}}}; 
                      end
                    6'h32:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-2:0],{(4+2){1'b0}}}; 
                      end
                    6'h31:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-3:0],{(4+3){1'b0}}}; 
                      end
                    6'h30:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-4:0],{(4+4){1'b0}}}; 
                      end
                    6'h2f:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-5:0],{(4+5){1'b0}}}; 
                      end
                    6'h2e:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-6:0],{(4+6){1'b0}}}; 
                      end
                    6'h2d:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-7:0],{(4+7){1'b0}}}; 
                      end
                    6'h2c:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-8:0],{(4+8){1'b0}}}; 
                      end
                    6'h2b:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-9:0],{(4+9){1'b0}}}; 
                      end
                    6'h2a:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-10:0],{(4+10){1'b0}}}; 
                      end
                    6'h29:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-11:0],{(4+11){1'b0}}}; 
                      end
                    6'h28:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-12:0],{(4+12){1'b0}}}; 
                      end
                    6'h27:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-13:0],{(4+13){1'b0}}}; 
                      end
                    6'h26:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-14:0],{(4+14){1'b0}}}; 
                      end
                    6'h25:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-15:0],{(4+15){1'b0}}}; 
                      end
                    6'h24:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-16:0],{(4+16){1'b0}}}; 
                      end
                    6'h23:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-17:0],{(4+17){1'b0}}}; 
                      end
                    6'h22:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-18:0],{(4+18){1'b0}}}; 
                      end
                    6'h21:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-19:0],{(4+19){1'b0}}}; 
                      end
                    6'h20:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-20:0],{(4+20){1'b0}}}; 
                      end
                    6'h1f:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-21:0],{(4+21){1'b0}}}; 
                      end
                    6'h1e:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-22:0],{(4+22){1'b0}}}; 
                      end
                    6'h1d:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-23:0],{(4+23){1'b0}}}; 
                      end
                    6'h1c:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-24:0],{(4+24){1'b0}}}; 
                      end
                    6'h1b:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-25:0],{(4+25){1'b0}}}; 
                      end
                    6'h1a:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-26:0],{(4+26){1'b0}}}; 
                      end
                    6'h19:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-27:0],{(4+27){1'b0}}}; 
                      end
                    6'h18:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-28:0],{(4+28){1'b0}}}; 
                      end
                    6'h17:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-29:0],{(4+29){1'b0}}}; 
                      end
                    6'h16:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-30:0],{(4+30){1'b0}}}; 
                      end
                    6'h15:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-31:0],{(4+31){1'b0}}}; 
                      end
                    6'h14:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-32:0],{(4+32){1'b0}}}; 
                      end
                    6'h13:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-33:0],{(4+33){1'b0}}}; 
                      end
                    6'h12:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-34:0],{(4+34){1'b0}}}; 
                      end
                    6'h11:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-35:0],{(4+35){1'b0}}}; 
                      end
                    6'h10:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-36:0],{(4+36){1'b0}}}; 
                      end
                    6'h0f:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-37:0],{(4+37){1'b0}}}; 
                      end
                    6'h0e:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-38:0],{(4+38){1'b0}}}; 
                      end
                    6'h0d:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-39:0],{(4+39){1'b0}}}; 
                      end
                    6'h0c:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-40:0],{(4+40){1'b0}}}; 
                      end
                    6'h0b:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-41:0],{(4+41){1'b0}}}; 
                      end
                    6'h0a:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-42:0],{(4+42){1'b0}}}; 
                      end
                    6'h09:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-43:0],{(4+43){1'b0}}}; 
                      end
                    6'h08:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-44:0],{(4+44){1'b0}}}; 
                      end
                    6'h07:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-45:0],{(4+45){1'b0}}}; 
                      end
                    default:
                      begin
                        Mant_result_prenorm_DO = Quotient_DP[C_MANT_FP64+4:0]; 
                      end
                  endcase
                end
              2'b10:
                begin
                  case (Precision_ctl_S)
                    6'b00:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16+4:0],{(C_MANT_FP64-C_MANT_FP16){1'b0}}}; 
                      end
                    6'h0a:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16:0],{(C_MANT_FP64-C_MANT_FP16+4){1'b0}}}; 
                      end
                    6'h09:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16-1:0],{(C_MANT_FP64-C_MANT_FP16+4+1){1'b0}}}; 
                      end
                    6'h08:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16-2:0],{(C_MANT_FP64-C_MANT_FP16+4+2){1'b0}}}; 
                      end
                    6'h07:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16-3:0],{(C_MANT_FP64-C_MANT_FP16+4+3){1'b0}}}; 
                      end
                    default :
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16+4:0],{(C_MANT_FP64-C_MANT_FP16){1'b0}}}; 
                      end
                  endcase
                end
              2'b11:
                begin
                  case (Precision_ctl_S)
                    6'b00:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16ALT+4:0],{(C_MANT_FP64-C_MANT_FP16ALT){1'b0}}}; 
                      end
                    6'h07:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16ALT:0],{(C_MANT_FP64-C_MANT_FP16ALT+4){1'b0}}}; 
                      end
                    default :
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16ALT+4:0],{(C_MANT_FP64-C_MANT_FP16ALT){1'b0}}}; 
                      end
                  endcase
                end
            endcase
          end
        end
      endgenerate
   generate
     if(Iteration_unit_num_S==2'b01)
       begin
        always_comb
          begin
            case (Format_sel_S)
              2'b00:
                begin
                  case (Precision_ctl_S)
                    6'h00:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32+4:0],{(C_MANT_FP64-C_MANT_FP32){1'b0}}}; 
                      end
                    6'h17,6'h16:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32:0],{(C_MANT_FP64-C_MANT_FP32+4){1'b0}}}; 
                      end
                    6'h15,6'h14:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-2:0],{(C_MANT_FP64-C_MANT_FP32+4+2){1'b0}}}; 
                      end
                    6'h13,6'h12:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-4:0],{(C_MANT_FP64-C_MANT_FP32+4+4){1'b0}}}; 
                      end
                    6'h11,6'h10:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-6:0],{(C_MANT_FP64-C_MANT_FP32+4+6){1'b0}}}; 
                      end
                    6'h0f,6'h0e:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-8:0],{(C_MANT_FP64-C_MANT_FP32+4+8){1'b0}}}; 
                      end
                    6'h0d,6'h0c:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-10:0],{(C_MANT_FP64-C_MANT_FP32+4+10){1'b0}}}; 
                      end
                    6'h0b,6'h0a:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-12:0],{(C_MANT_FP64-C_MANT_FP32+4+12){1'b0}}}; 
                      end
                    6'h09,6'h08:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-14:0],{(C_MANT_FP64-C_MANT_FP32+4+14){1'b0}}}; 
                      end
                    6'h07,6'h06:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-16:0],{(C_MANT_FP64-C_MANT_FP32+4+16){1'b0}}}; 
                      end
                    default:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32+4:0],{(C_MANT_FP64-C_MANT_FP32){1'b0}}}; 
                      end
                  endcase
                end
              2'b01:
                begin
                  case (Precision_ctl_S)
                    6'h00:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64+3:0],1'b0}; 
                      end
                    6'h34:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64+1:1],{(4){1'b0}} }; 
                      end
                    6'h33,6'h32:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-1:0],{(4+1){1'b0}} }; 
                      end
                    6'h31,6'h30:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-3:0],{(4+3){1'b0}} }; 
                      end
                    6'h2f,6'h2e:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-5:0],{(4+5){1'b0}} }; 
                      end
                    6'h2d,6'h2c:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-7:0],{(4+7){1'b0}} }; 
                      end
                    6'h2b,6'h2a:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-9:0],{(4+9){1'b0}} }; 
                      end
                    6'h29,6'h28:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-11:0],{(4+11){1'b0}} }; 
                      end
                    6'h27,6'h26:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-13:0],{(4+13){1'b0}} }; 
                      end
                    6'h25,6'h24:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-15:0],{(4+15){1'b0}} }; 
                      end
                    6'h23,6'h22:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-17:0],{(4+17){1'b0}} }; 
                      end
                    6'h21,6'h20:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-19:0],{(4+19){1'b0}} }; 
                      end
                    6'h1f,6'h1e:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-21:0],{(4+21){1'b0}} }; 
                      end
                    6'h1d,6'h1c:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-23:0],{(4+23){1'b0}} }; 
                      end
                    6'h1b,6'h1a:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-25:0],{(4+25){1'b0}} }; 
                      end
                    6'h19,6'h18:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-27:0],{(4+27){1'b0}} }; 
                      end
                    6'h17,6'h16:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-29:0],{(4+29){1'b0}} }; 
                      end
                    6'h15,6'h14:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-31:0],{(4+31){1'b0}} }; 
                      end
                    6'h13,6'h12:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-33:0],{(4+33){1'b0}} }; 
                      end
                    6'h11,6'h10:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-35:0],{(4+35){1'b0}} }; 
                      end
                    6'h0f,6'h0e:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-37:0],{(4+37){1'b0}} }; 
                      end
                    6'h0d,6'h0c:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-39:0],{(4+39){1'b0}} }; 
                      end
                    6'h0b,6'h0a:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-41:0],{(4+41){1'b0}} }; 
                      end
                    6'h09,6'h08:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-43:0],{(4+43){1'b0}} }; 
                      end
                    6'h07:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-45:0],{(4+45){1'b0}} }; 
                      end
                    default:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64+3:0],1'b0}; 
                      end
                  endcase
                end
              2'b10:
                begin
                  case (Precision_ctl_S)
                    6'b00:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16+3:0],{(C_MANT_FP64-C_MANT_FP16+1){1'b0}} }; 
                      end
                    6'h0a:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16+1:1],{(C_MANT_FP64-C_MANT_FP16+4){1'b0}} }; 
                      end
                    6'h09,6'h08:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16-1:0],{(C_MANT_FP64-C_MANT_FP16+4+1){1'b0}} }; 
                      end
                    6'h07:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16-3:0],{(C_MANT_FP64-C_MANT_FP16+4+3){1'b0}} }; 
                      end
                    default :
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16+4:0],{(C_MANT_FP64-C_MANT_FP16){1'b0}} }; 
                      end
                  endcase
                end
              2'b11:
                begin
                  case (Precision_ctl_S)
                    6'b00:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16ALT+4:0],{(C_MANT_FP64-C_MANT_FP16ALT){1'b0}} }; 
                      end
                    6'h07:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16ALT:0],{(C_MANT_FP64-C_MANT_FP16ALT+4){1'b0}} }; 
                      end
                    default :
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16ALT+4:0],{(C_MANT_FP64-C_MANT_FP16ALT){1'b0}} }; 
                      end
                  endcase
                end
            endcase
          end
       end
     endgenerate
   generate
     if(Iteration_unit_num_S==2'b10)
       begin
        always_comb
          begin
            case (Format_sel_S)
              2'b00:
                begin
                  case (Precision_ctl_S)
                    6'h00:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32+3:0],{(C_MANT_FP64-C_MANT_FP32+1){1'b0}}}; 
                      end
                    6'h17,6'h16,6'h15:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32:0],{(C_MANT_FP64-C_MANT_FP32+4){1'b0}}}; 
                      end
                    6'h14,6'h13,6'h12:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-3:0],{(C_MANT_FP64-C_MANT_FP32+4+3){1'b0}}}; 
                      end
                    6'h11,6'h10,6'h0f:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-6:0],{(C_MANT_FP64-C_MANT_FP32+4+6){1'b0}}}; 
                      end
                    6'h0e,6'h0d,6'h0c:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-9:0],{(C_MANT_FP64-C_MANT_FP32+4+9){1'b0}}}; 
                      end
                    6'h0b,6'h0a,6'h09:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-12:0],{(C_MANT_FP64-C_MANT_FP32+4+12){1'b0}}}; 
                      end
                    6'h08,6'h07,6'h06:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-15:0],{(C_MANT_FP64-C_MANT_FP32+4+15){1'b0}}}; 
                      end
                    default:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32+3:0],{(C_MANT_FP64-C_MANT_FP32+1){1'b0}}}; 
                      end
                  endcase
                end
              2'b01:
                begin
                  case (Precision_ctl_S)
                    6'h00:
                      begin
                        Mant_result_prenorm_DO = Quotient_DP[C_MANT_FP64+4:0]; 
                      end
                    6'h34,6'h33:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64+1:1],{(4){1'b0}} }; 
                      end
                    6'h32,6'h31,6'h30:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-2:0],{(4+2){1'b0}} }; 
                      end
                    6'h2f,6'h2e,6'h2d:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-5:0],{(4+5){1'b0}} }; 
                      end
                    6'h2c,6'h2b,6'h2a:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-8:0],{(4+8){1'b0}} }; 
                      end
                    6'h29,6'h28,6'h27:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-11:0],{(4+11){1'b0}} }; 
                      end
                    6'h26,6'h25,6'h24:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-14:0],{(4+14){1'b0}} }; 
                      end
                    6'h23,6'h22,6'h21:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-17:0],{(4+17){1'b0}} }; 
                      end
                    6'h20,6'h1f,6'h1e:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-20:0],{(4+20){1'b0}} }; 
                      end
                    6'h1d,6'h1c,6'h1b:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-23:0],{(4+23){1'b0}} }; 
                      end
                    6'h1a,6'h19,6'h18:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-26:0],{(4+26){1'b0}} }; 
                      end
                    6'h17,6'h16,6'h15:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-29:0],{(4+29){1'b0}} }; 
                      end
                    6'h14,6'h13,6'h12:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-32:0],{(4+32){1'b0}} }; 
                      end
                    6'h11,6'h10,6'h0f:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-35:0],{(4+35){1'b0}} }; 
                      end
                    6'h0e,6'h0d,6'h0c:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-38:0],{(4+38){1'b0}} }; 
                      end
                    6'h0b,6'h0a,6'h09:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-41:0],{(4+41){1'b0}} }; 
                      end
                    6'h08,6'h07,6'h06:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-44:0],{(4+44){1'b0}} }; 
                      end
                    default:
                      begin
                        Mant_result_prenorm_DO = Quotient_DP[C_MANT_FP64+4:0]; 
                      end
                  endcase
                end
              2'b10:
                begin
                  case (Precision_ctl_S)
                    6'b00:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16+4:0],{(C_MANT_FP64-C_MANT_FP16){1'b0}} }; 
                      end
                    6'h0a,6'h09:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16+1:1],{(C_MANT_FP64-C_MANT_FP16+4){1'b0}} }; 
                      end
                    6'h08,6'h07,6'h06:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16-2:0],{(C_MANT_FP64-C_MANT_FP16+4+2){1'b0}} }; 
                      end
                    default :
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16+4:0],{(C_MANT_FP64-C_MANT_FP16){1'b0}} }; 
                      end
                  endcase
                end
              2'b11:
                begin
                  case (Precision_ctl_S)
                    6'b00:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16ALT+4:0],{(C_MANT_FP64-C_MANT_FP16ALT){1'b0}} }; 
                      end
                    6'h07,6'h06:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16ALT+1:1],{(C_MANT_FP64-C_MANT_FP16ALT+4){1'b0}} }; 
                      end
                    default :
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16ALT+4:0],{(C_MANT_FP64-C_MANT_FP16ALT){1'b0}} }; 
                      end
                  endcase
                end
            endcase
          end
        end
      endgenerate
   generate
     if(Iteration_unit_num_S==2'b11)
       begin
        always_comb
          begin
            case (Format_sel_S)
              2'b00:
                begin
                  case (Precision_ctl_S)
                    6'h00:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32+4:0],{(C_MANT_FP64-C_MANT_FP32){1'b0}}}; 
                      end
                    6'h17,6'h16,6'h15,6'h14:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32:0],{(C_MANT_FP64-C_MANT_FP32+4){1'b0}}}; 
                      end
                    6'h13,6'h12,6'h11,6'h10:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-4:0],{(C_MANT_FP64-C_MANT_FP32+4+4){1'b0}}}; 
                      end
                    6'h0f,6'h0e,6'h0d,6'h0c:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-8:0],{(C_MANT_FP64-C_MANT_FP32+4+8){1'b0}}}; 
                      end
                    6'h0b,6'h0a,6'h09,6'h08:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-12:0],{(C_MANT_FP64-C_MANT_FP32+4+12){1'b0}}}; 
                      end
                    6'h07,6'h06:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32-16:0],{(C_MANT_FP64-C_MANT_FP32+4+16){1'b0}}}; 
                      end
                    default:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP32+4:0],{(C_MANT_FP64-C_MANT_FP32){1'b0}}}; 
                      end
                  endcase
                end
              2'b01:
                begin
                  case (Precision_ctl_S)
                    6'h00:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64+3:0],{(1){1'b0}}}; 
                      end
                    6'h34:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64+3:0],{(1){1'b0}} }; 
                      end
                    6'h33,6'h32,6'h31,6'h30:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-1:0],{(5){1'b0}} }; 
                      end
                    6'h2f,6'h2e,6'h2d,6'h2c:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-5:0],{(9){1'b0}} }; 
                      end
                    6'h2b,6'h2a,6'h29,6'h28:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-9:0],{(13){1'b0}} }; 
                      end
                    6'h27,6'h26,6'h25,6'h24:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-13:0],{(17){1'b0}} }; 
                      end
                    6'h23,6'h22,6'h21,6'h20:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-17:0],{(21){1'b0}} }; 
                      end
                    6'h1f,6'h1e,6'h1d,6'h1c:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-21:0],{(25){1'b0}} }; 
                      end
                    6'h1b,6'h1a,6'h19,6'h18:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-25:0],{(29){1'b0}} }; 
                      end
                    6'h17,6'h16,6'h15,6'h14:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-29:0],{(33){1'b0}} }; 
                      end
                    6'h13,6'h12,6'h11,6'h10:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-33:0],{(37){1'b0}} }; 
                      end
                    6'h0f,6'h0e,6'h0d,6'h0c:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-37:0],{(41){1'b0}} }; 
                      end
                    6'h0b,6'h0a,6'h09,6'h08:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-41:0],{(45){1'b0}} }; 
                      end
                    6'h07,6'h06:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64-45:0],{(49){1'b0}} }; 
                      end
                    default:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP64+3:0],{(1){1'b0}}}; 
                      end
                  endcase
                end
              2'b10:
                begin
                  case (Precision_ctl_S)
                    6'b00:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16+5:0],{(C_MANT_FP64-C_MANT_FP16-1){1'b0}} }; 
                      end
                    6'h0a,6'h09,6'h08:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16+1:1],{(C_MANT_FP64-C_MANT_FP16+4){1'b0}} }; 
                      end
                    6'h07,6'h06:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16+1-4:0],{(C_MANT_FP64-C_MANT_FP16+4+3){1'b0}} }; 
                      end
                    default :
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16+5:0],{(C_MANT_FP64-C_MANT_FP16-1){1'b0}} }; 
                      end
                  endcase
                end
              2'b11:
                begin
                  case (Precision_ctl_S)
                    6'b00:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16ALT+4:0],{(C_MANT_FP64-C_MANT_FP16ALT){1'b0}} }; 
                      end
                    6'h07,6'h06:
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16ALT:0],{(C_MANT_FP64-C_MANT_FP16ALT+4){1'b0}} }; 
                      end
                    default :
                      begin
                        Mant_result_prenorm_DO = {Quotient_DP[C_MANT_FP16ALT+4:0],{(C_MANT_FP64-C_MANT_FP16ALT){1'b0}} }; 
                      end
                  endcase
                end
            endcase
          end
        end
      endgenerate
   logic   [C_EXP_FP64+1:0]    Exp_result_prenorm_DN,Exp_result_prenorm_DP;
   logic   [C_EXP_FP64+1:0]                                Exp_add_a_D;
   logic   [C_EXP_FP64+1:0]                                Exp_add_b_D;
   logic   [C_EXP_FP64+1:0]                                Exp_add_c_D;
  integer                                                 C_BIAS_AONE, C_HALF_BIAS;
  always_comb
    begin  
      case (Format_sel_S)
        2'b00:
          begin
            C_BIAS_AONE =C_BIAS_AONE_FP32;
            C_HALF_BIAS =C_HALF_BIAS_FP32;
          end
        2'b01:
          begin
            C_BIAS_AONE =C_BIAS_AONE_FP64;
            C_HALF_BIAS =C_HALF_BIAS_FP64;
          end
        2'b10:
          begin
            C_BIAS_AONE =C_BIAS_AONE_FP16;
            C_HALF_BIAS =C_HALF_BIAS_FP16;
          end
        2'b11:
          begin
            C_BIAS_AONE =C_BIAS_AONE_FP16ALT;
            C_HALF_BIAS =C_HALF_BIAS_FP16ALT;
          end
        endcase
    end
  assign Exp_add_a_D = {Sqrt_start_dly_S?{Exp_num_DI[C_EXP_FP64],Exp_num_DI[C_EXP_FP64],Exp_num_DI[C_EXP_FP64],Exp_num_DI[C_EXP_FP64:1]}:{Exp_num_DI[C_EXP_FP64],Exp_num_DI[C_EXP_FP64],Exp_num_DI}};
  assign Exp_add_b_D = {Sqrt_start_dly_S?{1'b0,{C_EXP_ZERO_FP64},Exp_num_DI[0]}:{~Exp_den_DI[C_EXP_FP64],~Exp_den_DI[C_EXP_FP64],~Exp_den_DI}};
  assign Exp_add_c_D = {Div_start_dly_S?{{C_BIAS_AONE}}:{{C_HALF_BIAS}}};
  assign Exp_result_prenorm_DN  = (Start_dly_S)?{Exp_add_a_D + Exp_add_b_D + Exp_add_c_D}:Exp_result_prenorm_DP;
  always_ff @(posedge Clk_CI, negedge Rst_RBI)
   begin
      if(~Rst_RBI)
        begin
          Exp_result_prenorm_DP <= '0;
        end
      else
        begin
          Exp_result_prenorm_DP<=  Exp_result_prenorm_DN;
        end
   end
  assign Exp_result_prenorm_DO = Exp_result_prenorm_DP;
endmodule
import defs_div_sqrt_mvp::*;
module div_sqrt_mvp_wrapper
#(
   parameter   PrePipeline_depth_S             =        0,  
   parameter   PostPipeline_depth_S            =        2  
)
  (
   input logic                            Clk_CI,
   input logic                            Rst_RBI,
   input logic                            Div_start_SI,
   input logic                            Sqrt_start_SI,
   
   input logic [C_OP_FP64-1:0]            Operand_a_DI,
   input logic [C_OP_FP64-1:0]            Operand_b_DI,
   
   input logic [C_RM-1:0]                 RM_SI,    
   input logic [C_PC-1:0]                 Precision_ctl_SI, 
   input logic [C_FS-1:0]                 Format_sel_SI,  
   input logic                            Kill_SI,
   
   output logic [C_OP_FP64-1:0]           Result_DO,
   
   output logic [4:0]                     Fflags_SO,
   output logic                           Ready_SO,
   output logic                           Done_SO
 );
   logic                                 Div_start_S_S,Sqrt_start_S_S;
   logic [C_OP_FP64-1:0]                 Operand_a_S_D;
   logic [C_OP_FP64-1:0]                 Operand_b_S_D;
   
   logic [C_RM-1:0]                      RM_S_S;    
   logic [C_PC-1:0]                      Precision_ctl_S_S; 
   logic [C_FS-1:0]                      Format_sel_S_S;  
   logic                                 Kill_S_S;
  logic [C_OP_FP64-1:0]                  Result_D;
  logic                                  Ready_S;
  logic                                  Done_S;
  logic [4:0]                            Fflags_S;
  generate
    if(PrePipeline_depth_S==1)
      begin
         div_sqrt_top_mvp  div_top_U0  
          (
           .Clk_CI                 (Clk_CI),
           .Rst_RBI                (Rst_RBI),
           .Div_start_SI           (Div_start_S_S),
           .Sqrt_start_SI          (Sqrt_start_S_S),
           
           .Operand_a_DI          (Operand_a_S_D),
           .Operand_b_DI          (Operand_b_S_D),
           .RM_SI                 (RM_S_S),    
           .Precision_ctl_SI      (Precision_ctl_S_S),
           .Format_sel_SI         (Format_sel_S_S),
           .Kill_SI               (Kill_S_S),
           .Result_DO             (Result_D),
           .Fflags_SO             (Fflags_S),
           .Ready_SO              (Ready_S),
           .Done_SO               (Done_S)
         );
           always_ff @(posedge Clk_CI, negedge Rst_RBI)
             begin
                if(~Rst_RBI)
                  begin
                    Div_start_S_S<='0;
                    Sqrt_start_S_S<=1'b0;
                    Operand_a_S_D<='0;
                    Operand_b_S_D<='0;
                    RM_S_S <=1'b0;
                    Precision_ctl_S_S<='0;
                    Format_sel_S_S<='0;
                    Kill_S_S<='0;
                  end
                else
                  begin
                    Div_start_S_S<=Div_start_SI;
                    Sqrt_start_S_S<=Sqrt_start_SI;
                    Operand_a_S_D<=Operand_a_DI;
                    Operand_b_S_D<=Operand_b_DI;
                    RM_S_S <=RM_SI;
                    Precision_ctl_S_S<=Precision_ctl_SI;
                    Format_sel_S_S<=Format_sel_SI;
                    Kill_S_S<=Kill_SI;
                  end
            end
     end
     else
      begin
          div_sqrt_top_mvp  div_top_U0  
          (
           .Clk_CI                 (Clk_CI),
           .Rst_RBI                (Rst_RBI),
           .Div_start_SI           (Div_start_SI),
           .Sqrt_start_SI          (Sqrt_start_SI),
           
           .Operand_a_DI          (Operand_a_DI),
           .Operand_b_DI          (Operand_b_DI),
           .RM_SI                 (RM_SI),    
           .Precision_ctl_SI      (Precision_ctl_SI),
           .Format_sel_SI         (Format_sel_SI),
           .Kill_SI               (Kill_SI),
           .Result_DO             (Result_D),
           .Fflags_SO             (Fflags_S),
           .Ready_SO              (Ready_S),
           .Done_SO               (Done_S)
         );
      end
  endgenerate
   
   
   
  logic [C_OP_FP64-1:0]         Result_dly_S_D;
  logic                         Ready_dly_S_S;
  logic                         Done_dly_S_S;
  logic [4:0]                   Fflags_dly_S_S;
   always_ff @(posedge Clk_CI, negedge Rst_RBI)
     begin
        if(~Rst_RBI)
          begin
            Result_dly_S_D<='0;
            Ready_dly_S_S<=1'b0;
            Done_dly_S_S<=1'b0;
            Fflags_dly_S_S<=1'b0;
          end
        else
          begin
            Result_dly_S_D<=Result_D;
            Ready_dly_S_S<=Ready_S;
            Done_dly_S_S<=Done_S;
            Fflags_dly_S_S<=Fflags_S;
          end
    end
   
   
   
  logic [C_OP_FP64-1:0]         Result_dly_D_D;
  logic                         Ready_dly_D_S;
  logic                         Done_dly_D_S;
  logic [4:0]                   Fflags_dly_D_S;
  generate
    if(PostPipeline_depth_S==2)
      begin
        always_ff @(posedge Clk_CI, negedge Rst_RBI)
          begin
            if(~Rst_RBI)
              begin
                Result_dly_D_D<='0;
                Ready_dly_D_S<=1'b0;
                Done_dly_D_S<=1'b0;
                Fflags_dly_D_S<=1'b0;
              end
           else
             begin
               Result_dly_D_D<=Result_dly_S_D;
               Ready_dly_D_S<=Ready_dly_S_S;
               Done_dly_D_S<=Done_dly_S_S;
               Fflags_dly_D_S<=Fflags_dly_S_S;
             end
          end
        assign  Result_DO = Result_dly_D_D;
        assign  Ready_SO  = Ready_dly_D_S;
        assign  Done_SO  = Done_dly_D_S;
        assign  Fflags_SO=Fflags_dly_D_S;
       end
     else
       begin
         assign  Result_DO = Result_dly_S_D;
         assign  Ready_SO  = Ready_dly_S_S;
         assign  Done_SO   = Done_dly_S_S;
         assign  Fflags_SO  = Fflags_dly_S_S;
       end
   endgenerate
endmodule 
import defs_div_sqrt_mvp::*;
module div_sqrt_top_mvp
  (
   input logic                            Clk_CI,
   input logic                            Rst_RBI,
   input logic                            Div_start_SI,
   input logic                            Sqrt_start_SI,
   
   input logic [C_OP_FP64-1:0]            Operand_a_DI,
   input logic [C_OP_FP64-1:0]            Operand_b_DI,
   
   input logic [C_RM-1:0]                 RM_SI,    
   input logic [C_PC-1:0]                 Precision_ctl_SI, 
   input logic [C_FS-1:0]                 Format_sel_SI,  
   input logic                            Kill_SI,
   
   output logic [C_OP_FP64-1:0]           Result_DO,
   
   output logic [4:0]                     Fflags_SO,
   output logic                           Ready_SO,
   output logic                           Done_SO
 );
   
   logic [C_EXP_FP64:0]                 Exp_a_D;
   logic [C_EXP_FP64:0]                 Exp_b_D;
   logic [C_MANT_FP64:0]                Mant_a_D;
   logic [C_MANT_FP64:0]                Mant_b_D;
   logic [C_EXP_FP64+1:0]               Exp_z_D;
   logic [C_MANT_FP64+4:0]              Mant_z_D;
   logic                                Sign_z_D;
   logic                                Start_S;
   logic [C_RM-1:0]                     RM_dly_S;
   logic                                Div_enable_S;
   logic                                Sqrt_enable_S;
   logic                                Inf_a_S;
   logic                                Inf_b_S;
   logic                                Zero_a_S;
   logic                                Zero_b_S;
   logic                                NaN_a_S;
   logic                                NaN_b_S;
   logic                                SNaN_S;
   logic                                Special_case_SB,Special_case_dly_SB;
   logic Full_precision_S;
   logic FP32_S;
   logic FP64_S;
   logic FP16_S;
   logic FP16ALT_S;
 preprocess_mvp  preprocess_U0
 (
   .Clk_CI                (Clk_CI             ),
   .Rst_RBI               (Rst_RBI            ),
   .Div_start_SI          (Div_start_SI       ),
   .Sqrt_start_SI         (Sqrt_start_SI      ),
   .Ready_SI              (Ready_SO           ),
   .Operand_a_DI          (Operand_a_DI       ),
   .Operand_b_DI          (Operand_b_DI       ),
   .RM_SI                 (RM_SI              ),
   .Format_sel_SI         (Format_sel_SI      ),
   .Start_SO              (Start_S            ),
   .Exp_a_DO_norm         (Exp_a_D            ),
   .Exp_b_DO_norm         (Exp_b_D            ),
   .Mant_a_DO_norm        (Mant_a_D           ),
   .Mant_b_DO_norm        (Mant_b_D           ),
   .RM_dly_SO             (RM_dly_S           ),
   .Sign_z_DO             (Sign_z_D           ),
   .Inf_a_SO              (Inf_a_S            ),
   .Inf_b_SO              (Inf_b_S            ),
   .Zero_a_SO             (Zero_a_S           ),
   .Zero_b_SO             (Zero_b_S           ),
   .NaN_a_SO              (NaN_a_S            ),
   .NaN_b_SO              (NaN_b_S            ),
   .SNaN_SO               (SNaN_S             ),
   .Special_case_SBO      (Special_case_SB    ),
   .Special_case_dly_SBO  (Special_case_dly_SB)
   );
 nrbd_nrsc_mvp   nrbd_nrsc_U0
  (
   .Clk_CI                (Clk_CI             ),
   .Rst_RBI               (Rst_RBI            ),
   .Div_start_SI          (Div_start_SI       ) ,
   .Sqrt_start_SI         (Sqrt_start_SI      ),
   .Start_SI              (Start_S            ),
   .Kill_SI               (Kill_SI            ),
   .Special_case_SBI      (Special_case_SB    ),
   .Special_case_dly_SBI  (Special_case_dly_SB),
   .Div_enable_SO         (Div_enable_S       ),
   .Sqrt_enable_SO        (Sqrt_enable_S      ),
   .Precision_ctl_SI      (Precision_ctl_SI   ),
   .Format_sel_SI         (Format_sel_SI      ),
   .Exp_a_DI              (Exp_a_D            ),
   .Exp_b_DI              (Exp_b_D            ),
   .Mant_a_DI             (Mant_a_D           ),
   .Mant_b_DI             (Mant_b_D           ),
   .Full_precision_SO     (Full_precision_S   ),
   .FP32_SO               (FP32_S             ),
   .FP64_SO               (FP64_S             ),
   .FP16_SO               (FP16_S             ),
   .FP16ALT_SO            (FP16ALT_S          ),
   .Ready_SO              (Ready_SO           ),
   .Done_SO               (Done_SO            ),
   .Exp_z_DO              (Exp_z_D            ),
   .Mant_z_DO             (Mant_z_D           )
    );
 norm_div_sqrt_mvp  fpu_norm_U0
  (
   .Mant_in_DI            (Mant_z_D           ),
   .Exp_in_DI             (Exp_z_D            ),
   .Sign_in_DI            (Sign_z_D           ),
   .Div_enable_SI         (Div_enable_S       ),
   .Sqrt_enable_SI        (Sqrt_enable_S      ),
   .Inf_a_SI              (Inf_a_S            ),
   .Inf_b_SI              (Inf_b_S            ),
   .Zero_a_SI             (Zero_a_S           ),
   .Zero_b_SI             (Zero_b_S           ),
   .NaN_a_SI              (NaN_a_S            ),
   .NaN_b_SI              (NaN_b_S            ),
   .SNaN_SI               (SNaN_S             ),
   .RM_SI                 (RM_dly_S           ),
   .Full_precision_SI     (Full_precision_S   ),
   .FP32_SI               (FP32_S             ),
   .FP64_SI               (FP64_S             ),
   .FP16_SI               (FP16_S             ),
   .FP16ALT_SI            (FP16ALT_S          ),
   .Result_DO             (Result_DO          ),
   .Fflags_SO             (Fflags_SO          ) 
   );
endmodule
module iteration_div_sqrt_mvp
#(
   parameter   WIDTH=25
)
  (
   input logic [WIDTH-1:0]      A_DI,
   input logic [WIDTH-1:0]      B_DI,
   input logic                  Div_enable_SI,
   input logic                  Div_start_dly_SI,
   input logic                  Sqrt_enable_SI,
   input logic [1:0]            D_DI,
   output logic [1:0]           D_DO,
   output logic [WIDTH-1:0]     Sum_DO,
   output logic                 Carry_out_DO
    );
   logic                        D_carry_D;
   logic                        Sqrt_cin_D;
   logic                        Cin_D;
   assign D_DO[0]=~D_DI[0];
   assign D_DO[1]=~(D_DI[1] ^ D_DI[0]);
   assign D_carry_D=D_DI[1] | D_DI[0];
   assign Sqrt_cin_D=Sqrt_enable_SI&&D_carry_D;
   assign Cin_D=Div_enable_SI?1'b0:Sqrt_cin_D;
   assign {Carry_out_DO,Sum_DO}=A_DI+B_DI+Cin_D;
endmodule
import defs_div_sqrt_mvp::*;
module norm_div_sqrt_mvp
  (
   input logic [C_MANT_FP64+4:0]                Mant_in_DI,  
   input logic signed [C_EXP_FP64+1:0]          Exp_in_DI,
   input logic                                  Sign_in_DI,
   input logic                                  Div_enable_SI,
   input logic                                  Sqrt_enable_SI,
   input logic                                  Inf_a_SI,
   input logic                                  Inf_b_SI,
   input logic                                  Zero_a_SI,
   input logic                                  Zero_b_SI,
   input logic                                  NaN_a_SI,
   input logic                                  NaN_b_SI,
   input logic                                  SNaN_SI,
   input logic [C_RM-1:0]                       RM_SI,
   input logic                                  Full_precision_SI,
   input logic                                  FP32_SI,
   input logic                                  FP64_SI,
   input logic                                  FP16_SI,
   input logic                                  FP16ALT_SI,
   
   output logic [C_EXP_FP64+C_MANT_FP64:0]      Result_DO,
   output logic [4:0]                           Fflags_SO 
   );
   logic                                        Sign_res_D;
   logic                                        NV_OP_S;
   logic                                        Exp_OF_S;
   logic                                        Exp_UF_S;
   logic                                        Div_Zero_S;
   logic                                        In_Exact_S;
   
   
   
   logic [C_MANT_FP64:0]                        Mant_res_norm_D;
   logic [C_EXP_FP64-1:0]                       Exp_res_norm_D;
   
   
   
  logic  [C_EXP_FP64+1:0]                       Exp_Max_RS_FP64_D;
  logic  [C_EXP_FP32+1:0]                       Exp_Max_RS_FP32_D;
  logic  [C_EXP_FP16+1:0]                       Exp_Max_RS_FP16_D;
  logic  [C_EXP_FP16ALT+1:0]                    Exp_Max_RS_FP16ALT_D;
  
  assign Exp_Max_RS_FP64_D=Exp_in_DI[C_EXP_FP64:0]+C_MANT_FP64+1; 
  assign Exp_Max_RS_FP32_D=Exp_in_DI[C_EXP_FP32:0]+C_MANT_FP32+1; 
  assign Exp_Max_RS_FP16_D=Exp_in_DI[C_EXP_FP16:0]+C_MANT_FP16+1; 
  assign Exp_Max_RS_FP16ALT_D=Exp_in_DI[C_EXP_FP16ALT:0]+C_MANT_FP16ALT+1; 
  logic  [C_EXP_FP64+1:0]                       Num_RS_D;
  assign Num_RS_D=~Exp_in_DI+1+1;            
  logic  [C_MANT_FP64:0]                        Mant_RS_D;
  logic  [C_MANT_FP64+4:0]                      Mant_forsticky_D;
  assign  {Mant_RS_D,Mant_forsticky_D} ={Mant_in_DI,{(C_MANT_FP64+1){1'b0}} } >>(Num_RS_D); 
  logic [C_EXP_FP64+1:0]                        Exp_subOne_D;
  assign Exp_subOne_D = Exp_in_DI -1;
   
   logic [1:0]                                  Mant_lower_D;
   logic                                        Mant_sticky_bit_D;
   logic [C_MANT_FP64+4:0]                      Mant_forround_D;
   always_comb
     begin
       if(NaN_a_SI)  
         begin
           Div_Zero_S=1'b0;
           Exp_OF_S=1'b0;
           Exp_UF_S=1'b0;
           Mant_res_norm_D={1'b0,C_MANT_NAN_FP64};
           Exp_res_norm_D='1;
           Mant_forround_D='0;
           Sign_res_D=1'b0;
           NV_OP_S = SNaN_SI;
         end
      else if(NaN_b_SI)   
        begin
          Div_Zero_S=1'b0;
          Exp_OF_S=1'b0;
          Exp_UF_S=1'b0;
          Mant_res_norm_D={1'b0,C_MANT_NAN_FP64};
          Exp_res_norm_D='1;
          Mant_forround_D='0;
          Sign_res_D=1'b0;
          NV_OP_S = SNaN_SI;
        end
      else if(Inf_a_SI)
        begin
          if(Div_enable_SI&&Inf_b_SI)                     
            begin
              Div_Zero_S=1'b0;
              Exp_OF_S=1'b0;
              Exp_UF_S=1'b0;
              Mant_res_norm_D={1'b0,C_MANT_NAN_FP64};
              Exp_res_norm_D='1;
              Mant_forround_D='0;
              Sign_res_D=1'b0;
              NV_OP_S = 1'b1;
            end
          else if (Sqrt_enable_SI && Sign_in_DI) begin 
            Div_Zero_S=1'b0;
            Exp_OF_S=1'b0;
            Exp_UF_S=1'b0;
            Mant_res_norm_D={1'b0,C_MANT_NAN_FP64};
            Exp_res_norm_D='1;
            Mant_forround_D='0;
            Sign_res_D=1'b0;
            NV_OP_S = 1'b1;
          end else begin
            Div_Zero_S=1'b0;
            Exp_OF_S=1'b1;
            Exp_UF_S=1'b0;
            Mant_res_norm_D= '0;
            Exp_res_norm_D='1;
            Mant_forround_D='0;
            Sign_res_D=Sign_in_DI;
            NV_OP_S = 1'b0;
          end
        end
      else if(Div_enable_SI&&Inf_b_SI)
        begin
          Div_Zero_S=1'b0;
          Exp_OF_S=1'b1;
          Exp_UF_S=1'b0;
          Mant_res_norm_D= '0;
          Exp_res_norm_D='0;
          Mant_forround_D='0;
          Sign_res_D=Sign_in_DI;
          NV_OP_S = 1'b0;
        end
     else if(Zero_a_SI)
       begin
         if(Div_enable_SI&&Zero_b_SI)
           begin
              Div_Zero_S=1'b1;
              Exp_OF_S=1'b0;
              Exp_UF_S=1'b0;
              Mant_res_norm_D={1'b0,C_MANT_NAN_FP64};
              Exp_res_norm_D='1;
              Mant_forround_D='0;
              Sign_res_D=1'b0;
              NV_OP_S = 1'b1;
           end
         else
           begin
             Div_Zero_S=1'b0;
             Exp_OF_S=1'b0;
             Exp_UF_S=1'b0;
             Mant_res_norm_D='0;
             Exp_res_norm_D='0;
             Mant_forround_D='0;
             Sign_res_D=Sign_in_DI;
             NV_OP_S = 1'b0;
           end
       end
     else  if(Div_enable_SI&&(Zero_b_SI))  
       begin
         Div_Zero_S=1'b1;
         Exp_OF_S=1'b0;
         Exp_UF_S=1'b0;
         Mant_res_norm_D='0;
         Exp_res_norm_D='1;
         Mant_forround_D='0;
         Sign_res_D=Sign_in_DI;
         NV_OP_S = 1'b0;
       end
      else if(Sign_in_DI&&Sqrt_enable_SI)   
        begin
          Div_Zero_S=1'b0;
          Exp_OF_S=1'b0;
          Exp_UF_S=1'b0;
          Mant_res_norm_D={1'b0,C_MANT_NAN_FP64};
          Exp_res_norm_D='1;
          Mant_forround_D='0;
          Sign_res_D=1'b0;
          NV_OP_S = 1'b1;
        end
     else if((Exp_in_DI[C_EXP_FP64:0]=='0))
       begin
         if(Mant_in_DI!='0)       
           begin
             Div_Zero_S=1'b0;
             Exp_OF_S=1'b0;
             Exp_UF_S=1'b1;
             Mant_res_norm_D={1'b0,Mant_in_DI[C_MANT_FP64+4:5]};
             Exp_res_norm_D='0;
             Mant_forround_D={Mant_in_DI[4:0],{(C_MANT_FP64){1'b0}} };
             Sign_res_D=Sign_in_DI;
             NV_OP_S = 1'b0;
           end
         else                 
           begin
             Div_Zero_S=1'b0;
             Exp_OF_S=1'b0;
             Exp_UF_S=1'b0;
             Mant_res_norm_D='0;
             Exp_res_norm_D='0;
             Mant_forround_D='0;
             Sign_res_D=Sign_in_DI;
             NV_OP_S = 1'b0;
           end
        end
      else if((Exp_in_DI[C_EXP_FP64:0]==C_EXP_ONE_FP64)&&(~Mant_in_DI[C_MANT_FP64+4]))  
        begin
          Div_Zero_S=1'b0;
          Exp_OF_S=1'b0;
          Exp_UF_S=1'b1;
          Mant_res_norm_D=Mant_in_DI[C_MANT_FP64+4:4];
          Exp_res_norm_D='0;
          Mant_forround_D={Mant_in_DI[3:0],{(C_MANT_FP64+1){1'b0}}};
          Sign_res_D=Sign_in_DI;
          NV_OP_S = 1'b0;
        end
      else if(Exp_in_DI[C_EXP_FP64+1])    
        begin
          if(((~Exp_Max_RS_FP32_D[C_EXP_FP32+1])&&FP32_SI) | ((~Exp_Max_RS_FP64_D[C_EXP_FP64+1])&&FP64_SI) | ((~Exp_Max_RS_FP16_D[C_EXP_FP16+1])&&FP16_SI) | ((~Exp_Max_RS_FP16ALT_D[C_EXP_FP16ALT+1])&&FP16ALT_SI) )    
            begin
              Div_Zero_S=1'b0;
              Exp_OF_S=1'b1;
              Exp_UF_S=1'b0;
              Mant_res_norm_D='0;
              Exp_res_norm_D='0;
              Mant_forround_D='0;
              Sign_res_D=Sign_in_DI;
              NV_OP_S = 1'b0;
            end
          else                    
            begin
              Div_Zero_S=1'b0;
              Exp_OF_S=1'b0;
              Exp_UF_S=1'b1;
              Mant_res_norm_D={Mant_RS_D[C_MANT_FP64:0]};
              Exp_res_norm_D='0;
              Mant_forround_D={Mant_forsticky_D[C_MANT_FP64+4:0]};   
              Sign_res_D=Sign_in_DI;
              NV_OP_S = 1'b0;
            end
        end
      else if( (Exp_in_DI[C_EXP_FP32]&&FP32_SI) | (Exp_in_DI[C_EXP_FP64]&&FP64_SI) | (Exp_in_DI[C_EXP_FP16]&&FP16_SI) | (Exp_in_DI[C_EXP_FP16ALT]&&FP16ALT_SI) )            
        begin
          Div_Zero_S=1'b0;
          Exp_OF_S=1'b1;
          Exp_UF_S=1'b0;
          Mant_res_norm_D='0;
          Exp_res_norm_D='1;
          Mant_forround_D='0;
          Sign_res_D=Sign_in_DI;
          NV_OP_S = 1'b0;
        end
      else if( ((Exp_in_DI[C_EXP_FP32-1:0]=='1)&&FP32_SI) | ((Exp_in_DI[C_EXP_FP64-1:0]=='1)&&FP64_SI) |  ((Exp_in_DI[C_EXP_FP16-1:0]=='1)&&FP16_SI) | ((Exp_in_DI[C_EXP_FP16ALT-1:0]=='1)&&FP16ALT_SI) )
        begin
          if(~Mant_in_DI[C_MANT_FP64+4]) 
            begin
              Div_Zero_S=1'b0;
              Exp_OF_S=1'b0;
              Exp_UF_S=1'b0;
              Mant_res_norm_D=Mant_in_DI[C_MANT_FP64+3:3];
              Exp_res_norm_D=Exp_subOne_D;
              Mant_forround_D={Mant_in_DI[2:0],{(C_MANT_FP64+2){1'b0}}};
              Sign_res_D=Sign_in_DI;
              NV_OP_S = 1'b0;
            end
          else if(Mant_in_DI!='0)         
            begin
              Div_Zero_S=1'b0;
              Exp_OF_S=1'b1;
              Exp_UF_S=1'b0;
              Mant_res_norm_D= '0;
              Exp_res_norm_D='1;
              Mant_forround_D='0;
              Sign_res_D=Sign_in_DI;
              NV_OP_S = 1'b0;
            end
          else                         
            begin
              Div_Zero_S=1'b0;
              Exp_OF_S=1'b1;
              Exp_UF_S=1'b0;
              Mant_res_norm_D= '0;
              Exp_res_norm_D='1;
              Mant_forround_D='0;
              Sign_res_D=Sign_in_DI;
              NV_OP_S = 1'b0;
            end
         end
      else if(Mant_in_DI[C_MANT_FP64+4])  
        begin
           Div_Zero_S=1'b0;
           Exp_OF_S=1'b0;
           Exp_UF_S=1'b0;
           Mant_res_norm_D= Mant_in_DI[C_MANT_FP64+4:4];
           Exp_res_norm_D=Exp_in_DI[C_EXP_FP64-1:0];
           Mant_forround_D={Mant_in_DI[3:0],{(C_MANT_FP64+1){1'b0}}};
           Sign_res_D=Sign_in_DI;
           NV_OP_S = 1'b0;
        end
      else                                   
         begin
           Div_Zero_S=1'b0;
           Exp_OF_S=1'b0;
           Exp_UF_S=1'b0;
           Mant_res_norm_D=Mant_in_DI[C_MANT_FP64+3:3];
           Exp_res_norm_D=Exp_subOne_D;
           Mant_forround_D={Mant_in_DI[2:0],{(C_MANT_FP64+2){1'b0}}};
           Sign_res_D=Sign_in_DI;
           NV_OP_S = 1'b0;
         end
     end
   
   
   
   logic [C_MANT_FP64:0]                   Mant_upper_D;
   logic [C_MANT_FP64+1:0]                 Mant_upperRounded_D;
   logic                                   Mant_roundUp_S;
   logic                                   Mant_rounded_S;
  always_comb 
    begin
      if(FP32_SI)
        begin
          Mant_upper_D = {Mant_res_norm_D[C_MANT_FP64:C_MANT_FP64-C_MANT_FP32], {(C_MANT_FP64-C_MANT_FP32){1'b0}} };
          Mant_lower_D = Mant_res_norm_D[C_MANT_FP64-C_MANT_FP32-1:C_MANT_FP64-C_MANT_FP32-2];
          Mant_sticky_bit_D = | Mant_res_norm_D[C_MANT_FP64-C_MANT_FP32-3:0];
        end
      else if(FP64_SI)
        begin
          Mant_upper_D = Mant_res_norm_D[C_MANT_FP64:0];
          Mant_lower_D = Mant_forround_D[C_MANT_FP64+4:C_MANT_FP64+3];
          Mant_sticky_bit_D = | Mant_forround_D[C_MANT_FP64+3:0];
        end
      else if(FP16_SI)
        begin
          Mant_upper_D = {Mant_res_norm_D[C_MANT_FP64:C_MANT_FP64-C_MANT_FP16], {(C_MANT_FP64-C_MANT_FP16){1'b0}} };
          Mant_lower_D = Mant_res_norm_D[C_MANT_FP64-C_MANT_FP16-1:C_MANT_FP64-C_MANT_FP16-2];
          Mant_sticky_bit_D = | Mant_res_norm_D[C_MANT_FP64-C_MANT_FP16-3:30];
        end
      else  
      begin
          Mant_upper_D = {Mant_res_norm_D[C_MANT_FP64:C_MANT_FP64-C_MANT_FP16ALT], {(C_MANT_FP64-C_MANT_FP16ALT){1'b0}} };
          Mant_lower_D = Mant_res_norm_D[C_MANT_FP64-C_MANT_FP16ALT-1:C_MANT_FP64-C_MANT_FP16ALT-2];
          Mant_sticky_bit_D = | Mant_res_norm_D[C_MANT_FP64-C_MANT_FP16ALT-3:30];
      end
    end
   assign Mant_rounded_S = (|(Mant_lower_D))| Mant_sticky_bit_D;
   always_comb 
     begin
        Mant_roundUp_S = 1'b0;
        case (RM_SI)
          C_RM_NEAREST :
            Mant_roundUp_S = Mant_lower_D[1] && ((Mant_lower_D[0] | Mant_sticky_bit_D )| ( (FP32_SI&&Mant_upper_D[C_MANT_FP64-C_MANT_FP32]) | (FP64_SI&&Mant_upper_D[0]) | (FP16_SI&&Mant_upper_D[C_MANT_FP64-C_MANT_FP16]) | (FP16ALT_SI&&Mant_upper_D[C_MANT_FP64-C_MANT_FP16ALT]) ) );
          C_RM_TRUNC   :
            Mant_roundUp_S = 0;
          C_RM_PLUSINF :
            Mant_roundUp_S = Mant_rounded_S & ~Sign_in_DI;
          C_RM_MINUSINF:
            Mant_roundUp_S = Mant_rounded_S & Sign_in_DI;
          default          :
            Mant_roundUp_S = 0;
        endcase 
     end 
  logic                                 Mant_renorm_S;
  logic  [C_MANT_FP64:0]                Mant_roundUp_Vector_S; 
  assign Mant_roundUp_Vector_S={7'h0,(FP16ALT_SI&&Mant_roundUp_S),2'h0,(FP16_SI&&Mant_roundUp_S),12'h0,(FP32_SI&&Mant_roundUp_S),28'h0,(FP64_SI&&Mant_roundUp_S)};
  assign Mant_upperRounded_D = Mant_upper_D + Mant_roundUp_Vector_S;
  assign Mant_renorm_S       = Mant_upperRounded_D[C_MANT_FP64+1];
  
  
  
  logic [C_MANT_FP64-1:0]               Mant_res_round_D;
  logic [C_EXP_FP64-1:0]                Exp_res_round_D;
  assign Mant_res_round_D = (Mant_renorm_S)?Mant_upperRounded_D[C_MANT_FP64:1]:Mant_upperRounded_D[C_MANT_FP64-1:0]; 
  assign Exp_res_round_D  = Exp_res_norm_D+Mant_renorm_S;
  
  
  
  logic [C_MANT_FP64-1:0]               Mant_before_format_ctl_D;
  logic [C_EXP_FP64-1:0]                Exp_before_format_ctl_D;
  assign Mant_before_format_ctl_D = Full_precision_SI ? Mant_res_round_D : Mant_res_norm_D;
  assign Exp_before_format_ctl_D = Full_precision_SI ? Exp_res_round_D : Exp_res_norm_D;
  always_comb    
    begin  
      if(FP32_SI)
          begin
            Result_DO ={32'hffff_ffff,Sign_res_D,Exp_before_format_ctl_D[C_EXP_FP32-1:0],Mant_before_format_ctl_D[C_MANT_FP64-1:C_MANT_FP64-C_MANT_FP32]};
          end
       else if(FP64_SI)
          begin
            Result_DO ={Sign_res_D,Exp_before_format_ctl_D[C_EXP_FP64-1:0],Mant_before_format_ctl_D[C_MANT_FP64-1:0]};
          end
      else if(FP16_SI)
          begin
            Result_DO ={48'hffff_ffff_ffff,Sign_res_D,Exp_before_format_ctl_D[C_EXP_FP16-1:0],Mant_before_format_ctl_D[C_MANT_FP64-1:C_MANT_FP64-C_MANT_FP16]};
          end
      else
          begin
            Result_DO ={48'hffff_ffff_ffff,Sign_res_D,Exp_before_format_ctl_D[C_EXP_FP16ALT-1:0],Mant_before_format_ctl_D[C_MANT_FP64-1:C_MANT_FP64-C_MANT_FP16ALT]};
          end
    end
assign In_Exact_S = (~Full_precision_SI) | Mant_rounded_S;
assign Fflags_SO = {NV_OP_S,Div_Zero_S,Exp_OF_S,Exp_UF_S,In_Exact_S}; 
endmodule 
import defs_div_sqrt_mvp::*;
module nrbd_nrsc_mvp
  (
   input logic                                 Clk_CI,
   input logic                                 Rst_RBI,
   input logic                                 Div_start_SI,
   input logic                                 Sqrt_start_SI,
   input logic                                 Start_SI,
   input logic                                 Kill_SI,
   input logic                                 Special_case_SBI,
   input logic                                 Special_case_dly_SBI,
   input logic [C_PC-1:0]                      Precision_ctl_SI,
   input logic [1:0]                           Format_sel_SI,
   input logic [C_MANT_FP64:0]                 Mant_a_DI,
   input logic [C_MANT_FP64:0]                 Mant_b_DI,
   input logic [C_EXP_FP64:0]                  Exp_a_DI,
   input logic [C_EXP_FP64:0]                  Exp_b_DI,
  
   output logic                                Div_enable_SO,
   output logic                                Sqrt_enable_SO,
   output logic                                Full_precision_SO,
   output logic                                FP32_SO,
   output logic                                FP64_SO,
   output logic                                FP16_SO,
   output logic                                FP16ALT_SO,
   output logic                                Ready_SO,
   output logic                                Done_SO,
   output logic  [C_MANT_FP64+4:0]             Mant_z_DO,
   output logic [C_EXP_FP64+1:0]               Exp_z_DO
    );
    logic                                     Div_start_dly_S,Sqrt_start_dly_S;
control_mvp         control_U0
(  .Clk_CI                                   (Clk_CI                          ),
   .Rst_RBI                                  (Rst_RBI                         ),
   .Div_start_SI                             (Div_start_SI                    ),
   .Sqrt_start_SI                            (Sqrt_start_SI                   ),
   .Start_SI                                 (Start_SI                        ),
   .Kill_SI                                  (Kill_SI                         ),
   .Special_case_SBI                         (Special_case_SBI                ),
   .Special_case_dly_SBI                     (Special_case_dly_SBI            ),
   .Precision_ctl_SI                         (Precision_ctl_SI                ),
   .Format_sel_SI                            (Format_sel_SI                   ),
   .Numerator_DI                             (Mant_a_DI                       ),
   .Exp_num_DI                               (Exp_a_DI                        ),
   .Denominator_DI                           (Mant_b_DI                       ),
   .Exp_den_DI                               (Exp_b_DI                        ),
   .Div_start_dly_SO                         (Div_start_dly_S                 ),
   .Sqrt_start_dly_SO                        (Sqrt_start_dly_S                ),
   .Div_enable_SO                            (Div_enable_SO                   ),
   .Sqrt_enable_SO                           (Sqrt_enable_SO                  ),
   .Full_precision_SO                        (Full_precision_SO               ),
   .FP32_SO                                  (FP32_SO                         ),
   .FP64_SO                                  (FP64_SO                         ),
   .FP16_SO                                  (FP16_SO                         ),
   .FP16ALT_SO                               (FP16ALT_SO                      ),
   .Ready_SO                                 (Ready_SO                        ),
   .Done_SO                                  (Done_SO                         ),
   .Mant_result_prenorm_DO                   (Mant_z_DO                       ),
   .Exp_result_prenorm_DO                    (Exp_z_DO                        )
);
endmodule
import defs_div_sqrt_mvp::*;
module preprocess_mvp
  (
   input logic                   Clk_CI,
   input logic                   Rst_RBI,
   input logic                   Div_start_SI,
   input logic                   Sqrt_start_SI,
   input logic                   Ready_SI,
   
   input logic [C_OP_FP64-1:0]   Operand_a_DI,
   input logic [C_OP_FP64-1:0]   Operand_b_DI,
   input logic [C_RM-1:0]        RM_SI,    
   input logic [C_FS-1:0]        Format_sel_SI,  
   
   output logic                  Start_SO,
   output logic [C_EXP_FP64:0]   Exp_a_DO_norm,
   output logic [C_EXP_FP64:0]   Exp_b_DO_norm,
   output logic [C_MANT_FP64:0]  Mant_a_DO_norm,
   output logic [C_MANT_FP64:0]  Mant_b_DO_norm,
   output logic [C_RM-1:0]       RM_dly_SO,
   output logic                  Sign_z_DO,
   output logic                  Inf_a_SO,
   output logic                  Inf_b_SO,
   output logic                  Zero_a_SO,
   output logic                  Zero_b_SO,
   output logic                  NaN_a_SO,
   output logic                  NaN_b_SO,
   output logic                  SNaN_SO,
   output logic                  Special_case_SBO,
   output logic                  Special_case_dly_SBO
   );
   
   logic                         Hb_a_D;
   logic                         Hb_b_D;
   logic [C_EXP_FP64-1:0]        Exp_a_D;
   logic [C_EXP_FP64-1:0]        Exp_b_D;
   logic [C_MANT_FP64-1:0]       Mant_a_NonH_D;
   logic [C_MANT_FP64-1:0]       Mant_b_NonH_D;
   logic [C_MANT_FP64:0]         Mant_a_D;
   logic [C_MANT_FP64:0]         Mant_b_D;
   
   
   
   logic                      Sign_a_D,Sign_b_D;
   logic                      Start_S;
     always_comb
       begin
         case(Format_sel_SI)
           2'b00:
             begin
               Sign_a_D = Operand_a_DI[C_OP_FP32-1];
               Sign_b_D = Operand_b_DI[C_OP_FP32-1];
               Exp_a_D  = {3'h0, Operand_a_DI[C_OP_FP32-2:C_MANT_FP32]};
               Exp_b_D  = {3'h0, Operand_b_DI[C_OP_FP32-2:C_MANT_FP32]};
               Mant_a_NonH_D = {Operand_a_DI[C_MANT_FP32-1:0],29'h0};
               Mant_b_NonH_D = {Operand_b_DI[C_MANT_FP32-1:0],29'h0};
             end
           2'b01:
             begin
               Sign_a_D = Operand_a_DI[C_OP_FP64-1];
               Sign_b_D = Operand_b_DI[C_OP_FP64-1];
               Exp_a_D  = Operand_a_DI[C_OP_FP64-2:C_MANT_FP64];
               Exp_b_D  = Operand_b_DI[C_OP_FP64-2:C_MANT_FP64];
               Mant_a_NonH_D = Operand_a_DI[C_MANT_FP64-1:0];
               Mant_b_NonH_D = Operand_b_DI[C_MANT_FP64-1:0];
             end
           2'b10:
             begin
               Sign_a_D = Operand_a_DI[C_OP_FP16-1];
               Sign_b_D = Operand_b_DI[C_OP_FP16-1];
               Exp_a_D  = {6'h00, Operand_a_DI[C_OP_FP16-2:C_MANT_FP16]};
               Exp_b_D  = {6'h00, Operand_b_DI[C_OP_FP16-2:C_MANT_FP16]};
               Mant_a_NonH_D = {Operand_a_DI[C_MANT_FP16-1:0],42'h0};
               Mant_b_NonH_D = {Operand_b_DI[C_MANT_FP16-1:0],42'h0};
             end
           2'b11:
             begin
               Sign_a_D = Operand_a_DI[C_OP_FP16ALT-1];
               Sign_b_D = Operand_b_DI[C_OP_FP16ALT-1];
               Exp_a_D  = {3'h0, Operand_a_DI[C_OP_FP16ALT-2:C_MANT_FP16ALT]};
               Exp_b_D  = {3'h0, Operand_b_DI[C_OP_FP16ALT-2:C_MANT_FP16ALT]};
               Mant_a_NonH_D = {Operand_a_DI[C_MANT_FP16ALT-1:0],45'h0};
               Mant_b_NonH_D = {Operand_b_DI[C_MANT_FP16ALT-1:0],45'h0};
             end
           endcase
       end
   assign Mant_a_D = {Hb_a_D,Mant_a_NonH_D};
   assign Mant_b_D = {Hb_b_D,Mant_b_NonH_D};
   assign Hb_a_D = | Exp_a_D; 
   assign Hb_b_D = | Exp_b_D; 
   assign Start_S= Div_start_SI | Sqrt_start_SI;
   
   
   
   logic               Mant_a_prenorm_zero_S;
   logic               Mant_b_prenorm_zero_S;
   logic               Exp_a_prenorm_zero_S;
   logic               Exp_b_prenorm_zero_S;
   assign Exp_a_prenorm_zero_S = ~Hb_a_D;
   assign Exp_b_prenorm_zero_S = ~Hb_b_D;
   logic               Exp_a_prenorm_Inf_NaN_S;
   logic               Exp_b_prenorm_Inf_NaN_S;
   logic               Mant_a_prenorm_QNaN_S;
   logic               Mant_a_prenorm_SNaN_S;
   logic               Mant_b_prenorm_QNaN_S;
   logic               Mant_b_prenorm_SNaN_S;
   assign Mant_a_prenorm_QNaN_S=Mant_a_NonH_D[C_MANT_FP64-1]&&(~(|Mant_a_NonH_D[C_MANT_FP64-2:0]));
   assign Mant_a_prenorm_SNaN_S=(~Mant_a_NonH_D[C_MANT_FP64-1])&&((|Mant_a_NonH_D[C_MANT_FP64-2:0]));
   assign Mant_b_prenorm_QNaN_S=Mant_b_NonH_D[C_MANT_FP64-1]&&(~(|Mant_b_NonH_D[C_MANT_FP64-2:0]));
   assign Mant_b_prenorm_SNaN_S=(~Mant_b_NonH_D[C_MANT_FP64-1])&&((|Mant_b_NonH_D[C_MANT_FP64-2:0]));
     always_comb
       begin
         case(Format_sel_SI)
           2'b00:
             begin
               Mant_a_prenorm_zero_S=(Operand_a_DI[C_MANT_FP32-1:0] == C_MANT_ZERO_FP32);
               Mant_b_prenorm_zero_S=(Operand_b_DI[C_MANT_FP32-1:0] == C_MANT_ZERO_FP32);
               Exp_a_prenorm_Inf_NaN_S=(Operand_a_DI[C_OP_FP32-2:C_MANT_FP32] == C_EXP_INF_FP32);
               Exp_b_prenorm_Inf_NaN_S=(Operand_b_DI[C_OP_FP32-2:C_MANT_FP32] == C_EXP_INF_FP32);
             end
           2'b01:
             begin
               Mant_a_prenorm_zero_S=(Operand_a_DI[C_MANT_FP64-1:0] == C_MANT_ZERO_FP64);
               Mant_b_prenorm_zero_S=(Operand_b_DI[C_MANT_FP64-1:0] == C_MANT_ZERO_FP64);
               Exp_a_prenorm_Inf_NaN_S=(Operand_a_DI[C_OP_FP64-2:C_MANT_FP64] == C_EXP_INF_FP64);
               Exp_b_prenorm_Inf_NaN_S=(Operand_b_DI[C_OP_FP64-2:C_MANT_FP64] == C_EXP_INF_FP64);
             end
           2'b10:
             begin
               Mant_a_prenorm_zero_S=(Operand_a_DI[C_MANT_FP16-1:0] == C_MANT_ZERO_FP16);
               Mant_b_prenorm_zero_S=(Operand_b_DI[C_MANT_FP16-1:0] == C_MANT_ZERO_FP16);
               Exp_a_prenorm_Inf_NaN_S=(Operand_a_DI[C_OP_FP16-2:C_MANT_FP16] == C_EXP_INF_FP16);
               Exp_b_prenorm_Inf_NaN_S=(Operand_b_DI[C_OP_FP16-2:C_MANT_FP16] == C_EXP_INF_FP16);
             end
           2'b11:
             begin
               Mant_a_prenorm_zero_S=(Operand_a_DI[C_MANT_FP16ALT-1:0] == C_MANT_ZERO_FP16ALT);
               Mant_b_prenorm_zero_S=(Operand_b_DI[C_MANT_FP16ALT-1:0] == C_MANT_ZERO_FP16ALT);
               Exp_a_prenorm_Inf_NaN_S=(Operand_a_DI[C_OP_FP16ALT-2:C_MANT_FP16ALT] == C_EXP_INF_FP16ALT);
               Exp_b_prenorm_Inf_NaN_S=(Operand_b_DI[C_OP_FP16ALT-2:C_MANT_FP16ALT] == C_EXP_INF_FP16ALT);
             end
           endcase
       end
   logic               Zero_a_SN,Zero_a_SP;
   logic               Zero_b_SN,Zero_b_SP;
   logic               Inf_a_SN,Inf_a_SP;
   logic               Inf_b_SN,Inf_b_SP;
   logic               NaN_a_SN,NaN_a_SP;
   logic               NaN_b_SN,NaN_b_SP;
   logic               SNaN_SN,SNaN_SP;
   assign Zero_a_SN = (Start_S&&Ready_SI)?(Exp_a_prenorm_zero_S&&Mant_a_prenorm_zero_S):Zero_a_SP;
   assign Zero_b_SN = (Start_S&&Ready_SI)?(Exp_b_prenorm_zero_S&&Mant_b_prenorm_zero_S):Zero_b_SP;
   assign Inf_a_SN = (Start_S&&Ready_SI)?(Exp_a_prenorm_Inf_NaN_S&&Mant_a_prenorm_zero_S):Inf_a_SP;
   assign Inf_b_SN = (Start_S&&Ready_SI)?(Exp_b_prenorm_Inf_NaN_S&&Mant_b_prenorm_zero_S):Inf_b_SP;
   assign NaN_a_SN = (Start_S&&Ready_SI)?(Exp_a_prenorm_Inf_NaN_S&&(~Mant_a_prenorm_zero_S)):NaN_a_SP;
   assign NaN_b_SN = (Start_S&&Ready_SI)?(Exp_b_prenorm_Inf_NaN_S&&(~Mant_b_prenorm_zero_S)):NaN_b_SP;
   assign SNaN_SN = (Start_S&&Ready_SI) ? ((Mant_a_prenorm_SNaN_S&&NaN_a_SN) | (Mant_b_prenorm_SNaN_S&&NaN_b_SN)) : SNaN_SP;
   always_ff @(posedge Clk_CI, negedge Rst_RBI)
     begin
        if(~Rst_RBI)
          begin
            Zero_a_SP <='0;
            Zero_b_SP <='0;
            Inf_a_SP <='0;
            Inf_b_SP <='0;
            NaN_a_SP <='0;
            NaN_b_SP <='0;
            SNaN_SP <= '0;
          end
        else
         begin
           Inf_a_SP <=Inf_a_SN;
           Inf_b_SP <=Inf_b_SN;
           Zero_a_SP <=Zero_a_SN;
           Zero_b_SP <=Zero_b_SN;
           NaN_a_SP <=NaN_a_SN;
           NaN_b_SP <=NaN_b_SN;
           SNaN_SP <= SNaN_SN;
         end
      end
   
   
   
   assign Special_case_SBO=(~{(Div_start_SI)?(Zero_a_SN | Zero_b_SN |  Inf_a_SN | Inf_b_SN | NaN_a_SN | NaN_b_SN): (Zero_a_SN | Inf_a_SN | NaN_a_SN | Sign_a_D) })&&(Start_S&&Ready_SI);
   always_ff @(posedge Clk_CI, negedge Rst_RBI)
     begin
       if(~Rst_RBI)
          begin
            Special_case_dly_SBO <= '0;
          end
       else if((Start_S&&Ready_SI))
         begin
            Special_case_dly_SBO <= Special_case_SBO;
         end
       else if(Special_case_dly_SBO)
         begin
         Special_case_dly_SBO <= 1'b1;
         end
      else
         begin
            Special_case_dly_SBO <= '0;
         end
    end
   
   
   
   logic                   Sign_z_DN;
   logic                   Sign_z_DP;
   always_comb
     begin
       if(Div_start_SI&&Ready_SI)
           Sign_z_DN = Sign_a_D ^ Sign_b_D;
       else if(Sqrt_start_SI&&Ready_SI)
           Sign_z_DN = Sign_a_D;
       else
           Sign_z_DN = Sign_z_DP;
    end
   always_ff @(posedge Clk_CI, negedge Rst_RBI)
     begin
       if(~Rst_RBI)
          begin
            Sign_z_DP <= '0;
          end
       else
         begin
            Sign_z_DP <= Sign_z_DN;
         end
    end
   logic [C_RM-1:0]                  RM_DN;
   logic [C_RM-1:0]                  RM_DP;
   always_comb
     begin
       if(Start_S&&Ready_SI)
           RM_DN = RM_SI;
       else
           RM_DN = RM_DP;
    end
   always_ff @(posedge Clk_CI, negedge Rst_RBI)
     begin
       if(~Rst_RBI)
          begin
            RM_DP <= '0;
          end
       else
         begin
            RM_DP <= RM_DN;
         end
    end
   assign RM_dly_SO = RM_DP;
   logic [5:0]                  Mant_leadingOne_a, Mant_leadingOne_b;
   logic                        Mant_zero_S_a,Mant_zero_S_b;
  lzc #(
    .WIDTH ( C_MANT_FP64+1 ),
    .MODE  ( 1             )
  ) LOD_Ua (
    .in_i    ( Mant_a_D          ),
    .cnt_o   ( Mant_leadingOne_a ),
    .empty_o ( Mant_zero_S_a     )
  );
   logic [C_MANT_FP64:0]            Mant_a_norm_DN,Mant_a_norm_DP;
   assign  Mant_a_norm_DN = ((Start_S&&Ready_SI))?(Mant_a_D<<(Mant_leadingOne_a)):Mant_a_norm_DP;
   always_ff @(posedge Clk_CI, negedge Rst_RBI)
     begin
        if(~Rst_RBI)
          begin
            Mant_a_norm_DP <= '0;
          end
        else
          begin
            Mant_a_norm_DP<=Mant_a_norm_DN;
          end
     end
   logic [C_EXP_FP64:0]            Exp_a_norm_DN,Exp_a_norm_DP;
   assign  Exp_a_norm_DN = ((Start_S&&Ready_SI))?(Exp_a_D-Mant_leadingOne_a+(|Mant_leadingOne_a)):Exp_a_norm_DP;  
   always_ff @(posedge Clk_CI, negedge Rst_RBI)
     begin
        if(~Rst_RBI)
          begin
            Exp_a_norm_DP <= '0;
          end
        else
          begin
            Exp_a_norm_DP<=Exp_a_norm_DN;
          end
     end
  lzc #(
    .WIDTH ( C_MANT_FP64+1 ),
    .MODE  ( 1             )
  ) LOD_Ub (
    .in_i    ( Mant_b_D          ),
    .cnt_o   ( Mant_leadingOne_b ),
    .empty_o ( Mant_zero_S_b     )
  );
   logic [C_MANT_FP64:0]            Mant_b_norm_DN,Mant_b_norm_DP;
   assign  Mant_b_norm_DN = ((Start_S&&Ready_SI))?(Mant_b_D<<(Mant_leadingOne_b)):Mant_b_norm_DP;
   always_ff @(posedge Clk_CI, negedge Rst_RBI)
     begin
        if(~Rst_RBI)
          begin
            Mant_b_norm_DP <= '0;
          end
        else
          begin
            Mant_b_norm_DP<=Mant_b_norm_DN;
          end
     end
   logic [C_EXP_FP64:0]            Exp_b_norm_DN,Exp_b_norm_DP;
   assign  Exp_b_norm_DN = ((Start_S&&Ready_SI))?(Exp_b_D-Mant_leadingOne_b+(|Mant_leadingOne_b)):Exp_b_norm_DP; 
   always_ff @(posedge Clk_CI, negedge Rst_RBI)
     begin
        if(~Rst_RBI)
          begin
            Exp_b_norm_DP <= '0;
          end
        else
          begin
            Exp_b_norm_DP<=Exp_b_norm_DN;
          end
     end
   
   
   
   assign Start_SO=Start_S;
   assign Exp_a_DO_norm=Exp_a_norm_DP;
   assign Exp_b_DO_norm=Exp_b_norm_DP;
   assign Mant_a_DO_norm=Mant_a_norm_DP;
   assign Mant_b_DO_norm=Mant_b_norm_DP;
   assign Sign_z_DO=Sign_z_DP;
   assign Inf_a_SO=Inf_a_SP;
   assign Inf_b_SO=Inf_b_SP;
   assign Zero_a_SO=Zero_a_SP;
   assign Zero_b_SO=Zero_b_SP;
   assign NaN_a_SO=NaN_a_SP;
   assign NaN_b_SO=NaN_b_SP;
   assign SNaN_SO=SNaN_SP;
endmodule
module fpnew_cast_multi #(
  parameter fpnew_pkg::fmt_logic_t   FpFmtConfig  = '1,
  parameter fpnew_pkg::ifmt_logic_t  IntFmtConfig = '1,
  
  parameter int unsigned             NumPipeRegs = 0,
  parameter fpnew_pkg::pipe_config_t PipeConfig  = fpnew_pkg::BEFORE,
  parameter type                     TagType     = logic,
  parameter type                     AuxType     = logic,
  
  localparam int unsigned WIDTH = fpnew_pkg::maximum(fpnew_pkg::max_fp_width(FpFmtConfig),
                                                     fpnew_pkg::max_int_width(IntFmtConfig)),
  localparam int unsigned NUM_FORMATS = fpnew_pkg::NUM_FP_FORMATS
) (
  input  logic                   clk_i,
  input  logic                   rst_ni,
  
  input  logic [WIDTH-1:0]       operands_i, 
  input  logic [NUM_FORMATS-1:0] is_boxed_i, 
  input  fpnew_pkg::roundmode_e  rnd_mode_i,
  input  fpnew_pkg::operation_e  op_i,
  input  logic                   op_mod_i,
  input  fpnew_pkg::fp_format_e  src_fmt_i,
  input  fpnew_pkg::fp_format_e  dst_fmt_i,
  input  fpnew_pkg::int_format_e int_fmt_i,
  input  TagType                 tag_i,
  input  AuxType                 aux_i,
  
  input  logic                   in_valid_i,
  output logic                   in_ready_o,
  input  logic                   flush_i,
  
  output logic [WIDTH-1:0]       result_o,
  output fpnew_pkg::status_t     status_o,
  output logic                   extension_bit_o,
  output TagType                 tag_o,
  output AuxType                 aux_o,
  
  output logic                   out_valid_o,
  input  logic                   out_ready_i,
  
  output logic                   busy_o
);
  
  
  
  localparam int unsigned NUM_INT_FORMATS = fpnew_pkg::NUM_INT_FORMATS;
  localparam int unsigned MAX_INT_WIDTH   = fpnew_pkg::max_int_width(IntFmtConfig);
  localparam fpnew_pkg::fp_encoding_t SUPER_FORMAT = fpnew_pkg::super_format(FpFmtConfig);
  localparam int unsigned SUPER_EXP_BITS = SUPER_FORMAT.exp_bits;
  localparam int unsigned SUPER_MAN_BITS = SUPER_FORMAT.man_bits;
  localparam int unsigned SUPER_BIAS     = 2**(SUPER_EXP_BITS - 1) - 1;
  
  localparam int unsigned INT_MAN_WIDTH = fpnew_pkg::maximum(SUPER_MAN_BITS + 1, MAX_INT_WIDTH);
  
  localparam int unsigned LZC_RESULT_WIDTH = $clog2(INT_MAN_WIDTH);
  
  
  localparam int unsigned INT_EXP_WIDTH = fpnew_pkg::maximum($clog2(MAX_INT_WIDTH),
      fpnew_pkg::maximum(SUPER_EXP_BITS, $clog2(SUPER_BIAS + SUPER_MAN_BITS))) + 1;
  
  localparam NUM_INP_REGS = PipeConfig == fpnew_pkg::BEFORE
                            ? NumPipeRegs
                            : (PipeConfig == fpnew_pkg::DISTRIBUTED
                               ? ((NumPipeRegs + 1) / 3) 
                               : 0); 
  localparam NUM_MID_REGS = PipeConfig == fpnew_pkg::INSIDE
                          ? NumPipeRegs
                          : (PipeConfig == fpnew_pkg::DISTRIBUTED
                             ? ((NumPipeRegs + 2) / 3) 
                             : 0); 
  localparam NUM_OUT_REGS = PipeConfig == fpnew_pkg::AFTER
                            ? NumPipeRegs
                            : (PipeConfig == fpnew_pkg::DISTRIBUTED
                               ? (NumPipeRegs / 3) 
                               : 0); 
  
  
  
  
  logic [WIDTH-1:0]       operands_q;
  logic [NUM_FORMATS-1:0] is_boxed_q;
  logic                   op_mod_q;
  fpnew_pkg::fp_format_e  src_fmt_q;
  fpnew_pkg::fp_format_e  dst_fmt_q;
  fpnew_pkg::int_format_e int_fmt_q;
  
  logic                   [0:NUM_INP_REGS][WIDTH-1:0]       inp_pipe_operands_q;
  logic                   [0:NUM_INP_REGS][NUM_FORMATS-1:0] inp_pipe_is_boxed_q;
  fpnew_pkg::roundmode_e  [0:NUM_INP_REGS]                  inp_pipe_rnd_mode_q;
  fpnew_pkg::operation_e  [0:NUM_INP_REGS]                  inp_pipe_op_q;
  logic                   [0:NUM_INP_REGS]                  inp_pipe_op_mod_q;
  fpnew_pkg::fp_format_e  [0:NUM_INP_REGS]                  inp_pipe_src_fmt_q;
  fpnew_pkg::fp_format_e  [0:NUM_INP_REGS]                  inp_pipe_dst_fmt_q;
  fpnew_pkg::int_format_e [0:NUM_INP_REGS]                  inp_pipe_int_fmt_q;
  TagType                 [0:NUM_INP_REGS]                  inp_pipe_tag_q;
  AuxType                 [0:NUM_INP_REGS]                  inp_pipe_aux_q;
  logic                   [0:NUM_INP_REGS]                  inp_pipe_valid_q;
  
  logic [0:NUM_INP_REGS] inp_pipe_ready;
  
  assign inp_pipe_operands_q[0] = operands_i;
  assign inp_pipe_is_boxed_q[0] = is_boxed_i;
  assign inp_pipe_rnd_mode_q[0] = rnd_mode_i;
  assign inp_pipe_op_q[0]       = op_i;
  assign inp_pipe_op_mod_q[0]   = op_mod_i;
  assign inp_pipe_src_fmt_q[0]  = src_fmt_i;
  assign inp_pipe_dst_fmt_q[0]  = dst_fmt_i;
  assign inp_pipe_int_fmt_q[0]  = int_fmt_i;
  assign inp_pipe_tag_q[0]      = tag_i;
  assign inp_pipe_aux_q[0]      = aux_i;
  assign inp_pipe_valid_q[0]    = in_valid_i;
  
  assign in_ready_o = inp_pipe_ready[0];
  
  for (genvar i = 0; i < NUM_INP_REGS; i++) begin : gen_input_pipeline
    
    logic reg_ena;
    
    
    
    assign inp_pipe_ready[i] = inp_pipe_ready[i+1] | ~inp_pipe_valid_q[i+1];
    
    
                           
                         
                            
  always_ff @(posedge (clk_i) or negedge (rst_ni)) begin                 
    if (!rst_ni) begin                                                   
      inp_pipe_valid_q[i+1] <= (1'b0);                                              
    end else begin                                                         
      inp_pipe_valid_q[i+1] <= (flush_i) ? (1'b0) : (inp_pipe_ready[i]) ? (inp_pipe_valid_q[i]) : (inp_pipe_valid_q[i+1]);       
    end                                                                    
  end
    
    assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
    
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_operands_q[i+1] <= ('0);                        
    end else begin                                   
      inp_pipe_operands_q[i+1] <= (reg_ena) ? (inp_pipe_operands_q[i]) : (inp_pipe_operands_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_is_boxed_q[i+1] <= ('0);                        
    end else begin                                   
      inp_pipe_is_boxed_q[i+1] <= (reg_ena) ? (inp_pipe_is_boxed_q[i]) : (inp_pipe_is_boxed_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_rnd_mode_q[i+1] <= (fpnew_pkg::RNE);                        
    end else begin                                   
      inp_pipe_rnd_mode_q[i+1] <= (reg_ena) ? (inp_pipe_rnd_mode_q[i]) : (inp_pipe_rnd_mode_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_op_q[i+1] <= (fpnew_pkg::FMADD);                        
    end else begin                                   
      inp_pipe_op_q[i+1] <= (reg_ena) ? (inp_pipe_op_q[i]) : (inp_pipe_op_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_op_mod_q[i+1] <= ('0);                        
    end else begin                                   
      inp_pipe_op_mod_q[i+1] <= (reg_ena) ? (inp_pipe_op_mod_q[i]) : (inp_pipe_op_mod_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_src_fmt_q[i+1] <= (fpnew_pkg::fp_format_e'(0));                        
    end else begin                                   
      inp_pipe_src_fmt_q[i+1] <= (reg_ena) ? (inp_pipe_src_fmt_q[i]) : (inp_pipe_src_fmt_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_dst_fmt_q[i+1] <= (fpnew_pkg::fp_format_e'(0));                        
    end else begin                                   
      inp_pipe_dst_fmt_q[i+1] <= (reg_ena) ? (inp_pipe_dst_fmt_q[i]) : (inp_pipe_dst_fmt_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_int_fmt_q[i+1] <= (fpnew_pkg::int_format_e'(0));                        
    end else begin                                   
      inp_pipe_int_fmt_q[i+1] <= (reg_ena) ? (inp_pipe_int_fmt_q[i]) : (inp_pipe_int_fmt_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_tag_q[i+1] <= (TagType'('0));                        
    end else begin                                   
      inp_pipe_tag_q[i+1] <= (reg_ena) ? (inp_pipe_tag_q[i]) : (inp_pipe_tag_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_aux_q[i+1] <= (AuxType'('0));                        
    end else begin                                   
      inp_pipe_aux_q[i+1] <= (reg_ena) ? (inp_pipe_aux_q[i]) : (inp_pipe_aux_q[i+1]);               
    end                                              
  end
  end
  
  assign operands_q = inp_pipe_operands_q[NUM_INP_REGS];
  assign is_boxed_q = inp_pipe_is_boxed_q[NUM_INP_REGS];
  assign op_mod_q   = inp_pipe_op_mod_q[NUM_INP_REGS];
  assign src_fmt_q  = inp_pipe_src_fmt_q[NUM_INP_REGS];
  assign dst_fmt_q  = inp_pipe_dst_fmt_q[NUM_INP_REGS];
  assign int_fmt_q  = inp_pipe_int_fmt_q[NUM_INP_REGS];
  
  
  
  logic src_is_int, dst_is_int; 
  assign src_is_int = (inp_pipe_op_q[NUM_INP_REGS] == fpnew_pkg::I2F);
  assign dst_is_int = (inp_pipe_op_q[NUM_INP_REGS] == fpnew_pkg::F2I);
  logic [INT_MAN_WIDTH-1:0] encoded_mant; 
  logic        [NUM_FORMATS-1:0]                    fmt_sign;
  logic signed [NUM_FORMATS-1:0][INT_EXP_WIDTH-1:0] fmt_exponent;
  logic        [NUM_FORMATS-1:0][INT_MAN_WIDTH-1:0] fmt_mantissa;
  logic signed [NUM_FORMATS-1:0][INT_EXP_WIDTH-1:0] fmt_shift_compensation; 
  fpnew_pkg::fp_info_t [NUM_FORMATS-1:0] info;
  logic [NUM_INT_FORMATS-1:0][INT_MAN_WIDTH-1:0] ifmt_input_val;
  logic                                          int_sign;
  logic [INT_MAN_WIDTH-1:0]                      int_value, int_mantissa;
  
  for (genvar fmt = 0; fmt < int'(NUM_FORMATS); fmt++) begin : fmt_init_inputs
    
    localparam int unsigned FP_WIDTH = fpnew_pkg::fp_width(fpnew_pkg::fp_format_e'(fmt));
    localparam int unsigned EXP_BITS = fpnew_pkg::exp_bits(fpnew_pkg::fp_format_e'(fmt));
    localparam int unsigned MAN_BITS = fpnew_pkg::man_bits(fpnew_pkg::fp_format_e'(fmt));
    if (FpFmtConfig[fmt]) begin : active_format
      
      fpnew_classifier #(
        .FpFormat    ( fpnew_pkg::fp_format_e'(fmt) ),
        .NumOperands ( 1                            )
      ) i_fpnew_classifier (
        .operands_i ( operands_q[FP_WIDTH-1:0] ),
        .is_boxed_i ( is_boxed_q[fmt]          ),
        .info_o     ( info[fmt]                )
      );
      assign fmt_sign[fmt]     = operands_q[FP_WIDTH-1];
      assign fmt_exponent[fmt] = signed'({1'b0, operands_q[MAN_BITS+:EXP_BITS]});
      assign fmt_mantissa[fmt] = {info[fmt].is_normal, operands_q[MAN_BITS-1:0]}; 
      
      assign fmt_shift_compensation[fmt] = signed'(INT_MAN_WIDTH - 1 - MAN_BITS);
    end else begin : inactive_format
      assign info[fmt]                   = '{default: fpnew_pkg::DONT_CARE}; 
      assign fmt_sign[fmt]               = fpnew_pkg::DONT_CARE;             
      assign fmt_exponent[fmt]           = '{default: fpnew_pkg::DONT_CARE}; 
      assign fmt_mantissa[fmt]           = '{default: fpnew_pkg::DONT_CARE}; 
      assign fmt_shift_compensation[fmt] = '{default: fpnew_pkg::DONT_CARE}; 
    end
  end
  
  for (genvar ifmt = 0; ifmt < int'(NUM_INT_FORMATS); ifmt++) begin : gen_sign_extend_int
    
    localparam int unsigned INT_WIDTH = fpnew_pkg::int_width(fpnew_pkg::int_format_e'(ifmt));
    if (IntFmtConfig[ifmt]) begin : active_format 
      always_comb begin : sign_ext_input
        
        ifmt_input_val[ifmt]                = '{default: operands_q[INT_WIDTH-1] & ~op_mod_q};
        ifmt_input_val[ifmt][INT_WIDTH-1:0] = operands_q[INT_WIDTH-1:0];
      end
    end else begin : inactive_format
      assign ifmt_input_val[ifmt] = '{default: fpnew_pkg::DONT_CARE}; 
    end
  end
  
  assign int_value    = ifmt_input_val[int_fmt_q];
  assign int_sign     = int_value[INT_MAN_WIDTH-1] & ~op_mod_q; 
  assign int_mantissa = int_sign ? unsigned'(-int_value) : int_value; 
  
  assign encoded_mant = src_is_int ? int_mantissa : fmt_mantissa[src_fmt_q];
  
  
  
  logic signed [INT_EXP_WIDTH-1:0] src_bias;      
  logic signed [INT_EXP_WIDTH-1:0] src_exp;       
  logic signed [INT_EXP_WIDTH-1:0] src_subnormal; 
  logic signed [INT_EXP_WIDTH-1:0] src_offset;    
  assign src_bias      = signed'(fpnew_pkg::bias(src_fmt_q));
  assign src_exp       = fmt_exponent[src_fmt_q];
  assign src_subnormal = signed'({1'b0, info[src_fmt_q].is_subnormal});
  assign src_offset    = fmt_shift_compensation[src_fmt_q];
  logic                            input_sign;   
  logic signed [INT_EXP_WIDTH-1:0] input_exp;    
  logic        [INT_MAN_WIDTH-1:0] input_mant;   
  logic                            mant_is_zero; 
  logic signed [INT_EXP_WIDTH-1:0] fp_input_exp;
  logic signed [INT_EXP_WIDTH-1:0] int_input_exp;
  
  logic [LZC_RESULT_WIDTH-1:0] renorm_shamt;     
  logic [LZC_RESULT_WIDTH:0]   renorm_shamt_sgn; 
  
  lzc #(
    .WIDTH ( INT_MAN_WIDTH ),
    .MODE  ( 1             ) 
  ) i_lzc (
    .in_i    ( encoded_mant ),
    .cnt_o   ( renorm_shamt ),
    .empty_o ( mant_is_zero )
  );
  assign renorm_shamt_sgn = signed'({1'b0, renorm_shamt});
  
  assign input_sign = src_is_int ? int_sign : fmt_sign[src_fmt_q];
  
  assign input_mant = encoded_mant << renorm_shamt;
  
  assign fp_input_exp  = signed'(src_exp + src_subnormal - src_bias -
                                 renorm_shamt_sgn + src_offset); 
  assign int_input_exp = signed'(INT_MAN_WIDTH - 1 - renorm_shamt_sgn);
  assign input_exp     = src_is_int ? int_input_exp : fp_input_exp;
  logic signed [INT_EXP_WIDTH-1:0] destination_exp;  
  
  assign destination_exp = input_exp + signed'(fpnew_pkg::bias(dst_fmt_q));
  
  
  
  
  logic                            input_sign_q;
  logic signed [INT_EXP_WIDTH-1:0] input_exp_q;
  logic [INT_MAN_WIDTH-1:0]        input_mant_q;
  logic signed [INT_EXP_WIDTH-1:0] destination_exp_q;
  logic                            src_is_int_q;
  logic                            dst_is_int_q;
  fpnew_pkg::fp_info_t             info_q;
  logic                            mant_is_zero_q;
  logic                            op_mod_q2;
  fpnew_pkg::roundmode_e           rnd_mode_q;
  fpnew_pkg::fp_format_e           src_fmt_q2;
  fpnew_pkg::fp_format_e           dst_fmt_q2;
  fpnew_pkg::int_format_e          int_fmt_q2;
  
  logic                   [0:NUM_MID_REGS]                    mid_pipe_input_sign_q;
  logic signed            [0:NUM_MID_REGS][INT_EXP_WIDTH-1:0] mid_pipe_input_exp_q;
  logic                   [0:NUM_MID_REGS][INT_MAN_WIDTH-1:0] mid_pipe_input_mant_q;
  logic signed            [0:NUM_MID_REGS][INT_EXP_WIDTH-1:0] mid_pipe_dest_exp_q;
  logic                   [0:NUM_MID_REGS]                    mid_pipe_src_is_int_q;
  logic                   [0:NUM_MID_REGS]                    mid_pipe_dst_is_int_q;
  fpnew_pkg::fp_info_t    [0:NUM_MID_REGS]                    mid_pipe_info_q;
  logic                   [0:NUM_MID_REGS]                    mid_pipe_mant_zero_q;
  logic                   [0:NUM_MID_REGS]                    mid_pipe_op_mod_q;
  fpnew_pkg::roundmode_e  [0:NUM_MID_REGS]                    mid_pipe_rnd_mode_q;
  fpnew_pkg::fp_format_e  [0:NUM_MID_REGS]                    mid_pipe_src_fmt_q;
  fpnew_pkg::fp_format_e  [0:NUM_MID_REGS]                    mid_pipe_dst_fmt_q;
  fpnew_pkg::int_format_e [0:NUM_MID_REGS]                    mid_pipe_int_fmt_q;
  TagType                 [0:NUM_MID_REGS]                    mid_pipe_tag_q;
  AuxType                 [0:NUM_MID_REGS]                    mid_pipe_aux_q;
  logic                   [0:NUM_MID_REGS]                    mid_pipe_valid_q;
  
  logic [0:NUM_MID_REGS] mid_pipe_ready;
  
  assign mid_pipe_input_sign_q[0] = input_sign;
  assign mid_pipe_input_exp_q[0]  = input_exp;
  assign mid_pipe_input_mant_q[0] = input_mant;
  assign mid_pipe_dest_exp_q[0]   = destination_exp;
  assign mid_pipe_src_is_int_q[0] = src_is_int;
  assign mid_pipe_dst_is_int_q[0] = dst_is_int;
  assign mid_pipe_info_q[0]       = info[src_fmt_q];
  assign mid_pipe_mant_zero_q[0]  = mant_is_zero;
  assign mid_pipe_op_mod_q[0]     = op_mod_q;
  assign mid_pipe_rnd_mode_q[0]   = inp_pipe_rnd_mode_q[NUM_INP_REGS];
  assign mid_pipe_src_fmt_q[0]    = src_fmt_q;
  assign mid_pipe_dst_fmt_q[0]    = dst_fmt_q;
  assign mid_pipe_int_fmt_q[0]    = int_fmt_q;
  assign mid_pipe_tag_q[0]        = inp_pipe_tag_q[NUM_INP_REGS];
  assign mid_pipe_aux_q[0]        = inp_pipe_aux_q[NUM_INP_REGS];
  assign mid_pipe_valid_q[0]      = inp_pipe_valid_q[NUM_INP_REGS];
  
  assign inp_pipe_ready[NUM_INP_REGS] = mid_pipe_ready[0];
  
  for (genvar i = 0; i < NUM_MID_REGS; i++) begin : gen_inside_pipeline
    
    logic reg_ena;
    
    
    
    assign mid_pipe_ready[i] = mid_pipe_ready[i+1] | ~mid_pipe_valid_q[i+1];
    
    
                           
                         
                            
  always_ff @(posedge (clk_i) or negedge (rst_ni)) begin                 
    if (!rst_ni) begin                                                   
      mid_pipe_valid_q[i+1] <= (1'b0);                                              
    end else begin                                                         
      mid_pipe_valid_q[i+1] <= (flush_i) ? (1'b0) : (mid_pipe_ready[i]) ? (mid_pipe_valid_q[i]) : (mid_pipe_valid_q[i+1]);       
    end                                                                    
  end
    
    assign reg_ena = mid_pipe_ready[i] & mid_pipe_valid_q[i];
    
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_input_sign_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_input_sign_q[i+1] <= (reg_ena) ? (mid_pipe_input_sign_q[i]) : (mid_pipe_input_sign_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_input_exp_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_input_exp_q[i+1] <= (reg_ena) ? (mid_pipe_input_exp_q[i]) : (mid_pipe_input_exp_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_input_mant_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_input_mant_q[i+1] <= (reg_ena) ? (mid_pipe_input_mant_q[i]) : (mid_pipe_input_mant_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_dest_exp_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_dest_exp_q[i+1] <= (reg_ena) ? (mid_pipe_dest_exp_q[i]) : (mid_pipe_dest_exp_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_src_is_int_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_src_is_int_q[i+1] <= (reg_ena) ? (mid_pipe_src_is_int_q[i]) : (mid_pipe_src_is_int_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_dst_is_int_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_dst_is_int_q[i+1] <= (reg_ena) ? (mid_pipe_dst_is_int_q[i]) : (mid_pipe_dst_is_int_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_info_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_info_q[i+1] <= (reg_ena) ? (mid_pipe_info_q[i]) : (mid_pipe_info_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_mant_zero_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_mant_zero_q[i+1] <= (reg_ena) ? (mid_pipe_mant_zero_q[i]) : (mid_pipe_mant_zero_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_op_mod_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_op_mod_q[i+1] <= (reg_ena) ? (mid_pipe_op_mod_q[i]) : (mid_pipe_op_mod_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_rnd_mode_q[i+1] <= (fpnew_pkg::RNE);                        
    end else begin                                   
      mid_pipe_rnd_mode_q[i+1] <= (reg_ena) ? (mid_pipe_rnd_mode_q[i]) : (mid_pipe_rnd_mode_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_src_fmt_q[i+1] <= (fpnew_pkg::fp_format_e'(0));                        
    end else begin                                   
      mid_pipe_src_fmt_q[i+1] <= (reg_ena) ? (mid_pipe_src_fmt_q[i]) : (mid_pipe_src_fmt_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_dst_fmt_q[i+1] <= (fpnew_pkg::fp_format_e'(0));                        
    end else begin                                   
      mid_pipe_dst_fmt_q[i+1] <= (reg_ena) ? (mid_pipe_dst_fmt_q[i]) : (mid_pipe_dst_fmt_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_int_fmt_q[i+1] <= (fpnew_pkg::int_format_e'(0));                        
    end else begin                                   
      mid_pipe_int_fmt_q[i+1] <= (reg_ena) ? (mid_pipe_int_fmt_q[i]) : (mid_pipe_int_fmt_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_tag_q[i+1] <= (TagType'('0));                        
    end else begin                                   
      mid_pipe_tag_q[i+1] <= (reg_ena) ? (mid_pipe_tag_q[i]) : (mid_pipe_tag_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_aux_q[i+1] <= (AuxType'('0));                        
    end else begin                                   
      mid_pipe_aux_q[i+1] <= (reg_ena) ? (mid_pipe_aux_q[i]) : (mid_pipe_aux_q[i+1]);               
    end                                              
  end
  end
  
  assign input_sign_q      = mid_pipe_input_sign_q[NUM_MID_REGS];
  assign input_exp_q       = mid_pipe_input_exp_q[NUM_MID_REGS];
  assign input_mant_q      = mid_pipe_input_mant_q[NUM_MID_REGS];
  assign destination_exp_q = mid_pipe_dest_exp_q[NUM_MID_REGS];
  assign src_is_int_q      = mid_pipe_src_is_int_q[NUM_MID_REGS];
  assign dst_is_int_q      = mid_pipe_dst_is_int_q[NUM_MID_REGS];
  assign info_q            = mid_pipe_info_q[NUM_MID_REGS];
  assign mant_is_zero_q    = mid_pipe_mant_zero_q[NUM_MID_REGS];
  assign op_mod_q2         = mid_pipe_op_mod_q[NUM_MID_REGS];
  assign rnd_mode_q        = mid_pipe_rnd_mode_q[NUM_MID_REGS];
  assign src_fmt_q2        = mid_pipe_src_fmt_q[NUM_MID_REGS];
  assign dst_fmt_q2        = mid_pipe_dst_fmt_q[NUM_MID_REGS];
  assign int_fmt_q2        = mid_pipe_int_fmt_q[NUM_MID_REGS];
  
  
  
  logic [INT_EXP_WIDTH-1:0] final_exp;        
  logic [2*INT_MAN_WIDTH:0]  preshift_mant;    
  logic [2*INT_MAN_WIDTH:0]  destination_mant; 
  logic [SUPER_MAN_BITS-1:0] final_mant;       
  logic [MAX_INT_WIDTH-1:0]  final_int;        
  logic [$clog2(INT_MAN_WIDTH+1)-1:0] denorm_shamt; 
  logic [1:0] fp_round_sticky_bits, int_round_sticky_bits, round_sticky_bits;
  logic       of_before_round, uf_before_round;
  
  always_comb begin : cast_value
    
    final_exp       = unsigned'(destination_exp_q); 
    preshift_mant   = '0;  
    denorm_shamt    = SUPER_MAN_BITS - fpnew_pkg::man_bits(dst_fmt_q2); 
    of_before_round = 1'b0;
    uf_before_round = 1'b0;
    
    preshift_mant = input_mant_q << (INT_MAN_WIDTH + 1);
    
    if (dst_is_int_q) begin
      
      denorm_shamt = unsigned'(MAX_INT_WIDTH - 1 - input_exp_q);
      
      if (input_exp_q >= signed'(fpnew_pkg::int_width(int_fmt_q2) - 1 + op_mod_q2)) begin
        denorm_shamt    = '0; 
        of_before_round = 1'b1;
      
      end else if (input_exp_q < -1) begin
        denorm_shamt    = MAX_INT_WIDTH + 1; 
        uf_before_round = 1'b1;
      end
    
    end else begin
      
      if ((destination_exp_q >= signed'(2**fpnew_pkg::exp_bits(dst_fmt_q2))-1) ||
          (~src_is_int_q && info_q.is_inf)) begin
        final_exp       = unsigned'(2**fpnew_pkg::exp_bits(dst_fmt_q2)-2); 
        preshift_mant   = '1;                           
        of_before_round = 1'b1;
      
      end else if (destination_exp_q < 1 &&
                   destination_exp_q >= -signed'(fpnew_pkg::man_bits(dst_fmt_q2))) begin
        final_exp       = '0; 
        denorm_shamt    = unsigned'(denorm_shamt + 1 - destination_exp_q); 
        uf_before_round = 1'b1;
      
      end else if (destination_exp_q < -signed'(fpnew_pkg::man_bits(dst_fmt_q2))) begin
        final_exp       = '0; 
        denorm_shamt    = unsigned'(denorm_shamt + 2 + fpnew_pkg::man_bits(dst_fmt_q2)); 
        uf_before_round = 1'b1;
      end
    end
  end
  localparam NUM_FP_STICKY  = 2 * INT_MAN_WIDTH - SUPER_MAN_BITS - 1; 
  localparam NUM_INT_STICKY = 2 * INT_MAN_WIDTH - MAX_INT_WIDTH; 
  
  assign destination_mant = preshift_mant >> denorm_shamt;
  
  assign {final_mant, fp_round_sticky_bits[1]} =
      destination_mant[2*INT_MAN_WIDTH-1-:SUPER_MAN_BITS+1];
  assign {final_int, int_round_sticky_bits[1]} = destination_mant[2*INT_MAN_WIDTH-:MAX_INT_WIDTH+1];
  
  assign fp_round_sticky_bits[0]  = (| {destination_mant[NUM_FP_STICKY-1:0]});
  assign int_round_sticky_bits[0] = (| {destination_mant[NUM_INT_STICKY-1:0]});
  
  assign round_sticky_bits = dst_is_int_q ? int_round_sticky_bits : fp_round_sticky_bits;
  
  
  
  logic [WIDTH-1:0] pre_round_abs;  
  logic             of_after_round; 
  logic             uf_after_round; 
  logic [NUM_FORMATS-1:0][WIDTH-1:0] fmt_pre_round_abs; 
  logic [NUM_FORMATS-1:0]            fmt_of_after_round;
  logic [NUM_FORMATS-1:0]            fmt_uf_after_round;
  logic [NUM_INT_FORMATS-1:0][WIDTH-1:0] ifmt_pre_round_abs; 
  logic             rounded_sign;
  logic [WIDTH-1:0] rounded_abs; 
  logic             result_true_zero;
  logic [WIDTH-1:0] rounded_int_res; 
  logic             rounded_int_res_zero; 
  
  for (genvar fmt = 0; fmt < int'(NUM_FORMATS); fmt++) begin : gen_res_assemble
    
    localparam int unsigned EXP_BITS = fpnew_pkg::exp_bits(fpnew_pkg::fp_format_e'(fmt));
    localparam int unsigned MAN_BITS = fpnew_pkg::man_bits(fpnew_pkg::fp_format_e'(fmt));
    if (FpFmtConfig[fmt]) begin : active_format
      always_comb begin : assemble_result
        fmt_pre_round_abs[fmt] = {final_exp[EXP_BITS-1:0], final_mant[MAN_BITS-1:0]}; 
      end
    end else begin : inactive_format
      assign fmt_pre_round_abs[fmt] = '{default: fpnew_pkg::DONT_CARE};
    end
  end
  
  for (genvar ifmt = 0; ifmt < int'(NUM_INT_FORMATS); ifmt++) begin : gen_int_res_sign_ext
    
    localparam int unsigned INT_WIDTH = fpnew_pkg::int_width(fpnew_pkg::int_format_e'(ifmt));
    if (IntFmtConfig[ifmt]) begin : active_format
      always_comb begin : assemble_result
        
        ifmt_pre_round_abs[ifmt]                = '{default: final_int[INT_WIDTH-1]};
        ifmt_pre_round_abs[ifmt][INT_WIDTH-1:0] = final_int[INT_WIDTH-1:0];
      end
    end else begin : inactive_format
      assign ifmt_pre_round_abs[ifmt] = '{default: fpnew_pkg::DONT_CARE};
    end
  end
  
  assign pre_round_abs = dst_is_int_q ? ifmt_pre_round_abs[int_fmt_q2] : fmt_pre_round_abs[dst_fmt_q2];
  fpnew_rounding #(
    .AbsWidth ( WIDTH )
  ) i_fpnew_rounding (
    .abs_value_i             ( pre_round_abs     ),
    .sign_i                  ( input_sign_q      ), 
    .round_sticky_bits_i     ( round_sticky_bits ),
    .rnd_mode_i              ( rnd_mode_q        ),
    .effective_subtraction_i ( 1'b0              ), 
    .abs_rounded_o           ( rounded_abs       ),
    .sign_o                  ( rounded_sign      ),
    .exact_zero_o            ( result_true_zero  )
  );
  logic [NUM_FORMATS-1:0][WIDTH-1:0] fmt_result;
  
  for (genvar fmt = 0; fmt < int'(NUM_FORMATS); fmt++) begin : gen_sign_inject
    
    localparam int unsigned FP_WIDTH = fpnew_pkg::fp_width(fpnew_pkg::fp_format_e'(fmt));
    localparam int unsigned EXP_BITS = fpnew_pkg::exp_bits(fpnew_pkg::fp_format_e'(fmt));
    localparam int unsigned MAN_BITS = fpnew_pkg::man_bits(fpnew_pkg::fp_format_e'(fmt));
    if (FpFmtConfig[fmt]) begin : active_format
      always_comb begin : post_process
        
        fmt_uf_after_round[fmt] = rounded_abs[EXP_BITS+MAN_BITS-1:MAN_BITS] == '0; 
        fmt_of_after_round[fmt] = rounded_abs[EXP_BITS+MAN_BITS-1:MAN_BITS] == '1; 
        
        fmt_result[fmt]               = '1;
        fmt_result[fmt][FP_WIDTH-1:0] = src_is_int_q & mant_is_zero_q
                                        ? '0
                                        : {rounded_sign, rounded_abs[EXP_BITS+MAN_BITS-1:0]};
      end
    end else begin : inactive_format
      assign fmt_uf_after_round[fmt] = fpnew_pkg::DONT_CARE;
      assign fmt_of_after_round[fmt] = fpnew_pkg::DONT_CARE;
      assign fmt_result[fmt]         = '{default: fpnew_pkg::DONT_CARE};
    end
  end
  
  assign uf_after_round = fmt_uf_after_round[dst_fmt_q2];
  assign of_after_round = fmt_of_after_round[dst_fmt_q2];
  
  assign rounded_int_res      = rounded_sign ? unsigned'(-rounded_abs) : rounded_abs;
  assign rounded_int_res_zero = (rounded_int_res == '0);
  
  
  
  logic [WIDTH-1:0]   fp_special_result;
  fpnew_pkg::status_t fp_special_status;
  logic               fp_result_is_special;
  logic [NUM_FORMATS-1:0][WIDTH-1:0] fmt_special_result;
  
  for (genvar fmt = 0; fmt < int'(NUM_FORMATS); fmt++) begin : gen_special_results
    
    localparam int unsigned FP_WIDTH = fpnew_pkg::fp_width(fpnew_pkg::fp_format_e'(fmt));
    localparam int unsigned EXP_BITS = fpnew_pkg::exp_bits(fpnew_pkg::fp_format_e'(fmt));
    localparam int unsigned MAN_BITS = fpnew_pkg::man_bits(fpnew_pkg::fp_format_e'(fmt));
    localparam logic [EXP_BITS-1:0] QNAN_EXPONENT = '1;
    localparam logic [MAN_BITS-1:0] QNAN_MANTISSA = 2**(MAN_BITS-1);
    if (FpFmtConfig[fmt]) begin : active_format
      always_comb begin : special_results
        logic [FP_WIDTH-1:0] special_res;
        special_res = info_q.is_zero
                      ? input_sign_q << FP_WIDTH-1 
                      : {1'b0, QNAN_EXPONENT, QNAN_MANTISSA}; 
        
        fmt_special_result[fmt]               = '1;
        fmt_special_result[fmt][FP_WIDTH-1:0] = special_res;
      end
    end else begin : inactive_format
      assign fmt_special_result[fmt] = '{default: fpnew_pkg::DONT_CARE};
    end
  end
  
  assign fp_result_is_special = ~src_is_int_q & (info_q.is_zero |
                                                 info_q.is_nan |
                                                 ~info_q.is_boxed);
  
  assign fp_special_status = '{NV: info_q.is_signalling, default: 1'b0};
  
  assign fp_special_result = fmt_special_result[dst_fmt_q2]; 
  
  
  
  logic [WIDTH-1:0]   int_special_result;
  fpnew_pkg::status_t int_special_status;
  logic               int_result_is_special;
  logic [NUM_INT_FORMATS-1:0][WIDTH-1:0] ifmt_special_result;
  
  for (genvar ifmt = 0; ifmt < int'(NUM_INT_FORMATS); ifmt++) begin : gen_special_results_int
    
    localparam int unsigned INT_WIDTH = fpnew_pkg::int_width(fpnew_pkg::int_format_e'(ifmt));
    if (IntFmtConfig[ifmt]) begin : active_format
      always_comb begin : special_results
        automatic logic [INT_WIDTH-1:0] special_res;
        
        special_res[INT_WIDTH-2:0] = '1;       
        special_res[INT_WIDTH-1]   = op_mod_q2; 
        
        if (input_sign_q && !info_q.is_nan)
          special_res = ~special_res;
        
        ifmt_special_result[ifmt]                = '{default: special_res[INT_WIDTH-1]};
        ifmt_special_result[ifmt][INT_WIDTH-1:0] = special_res;
      end
    end else begin : inactive_format
      assign ifmt_special_result[ifmt] = '{default: fpnew_pkg::DONT_CARE};
    end
  end
  
  assign int_result_is_special = info_q.is_nan | info_q.is_inf |
                                 of_before_round | ~info_q.is_boxed |
                                 (input_sign_q & op_mod_q2 & ~rounded_int_res_zero);
  
  assign int_special_status = '{NV: 1'b1, default: 1'b0};
  
  assign int_special_result = ifmt_special_result[int_fmt_q2]; 
  
  
  
  fpnew_pkg::status_t int_regular_status, fp_regular_status;
  logic [WIDTH-1:0]   fp_result, int_result;
  fpnew_pkg::status_t fp_status, int_status;
  assign fp_regular_status.NV = src_is_int_q & (of_before_round | of_after_round); 
  assign fp_regular_status.DZ = 1'b0; 
  assign fp_regular_status.OF = ~src_is_int_q & (~info_q.is_inf & (of_before_round | of_after_round)); 
  assign fp_regular_status.UF = uf_after_round & fp_regular_status.NX;
  assign fp_regular_status.NX = src_is_int_q ? (| fp_round_sticky_bits) 
            : (| fp_round_sticky_bits) | (~info_q.is_inf & (of_before_round | of_after_round));
  assign int_regular_status = '{NX: (| int_round_sticky_bits), default: 1'b0};
  assign fp_result  = fp_result_is_special  ? fp_special_result  : fmt_result[dst_fmt_q2];
  assign fp_status  = fp_result_is_special  ? fp_special_status  : fp_regular_status;
  assign int_result = int_result_is_special ? int_special_result : rounded_int_res;
  assign int_status = int_result_is_special ? int_special_status : int_regular_status;
  
  logic [WIDTH-1:0]   result_d;
  fpnew_pkg::status_t status_d;
  logic               extension_bit;
  
  assign result_d = dst_is_int_q ? int_result : fp_result;
  assign status_d = dst_is_int_q ? int_status : fp_status;
  
  assign extension_bit = dst_is_int_q ? int_result[WIDTH-1] : 1'b1;
  
  
  
  
  logic               [0:NUM_OUT_REGS][WIDTH-1:0] out_pipe_result_q;
  fpnew_pkg::status_t [0:NUM_OUT_REGS]            out_pipe_status_q;
  logic               [0:NUM_OUT_REGS]            out_pipe_ext_bit_q;
  TagType             [0:NUM_OUT_REGS]            out_pipe_tag_q;
  AuxType             [0:NUM_OUT_REGS]            out_pipe_aux_q;
  logic               [0:NUM_OUT_REGS]            out_pipe_valid_q;
  
  logic [0:NUM_OUT_REGS] out_pipe_ready;
  
  assign out_pipe_result_q[0]  = result_d;
  assign out_pipe_status_q[0]  = status_d;
  assign out_pipe_ext_bit_q[0] = extension_bit;
  assign out_pipe_tag_q[0]     = mid_pipe_tag_q[NUM_MID_REGS];
  assign out_pipe_aux_q[0]     = mid_pipe_aux_q[NUM_MID_REGS];
  assign out_pipe_valid_q[0]   = mid_pipe_valid_q[NUM_MID_REGS];
  
  assign mid_pipe_ready[NUM_MID_REGS] = out_pipe_ready[0];
  
  for (genvar i = 0; i < NUM_OUT_REGS; i++) begin : gen_output_pipeline
    
    logic reg_ena;
    
    
    
    assign out_pipe_ready[i] = out_pipe_ready[i+1] | ~out_pipe_valid_q[i+1];
    
    
                           
                         
                            
  always_ff @(posedge (clk_i) or negedge (rst_ni)) begin                 
    if (!rst_ni) begin                                                   
      out_pipe_valid_q[i+1] <= (1'b0);                                              
    end else begin                                                         
      out_pipe_valid_q[i+1] <= (flush_i) ? (1'b0) : (out_pipe_ready[i]) ? (out_pipe_valid_q[i]) : (out_pipe_valid_q[i+1]);       
    end                                                                    
  end
    
    assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
    
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_result_q[i+1] <= ('0);                        
    end else begin                                   
      out_pipe_result_q[i+1] <= (reg_ena) ? (out_pipe_result_q[i]) : (out_pipe_result_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_status_q[i+1] <= ('0);                        
    end else begin                                   
      out_pipe_status_q[i+1] <= (reg_ena) ? (out_pipe_status_q[i]) : (out_pipe_status_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_ext_bit_q[i+1] <= ('0);                        
    end else begin                                   
      out_pipe_ext_bit_q[i+1] <= (reg_ena) ? (out_pipe_ext_bit_q[i]) : (out_pipe_ext_bit_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_tag_q[i+1] <= (TagType'('0));                        
    end else begin                                   
      out_pipe_tag_q[i+1] <= (reg_ena) ? (out_pipe_tag_q[i]) : (out_pipe_tag_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_aux_q[i+1] <= (AuxType'('0));                        
    end else begin                                   
      out_pipe_aux_q[i+1] <= (reg_ena) ? (out_pipe_aux_q[i]) : (out_pipe_aux_q[i+1]);               
    end                                              
  end
  end
  
  assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
  
  assign result_o        = out_pipe_result_q[NUM_OUT_REGS];
  assign status_o        = out_pipe_status_q[NUM_OUT_REGS];
  assign extension_bit_o = out_pipe_ext_bit_q[NUM_OUT_REGS];
  assign tag_o           = out_pipe_tag_q[NUM_OUT_REGS];
  assign aux_o           = out_pipe_aux_q[NUM_OUT_REGS];
  assign out_valid_o     = out_pipe_valid_q[NUM_OUT_REGS];
  assign busy_o          = (| {inp_pipe_valid_q, mid_pipe_valid_q, out_pipe_valid_q});
endmodule
module fpnew_classifier #(
  parameter fpnew_pkg::fp_format_e   FpFormat = fpnew_pkg::fp_format_e'(0),
  parameter int unsigned             NumOperands = 1,
  
  localparam int unsigned WIDTH = fpnew_pkg::fp_width(FpFormat)
) (
  input  logic                [NumOperands-1:0][WIDTH-1:0] operands_i,
  input  logic                [NumOperands-1:0]            is_boxed_i,
  output fpnew_pkg::fp_info_t [NumOperands-1:0]            info_o
);
  localparam int unsigned EXP_BITS = fpnew_pkg::exp_bits(FpFormat);
  localparam int unsigned MAN_BITS = fpnew_pkg::man_bits(FpFormat);
  
  typedef struct packed {
    logic                sign;
    logic [EXP_BITS-1:0] exponent;
    logic [MAN_BITS-1:0] mantissa;
  } fp_t;
  
  for (genvar op = 0; op < int'(NumOperands); op++) begin : gen_num_values
    fp_t value;
    logic is_boxed;
    logic is_normal;
    logic is_inf;
    logic is_nan;
    logic is_signalling;
    logic is_quiet;
    logic is_zero;
    logic is_subnormal;
    
    
    
    always_comb begin : classify_input
      value         = operands_i[op];
      is_boxed      = is_boxed_i[op];
      is_normal     = is_boxed && (value.exponent != '0) && (value.exponent != '1);
      is_zero       = is_boxed && (value.exponent == '0) && (value.mantissa == '0);
      is_subnormal  = is_boxed && (value.exponent == '0) && !is_zero;
      is_inf        = is_boxed && ((value.exponent == '1) && (value.mantissa == '0));
      is_nan        = !is_boxed || ((value.exponent == '1) && (value.mantissa != '0));
      is_signalling = is_boxed && is_nan && (value.mantissa[MAN_BITS-1] == 1'b0);
      is_quiet      = is_nan && !is_signalling;
      
      info_o[op].is_normal     = is_normal;
      info_o[op].is_subnormal  = is_subnormal;
      info_o[op].is_zero       = is_zero;
      info_o[op].is_inf        = is_inf;
      info_o[op].is_nan        = is_nan;
      info_o[op].is_signalling = is_signalling;
      info_o[op].is_quiet      = is_quiet;
      info_o[op].is_boxed      = is_boxed;
    end
  end
endmodule
                                      
module fpnew_divsqrt_multi #(
  parameter fpnew_pkg::fmt_logic_t   FpFmtConfig  = '1,
  
  parameter int unsigned             NumPipeRegs = 0,
  parameter fpnew_pkg::pipe_config_t PipeConfig  = fpnew_pkg::AFTER,
  parameter type                     TagType     = logic,
  parameter type                     AuxType     = logic,
  
  localparam int unsigned WIDTH       = fpnew_pkg::max_fp_width(FpFmtConfig),
  localparam int unsigned NUM_FORMATS = fpnew_pkg::NUM_FP_FORMATS
) (
  input  logic                        clk_i,
  input  logic                        rst_ni,
  
  input  logic [1:0][WIDTH-1:0]       operands_i, 
  input  logic [NUM_FORMATS-1:0][1:0] is_boxed_i, 
  input  fpnew_pkg::roundmode_e       rnd_mode_i,
  input  fpnew_pkg::operation_e       op_i,
  input  fpnew_pkg::fp_format_e       dst_fmt_i,
  input  TagType                      tag_i,
  input  AuxType                      aux_i,
  
  input  logic                        in_valid_i,
  output logic                        in_ready_o,
  input  logic                        flush_i,
  
  output logic [WIDTH-1:0]            result_o,
  output fpnew_pkg::status_t          status_o,
  output logic                        extension_bit_o,
  output TagType                      tag_o,
  output AuxType                      aux_o,
  
  output logic                        out_valid_o,
  input  logic                        out_ready_i,
  
  output logic                        busy_o
);
  
  
  
  
  localparam NUM_INP_REGS = (PipeConfig == fpnew_pkg::BEFORE)
                            ? NumPipeRegs
                            : (PipeConfig == fpnew_pkg::DISTRIBUTED
                               ? (NumPipeRegs / 2) 
                               : 0); 
  localparam NUM_OUT_REGS = (PipeConfig == fpnew_pkg::AFTER || PipeConfig == fpnew_pkg::INSIDE)
                            ? NumPipeRegs
                            : (PipeConfig == fpnew_pkg::DISTRIBUTED
                               ? ((NumPipeRegs + 1) / 2) 
                               : 0); 
  
  
  
  
  logic [1:0][WIDTH-1:0] operands_q;
  fpnew_pkg::roundmode_e rnd_mode_q;
  fpnew_pkg::operation_e op_q;
  fpnew_pkg::fp_format_e dst_fmt_q;
  logic                  in_valid_q;
  
  logic                  [0:NUM_INP_REGS][1:0][WIDTH-1:0]       inp_pipe_operands_q;
  fpnew_pkg::roundmode_e [0:NUM_INP_REGS]                       inp_pipe_rnd_mode_q;
  fpnew_pkg::operation_e [0:NUM_INP_REGS]                       inp_pipe_op_q;
  fpnew_pkg::fp_format_e [0:NUM_INP_REGS]                       inp_pipe_dst_fmt_q;
  TagType                [0:NUM_INP_REGS]                       inp_pipe_tag_q;
  AuxType                [0:NUM_INP_REGS]                       inp_pipe_aux_q;
  logic                  [0:NUM_INP_REGS]                       inp_pipe_valid_q;
  
  logic [0:NUM_INP_REGS] inp_pipe_ready;
  
  assign inp_pipe_operands_q[0] = operands_i;
  assign inp_pipe_rnd_mode_q[0] = rnd_mode_i;
  assign inp_pipe_op_q[0]       = op_i;
  assign inp_pipe_dst_fmt_q[0]  = dst_fmt_i;
  assign inp_pipe_tag_q[0]      = tag_i;
  assign inp_pipe_aux_q[0]      = aux_i;
  assign inp_pipe_valid_q[0]    = in_valid_i;
  
  assign in_ready_o = inp_pipe_ready[0];
  
  for (genvar i = 0; i < NUM_INP_REGS; i++) begin : gen_input_pipeline
    
    logic reg_ena;
    
    
    
    assign inp_pipe_ready[i] = inp_pipe_ready[i+1] | ~inp_pipe_valid_q[i+1];
    
    
                           
                         
                            
  always_ff @(posedge (clk_i) or negedge (rst_ni)) begin                 
    if (!rst_ni) begin                                                   
      inp_pipe_valid_q[i+1] <= (1'b0);                                              
    end else begin                                                         
      inp_pipe_valid_q[i+1] <= (flush_i) ? (1'b0) : (inp_pipe_ready[i]) ? (inp_pipe_valid_q[i]) : (inp_pipe_valid_q[i+1]);       
    end                                                                    
  end
    
    assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
    
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_operands_q[i+1] <= ('0);                        
    end else begin                                   
      inp_pipe_operands_q[i+1] <= (reg_ena) ? (inp_pipe_operands_q[i]) : (inp_pipe_operands_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_rnd_mode_q[i+1] <= (fpnew_pkg::RNE);                        
    end else begin                                   
      inp_pipe_rnd_mode_q[i+1] <= (reg_ena) ? (inp_pipe_rnd_mode_q[i]) : (inp_pipe_rnd_mode_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_op_q[i+1] <= (fpnew_pkg::FMADD);                        
    end else begin                                   
      inp_pipe_op_q[i+1] <= (reg_ena) ? (inp_pipe_op_q[i]) : (inp_pipe_op_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_dst_fmt_q[i+1] <= (fpnew_pkg::fp_format_e'(0));                        
    end else begin                                   
      inp_pipe_dst_fmt_q[i+1] <= (reg_ena) ? (inp_pipe_dst_fmt_q[i]) : (inp_pipe_dst_fmt_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_tag_q[i+1] <= (TagType'('0));                        
    end else begin                                   
      inp_pipe_tag_q[i+1] <= (reg_ena) ? (inp_pipe_tag_q[i]) : (inp_pipe_tag_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_aux_q[i+1] <= (AuxType'('0));                        
    end else begin                                   
      inp_pipe_aux_q[i+1] <= (reg_ena) ? (inp_pipe_aux_q[i]) : (inp_pipe_aux_q[i+1]);               
    end                                              
  end
  end
  
  assign operands_q = inp_pipe_operands_q[NUM_INP_REGS];
  assign rnd_mode_q = inp_pipe_rnd_mode_q[NUM_INP_REGS];
  assign op_q       = inp_pipe_op_q[NUM_INP_REGS];
  assign dst_fmt_q  = inp_pipe_dst_fmt_q[NUM_INP_REGS];
  assign in_valid_q = inp_pipe_valid_q[NUM_INP_REGS];
  
  
  
  logic [1:0]       divsqrt_fmt;
  logic [1:0][63:0] divsqrt_operands; 
  logic             input_is_fp8;
  
  always_comb begin : translate_fmt
    unique case (dst_fmt_q)
      fpnew_pkg::FP32:    divsqrt_fmt = 2'b00;
      fpnew_pkg::FP64:    divsqrt_fmt = 2'b01;
      fpnew_pkg::FP16:    divsqrt_fmt = 2'b10;
      fpnew_pkg::FP16ALT: divsqrt_fmt = 2'b11;
      default:            divsqrt_fmt = 2'b10; 
    endcase
    
    input_is_fp8 = FpFmtConfig[fpnew_pkg::FP8] & (dst_fmt_q == fpnew_pkg::FP8);
    
    divsqrt_operands[0] = input_is_fp8 ? operands_q[0] << 8 : operands_q[0];
    divsqrt_operands[1] = input_is_fp8 ? operands_q[1] << 8 : operands_q[1];
  end
  
  
  
  logic in_ready;               
  logic div_valid, sqrt_valid;  
  logic unit_ready, unit_done;  
  logic op_starting;            
  logic out_valid, out_ready;   
  logic hold_result;            
  logic data_is_held;           
  logic unit_busy;              
  
  typedef enum logic [1:0] {IDLE, BUSY, HOLD} fsm_state_e;
  fsm_state_e state_q, state_d;
  
  assign inp_pipe_ready[NUM_INP_REGS] = in_ready;
  
  assign div_valid   = in_valid_q & (op_q == fpnew_pkg::DIV) & in_ready & ~flush_i;
  assign sqrt_valid  = in_valid_q & (op_q != fpnew_pkg::DIV) & in_ready & ~flush_i;
  assign op_starting = div_valid | sqrt_valid;
  
  always_comb begin : flag_fsm
    
    in_ready     = 1'b0;
    out_valid    = 1'b0;
    hold_result  = 1'b0;
    data_is_held = 1'b0;
    unit_busy    = 1'b0;
    state_d      = state_q;
    unique case (state_q)
      
      IDLE: begin
        in_ready = 1'b1; 
        if (in_valid_q && unit_ready) begin 
          state_d = BUSY; 
        end
      end
      
      BUSY: begin
        unit_busy = 1'b1; 
        
        if (unit_done) begin
          out_valid = 1'b1; 
          
          if (out_ready) begin
            state_d = IDLE; 
            if (in_valid_q && unit_ready) begin 
              in_ready = 1'b1; 
              state_d  = BUSY; 
            end
          
          end else begin
            hold_result = 1'b1; 
            state_d     = HOLD; 
          end
        end
      end
      
      HOLD: begin
        unit_busy    = 1'b1; 
        data_is_held = 1'b1; 
        out_valid    = 1'b1; 
        
        if (out_ready) begin
          state_d = IDLE; 
          if (in_valid_q && unit_ready) begin 
            in_ready = 1'b1; 
            state_d  = BUSY; 
          end
        end
      end
      
      default: state_d = IDLE;
    endcase
    
    if (flush_i) begin
      unit_busy = 1'b0; 
      out_valid = 1'b0; 
      state_d   = IDLE; 
    end
  end
  
  
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      state_q <= (IDLE);                        
    end else begin                                   
      state_q <= (state_d);                                  
    end                                              
  end
  
  logic result_is_fp8_q;
  TagType result_tag_q;
  AuxType result_aux_q;
  
  
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      result_is_fp8_q <= ('0);                        
    end else begin                                   
      result_is_fp8_q <= (op_starting) ? (input_is_fp8) : (result_is_fp8_q);               
    end                                              
  end
  
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      result_tag_q <= ('0);                        
    end else begin                                   
      result_tag_q <= (op_starting) ? (inp_pipe_tag_q[NUM_INP_REGS]) : (result_tag_q);               
    end                                              
  end
  
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      result_aux_q <= ('0);                        
    end else begin                                   
      result_aux_q <= (op_starting) ? (inp_pipe_aux_q[NUM_INP_REGS]) : (result_aux_q);               
    end                                              
  end
  
  
  
  logic [63:0]        unit_result;
  logic [WIDTH-1:0]   adjusted_result, held_result_q;
  fpnew_pkg::status_t unit_status, held_status_q;
  div_sqrt_top_mvp i_divsqrt_lei (
   .Clk_CI           ( clk_i               ),
   .Rst_RBI          ( rst_ni              ),
   .Div_start_SI     ( div_valid           ),
   .Sqrt_start_SI    ( sqrt_valid          ),
   .Operand_a_DI     ( divsqrt_operands[0] ),
   .Operand_b_DI     ( divsqrt_operands[1] ),
   .RM_SI            ( rnd_mode_q          ),
   .Precision_ctl_SI ( '0                  ),
   .Format_sel_SI    ( divsqrt_fmt         ),
   .Kill_SI          ( flush_i             ),
   .Result_DO        ( unit_result         ),
   .Fflags_SO        ( unit_status         ),
   .Ready_SO         ( unit_ready          ),
   .Done_SO          ( unit_done           )
  );
  
  assign adjusted_result = result_is_fp8_q ? unit_result >> 8 : unit_result;
  
  
  always_ff @(posedge (clk_i)) begin   
    held_result_q <= (hold_result) ? (adjusted_result) : (held_result_q);   
  end
  
  always_ff @(posedge (clk_i)) begin   
    held_status_q <= (hold_result) ? (unit_status) : (held_status_q);   
  end
  
  
  
  logic [WIDTH-1:0]   result_d;
  fpnew_pkg::status_t status_d;
  
  assign result_d = data_is_held ? held_result_q : adjusted_result;
  assign status_d = data_is_held ? held_status_q : unit_status;
  
  
  
  
  logic               [0:NUM_OUT_REGS][WIDTH-1:0] out_pipe_result_q;
  fpnew_pkg::status_t [0:NUM_OUT_REGS]            out_pipe_status_q;
  TagType             [0:NUM_OUT_REGS]            out_pipe_tag_q;
  AuxType             [0:NUM_OUT_REGS]            out_pipe_aux_q;
  logic               [0:NUM_OUT_REGS]            out_pipe_valid_q;
  
  logic [0:NUM_OUT_REGS] out_pipe_ready;
  
  assign out_pipe_result_q[0] = result_d;
  assign out_pipe_status_q[0] = status_d;
  assign out_pipe_tag_q[0]    = result_tag_q;
  assign out_pipe_aux_q[0]    = result_aux_q;
  assign out_pipe_valid_q[0]  = out_valid;
  
  assign out_ready = out_pipe_ready[0];
  
  for (genvar i = 0; i < NUM_OUT_REGS; i++) begin : gen_output_pipeline
    
    logic reg_ena;
    
    
    
    assign out_pipe_ready[i] = out_pipe_ready[i+1] | ~out_pipe_valid_q[i+1];
    
    
                           
                         
                            
  always_ff @(posedge (clk_i) or negedge (rst_ni)) begin                 
    if (!rst_ni) begin                                                   
      out_pipe_valid_q[i+1] <= (1'b0);                                              
    end else begin                                                         
      out_pipe_valid_q[i+1] <= (flush_i) ? (1'b0) : (out_pipe_ready[i]) ? (out_pipe_valid_q[i]) : (out_pipe_valid_q[i+1]);       
    end                                                                    
  end
    
    assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
    
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_result_q[i+1] <= ('0);                        
    end else begin                                   
      out_pipe_result_q[i+1] <= (reg_ena) ? (out_pipe_result_q[i]) : (out_pipe_result_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_status_q[i+1] <= ('0);                        
    end else begin                                   
      out_pipe_status_q[i+1] <= (reg_ena) ? (out_pipe_status_q[i]) : (out_pipe_status_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_tag_q[i+1] <= (TagType'('0));                        
    end else begin                                   
      out_pipe_tag_q[i+1] <= (reg_ena) ? (out_pipe_tag_q[i]) : (out_pipe_tag_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_aux_q[i+1] <= (AuxType'('0));                        
    end else begin                                   
      out_pipe_aux_q[i+1] <= (reg_ena) ? (out_pipe_aux_q[i]) : (out_pipe_aux_q[i+1]);               
    end                                              
  end
  end
  
  assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
  
  assign result_o        = out_pipe_result_q[NUM_OUT_REGS];
  assign status_o        = out_pipe_status_q[NUM_OUT_REGS];
  assign extension_bit_o = 1'b1; 
  assign tag_o           = out_pipe_tag_q[NUM_OUT_REGS];
  assign aux_o           = out_pipe_aux_q[NUM_OUT_REGS];
  assign out_valid_o     = out_pipe_valid_q[NUM_OUT_REGS];
  assign busy_o          = (| {inp_pipe_valid_q, unit_busy, out_pipe_valid_q});
endmodule
                                      
module fpnew_fma_multi #(
  parameter fpnew_pkg::fmt_logic_t   FpFmtConfig = '1,
  parameter int unsigned             NumPipeRegs = 0,
  parameter fpnew_pkg::pipe_config_t PipeConfig  = fpnew_pkg::BEFORE,
  parameter type                     TagType     = logic,
  parameter type                     AuxType     = logic,
  
  localparam int unsigned WIDTH       = fpnew_pkg::max_fp_width(FpFmtConfig),
  localparam int unsigned NUM_FORMATS = fpnew_pkg::NUM_FP_FORMATS
) (
  input  logic                        clk_i,
  input  logic                        rst_ni,
  
  input  logic [2:0][WIDTH-1:0]       operands_i, 
  input  logic [NUM_FORMATS-1:0][2:0] is_boxed_i, 
  input  fpnew_pkg::roundmode_e       rnd_mode_i,
  input  fpnew_pkg::operation_e       op_i,
  input  logic                        op_mod_i,
  input  fpnew_pkg::fp_format_e       src_fmt_i, 
  input  fpnew_pkg::fp_format_e       dst_fmt_i, 
  input  TagType                      tag_i,
  input  AuxType                      aux_i,
  
  input  logic                        in_valid_i,
  output logic                        in_ready_o,
  input  logic                        flush_i,
  
  output logic [WIDTH-1:0]            result_o,
  output fpnew_pkg::status_t          status_o,
  output logic                        extension_bit_o,
  output TagType                      tag_o,
  output AuxType                      aux_o,
  
  output logic                        out_valid_o,
  input  logic                        out_ready_i,
  
  output logic                        busy_o
);
  
  
  
  
  localparam fpnew_pkg::fp_encoding_t SUPER_FORMAT = fpnew_pkg::super_format(FpFmtConfig);
  localparam int unsigned SUPER_EXP_BITS = SUPER_FORMAT.exp_bits;
  localparam int unsigned SUPER_MAN_BITS = SUPER_FORMAT.man_bits;
  
  localparam int unsigned PRECISION_BITS = SUPER_MAN_BITS + 1;
  
  localparam int unsigned LOWER_SUM_WIDTH  = 2 * PRECISION_BITS + 3;
  localparam int unsigned LZC_RESULT_WIDTH = $clog2(LOWER_SUM_WIDTH);
  
  
  
  localparam int unsigned EXP_WIDTH = fpnew_pkg::maximum(SUPER_EXP_BITS + 2, LZC_RESULT_WIDTH);
  
  localparam int unsigned SHIFT_AMOUNT_WIDTH = $clog2(3 * PRECISION_BITS + 3);
  
  localparam NUM_INP_REGS = PipeConfig == fpnew_pkg::BEFORE
                            ? NumPipeRegs
                            : (PipeConfig == fpnew_pkg::DISTRIBUTED
                               ? ((NumPipeRegs + 1) / 3) 
                               : 0); 
  localparam NUM_MID_REGS = PipeConfig == fpnew_pkg::INSIDE
                          ? NumPipeRegs
                          : (PipeConfig == fpnew_pkg::DISTRIBUTED
                             ? ((NumPipeRegs + 2) / 3) 
                             : 0); 
  localparam NUM_OUT_REGS = PipeConfig == fpnew_pkg::AFTER
                            ? NumPipeRegs
                            : (PipeConfig == fpnew_pkg::DISTRIBUTED
                               ? (NumPipeRegs / 3) 
                               : 0); 
  
  
  
  typedef struct packed {
    logic                      sign;
    logic [SUPER_EXP_BITS-1:0] exponent;
    logic [SUPER_MAN_BITS-1:0] mantissa;
  } fp_t;
  
  
  
  
  logic [2:0][WIDTH-1:0] operands_q;
  fpnew_pkg::fp_format_e src_fmt_q;
  fpnew_pkg::fp_format_e dst_fmt_q;
  
  logic                  [0:NUM_INP_REGS][2:0][WIDTH-1:0]       inp_pipe_operands_q;
  logic                  [0:NUM_INP_REGS][NUM_FORMATS-1:0][2:0] inp_pipe_is_boxed_q;
  fpnew_pkg::roundmode_e [0:NUM_INP_REGS]                       inp_pipe_rnd_mode_q;
  fpnew_pkg::operation_e [0:NUM_INP_REGS]                       inp_pipe_op_q;
  logic                  [0:NUM_INP_REGS]                       inp_pipe_op_mod_q;
  fpnew_pkg::fp_format_e [0:NUM_INP_REGS]                       inp_pipe_src_fmt_q;
  fpnew_pkg::fp_format_e [0:NUM_INP_REGS]                       inp_pipe_dst_fmt_q;
  TagType                [0:NUM_INP_REGS]                       inp_pipe_tag_q;
  AuxType                [0:NUM_INP_REGS]                       inp_pipe_aux_q;
  logic                  [0:NUM_INP_REGS]                       inp_pipe_valid_q;
  
  logic [0:NUM_INP_REGS] inp_pipe_ready;
  
  assign inp_pipe_operands_q[0] = operands_i;
  assign inp_pipe_is_boxed_q[0] = is_boxed_i;
  assign inp_pipe_rnd_mode_q[0] = rnd_mode_i;
  assign inp_pipe_op_q[0]       = op_i;
  assign inp_pipe_op_mod_q[0]   = op_mod_i;
  assign inp_pipe_src_fmt_q[0]  = src_fmt_i;
  assign inp_pipe_dst_fmt_q[0]  = dst_fmt_i;
  assign inp_pipe_tag_q[0]      = tag_i;
  assign inp_pipe_aux_q[0]      = aux_i;
  assign inp_pipe_valid_q[0]    = in_valid_i;
  
  assign in_ready_o = inp_pipe_ready[0];
  
  for (genvar i = 0; i < NUM_INP_REGS; i++) begin : gen_input_pipeline
    
    logic reg_ena;
    
    
    
    assign inp_pipe_ready[i] = inp_pipe_ready[i+1] | ~inp_pipe_valid_q[i+1];
    
    
                           
                         
                            
  always_ff @(posedge (clk_i) or negedge (rst_ni)) begin                 
    if (!rst_ni) begin                                                   
      inp_pipe_valid_q[i+1] <= (1'b0);                                              
    end else begin                                                         
      inp_pipe_valid_q[i+1] <= (flush_i) ? (1'b0) : (inp_pipe_ready[i]) ? (inp_pipe_valid_q[i]) : (inp_pipe_valid_q[i+1]);       
    end                                                                    
  end
    
    assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
    
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_operands_q[i+1] <= ('0);                        
    end else begin                                   
      inp_pipe_operands_q[i+1] <= (reg_ena) ? (inp_pipe_operands_q[i]) : (inp_pipe_operands_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_is_boxed_q[i+1] <= ('0);                        
    end else begin                                   
      inp_pipe_is_boxed_q[i+1] <= (reg_ena) ? (inp_pipe_is_boxed_q[i]) : (inp_pipe_is_boxed_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_rnd_mode_q[i+1] <= (fpnew_pkg::RNE);                        
    end else begin                                   
      inp_pipe_rnd_mode_q[i+1] <= (reg_ena) ? (inp_pipe_rnd_mode_q[i]) : (inp_pipe_rnd_mode_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_op_q[i+1] <= (fpnew_pkg::FMADD);                        
    end else begin                                   
      inp_pipe_op_q[i+1] <= (reg_ena) ? (inp_pipe_op_q[i]) : (inp_pipe_op_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_op_mod_q[i+1] <= ('0);                        
    end else begin                                   
      inp_pipe_op_mod_q[i+1] <= (reg_ena) ? (inp_pipe_op_mod_q[i]) : (inp_pipe_op_mod_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_src_fmt_q[i+1] <= (fpnew_pkg::fp_format_e'(0));                        
    end else begin                                   
      inp_pipe_src_fmt_q[i+1] <= (reg_ena) ? (inp_pipe_src_fmt_q[i]) : (inp_pipe_src_fmt_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_dst_fmt_q[i+1] <= (fpnew_pkg::fp_format_e'(0));                        
    end else begin                                   
      inp_pipe_dst_fmt_q[i+1] <= (reg_ena) ? (inp_pipe_dst_fmt_q[i]) : (inp_pipe_dst_fmt_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_tag_q[i+1] <= (TagType'('0));                        
    end else begin                                   
      inp_pipe_tag_q[i+1] <= (reg_ena) ? (inp_pipe_tag_q[i]) : (inp_pipe_tag_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_aux_q[i+1] <= (AuxType'('0));                        
    end else begin                                   
      inp_pipe_aux_q[i+1] <= (reg_ena) ? (inp_pipe_aux_q[i]) : (inp_pipe_aux_q[i+1]);               
    end                                              
  end
  end
  
  assign operands_q = inp_pipe_operands_q[NUM_INP_REGS];
  assign src_fmt_q  = inp_pipe_src_fmt_q[NUM_INP_REGS];
  assign dst_fmt_q  = inp_pipe_dst_fmt_q[NUM_INP_REGS];
  
  
  
  logic        [NUM_FORMATS-1:0][2:0]                     fmt_sign;
  logic signed [NUM_FORMATS-1:0][2:0][SUPER_EXP_BITS-1:0] fmt_exponent;
  logic        [NUM_FORMATS-1:0][2:0][SUPER_MAN_BITS-1:0] fmt_mantissa;
  fpnew_pkg::fp_info_t [NUM_FORMATS-1:0][2:0] info_q;
  
  for (genvar fmt = 0; fmt < int'(NUM_FORMATS); fmt++) begin : fmt_init_inputs
    
    localparam int unsigned FP_WIDTH = fpnew_pkg::fp_width(fpnew_pkg::fp_format_e'(fmt));
    localparam int unsigned EXP_BITS = fpnew_pkg::exp_bits(fpnew_pkg::fp_format_e'(fmt));
    localparam int unsigned MAN_BITS = fpnew_pkg::man_bits(fpnew_pkg::fp_format_e'(fmt));
    if (FpFmtConfig[fmt]) begin : active_format
      logic [2:0][FP_WIDTH-1:0] trimmed_ops;
      
      fpnew_classifier #(
        .FpFormat    ( fpnew_pkg::fp_format_e'(fmt) ),
        .NumOperands ( 3                            )
      ) i_fpnew_classifier (
        .operands_i ( trimmed_ops                            ),
        .is_boxed_i ( inp_pipe_is_boxed_q[NUM_INP_REGS][fmt] ),
        .info_o     ( info_q[fmt]                            )
      );
      for (genvar op = 0; op < 3; op++) begin : gen_operands
        assign trimmed_ops[op]       = operands_q[op][FP_WIDTH-1:0];
        assign fmt_sign[fmt][op]     = operands_q[op][FP_WIDTH-1];
        assign fmt_exponent[fmt][op] = signed'({1'b0, operands_q[op][MAN_BITS+:EXP_BITS]});
        assign fmt_mantissa[fmt][op] = {info_q[fmt][op].is_normal, operands_q[op][MAN_BITS-1:0]} <<
                                       (SUPER_MAN_BITS - MAN_BITS); 
      end
    end else begin : inactive_format
      assign info_q[fmt]                 = '{default: fpnew_pkg::DONT_CARE}; 
      assign fmt_sign[fmt]               = fpnew_pkg::DONT_CARE;             
      assign fmt_exponent[fmt]           = '{default: fpnew_pkg::DONT_CARE}; 
      assign fmt_mantissa[fmt]           = '{default: fpnew_pkg::DONT_CARE}; 
    end
  end
  fp_t                 operand_a, operand_b, operand_c;
  fpnew_pkg::fp_info_t info_a,    info_b,    info_c;
  
  
  
  
  
  
  
  
  
  
  
  
  always_comb begin : op_select
    
    operand_a = {fmt_sign[src_fmt_q][0], fmt_exponent[src_fmt_q][0], fmt_mantissa[src_fmt_q][0]};
    operand_b = {fmt_sign[src_fmt_q][1], fmt_exponent[src_fmt_q][1], fmt_mantissa[src_fmt_q][1]};
    operand_c = {fmt_sign[dst_fmt_q][2], fmt_exponent[dst_fmt_q][2], fmt_mantissa[dst_fmt_q][2]};
    info_a    = info_q[src_fmt_q][0];
    info_b    = info_q[src_fmt_q][1];
    info_c    = info_q[dst_fmt_q][2];
    
    operand_c.sign = operand_c.sign ^ inp_pipe_op_mod_q[NUM_INP_REGS];
    unique case (inp_pipe_op_q[NUM_INP_REGS])
      fpnew_pkg::FMADD:  ; 
      fpnew_pkg::FNMSUB: operand_a.sign = ~operand_a.sign; 
      fpnew_pkg::ADD: begin 
        operand_a = '{sign: 1'b0, exponent: fpnew_pkg::bias(src_fmt_q), mantissa: '0};
        info_a    = '{is_normal: 1'b1, is_boxed: 1'b1, default: 1'b0}; 
      end
      fpnew_pkg::MUL: begin 
        operand_c = '{sign: 1'b1, exponent: '0, mantissa: '0};
        info_c    = '{is_zero: 1'b1, is_boxed: 1'b1, default: 1'b0}; 
      end
      default: begin 
        operand_a  = '{default: fpnew_pkg::DONT_CARE};
        operand_b  = '{default: fpnew_pkg::DONT_CARE};
        operand_c  = '{default: fpnew_pkg::DONT_CARE};
        info_a     = '{default: fpnew_pkg::DONT_CARE};
        info_b     = '{default: fpnew_pkg::DONT_CARE};
        info_c     = '{default: fpnew_pkg::DONT_CARE};
      end
    endcase
  end
  
  
  
  logic any_operand_inf;
  logic any_operand_nan;
  logic signalling_nan;
  logic effective_subtraction;
  logic tentative_sign;
  
  assign any_operand_inf = (| {info_a.is_inf,        info_b.is_inf,        info_c.is_inf});
  assign any_operand_nan = (| {info_a.is_nan,        info_b.is_nan,        info_c.is_nan});
  assign signalling_nan  = (| {info_a.is_signalling, info_b.is_signalling, info_c.is_signalling});
  
  assign effective_subtraction = operand_a.sign ^ operand_b.sign ^ operand_c.sign;
  
  assign tentative_sign = operand_a.sign ^ operand_b.sign;
  
  
  
  logic [WIDTH-1:0]   special_result;
  fpnew_pkg::status_t special_status;
  logic               result_is_special;
  logic [NUM_FORMATS-1:0][WIDTH-1:0]    fmt_special_result;
  fpnew_pkg::status_t [NUM_FORMATS-1:0] fmt_special_status;
  logic [NUM_FORMATS-1:0]               fmt_result_is_special;
  for (genvar fmt = 0; fmt < int'(NUM_FORMATS); fmt++) begin : gen_special_results
    
    localparam int unsigned FP_WIDTH = fpnew_pkg::fp_width(fpnew_pkg::fp_format_e'(fmt));
    localparam int unsigned EXP_BITS = fpnew_pkg::exp_bits(fpnew_pkg::fp_format_e'(fmt));
    localparam int unsigned MAN_BITS = fpnew_pkg::man_bits(fpnew_pkg::fp_format_e'(fmt));
    localparam logic [EXP_BITS-1:0] QNAN_EXPONENT = '1;
    localparam logic [MAN_BITS-1:0] QNAN_MANTISSA = 2**(MAN_BITS-1);
    localparam logic [MAN_BITS-1:0] ZERO_MANTISSA = '0;
    if (FpFmtConfig[fmt]) begin : active_format
      always_comb begin : special_results
        logic [FP_WIDTH-1:0] special_res;
        
        special_res                = {1'b0, QNAN_EXPONENT, QNAN_MANTISSA}; 
        fmt_special_status[fmt]    = '0;
        fmt_result_is_special[fmt] = 1'b0;
        
        
        
        
        if ((info_a.is_inf && info_b.is_zero) || (info_a.is_zero && info_b.is_inf)) begin
          fmt_result_is_special[fmt] = 1'b1; 
          fmt_special_status[fmt].NV = 1'b1; 
        
        end else if (any_operand_nan) begin
          fmt_result_is_special[fmt] = 1'b1;           
          fmt_special_status[fmt].NV = signalling_nan; 
        
        end else if (any_operand_inf) begin
          fmt_result_is_special[fmt] = 1'b1; 
          
          if ((info_a.is_inf || info_b.is_inf) && info_c.is_inf && effective_subtraction)
            fmt_special_status[fmt].NV = 1'b1; 
          
          else if (info_a.is_inf || info_b.is_inf) begin
            
            special_res = {operand_a.sign ^ operand_b.sign, QNAN_EXPONENT, ZERO_MANTISSA};
          
          end else if (info_c.is_inf) begin
            
            special_res = {operand_c.sign, QNAN_EXPONENT, ZERO_MANTISSA};
          end
        end
        
        fmt_special_result[fmt]               = '1;
        fmt_special_result[fmt][FP_WIDTH-1:0] = special_res;
      end
    end else begin : inactive_format
      assign fmt_special_result[fmt] = '{default: fpnew_pkg::DONT_CARE};
    end
  end
  
  assign result_is_special = fmt_result_is_special[dst_fmt_q]; 
  
  assign special_status = fmt_special_status[dst_fmt_q];
  
  assign special_result = fmt_special_result[dst_fmt_q]; 
  
  
  
  logic signed [EXP_WIDTH-1:0] exponent_a, exponent_b, exponent_c;
  logic signed [EXP_WIDTH-1:0] exponent_addend, exponent_product, exponent_difference;
  logic signed [EXP_WIDTH-1:0] tentative_exponent;
  
  assign exponent_a = signed'({1'b0, operand_a.exponent});
  assign exponent_b = signed'({1'b0, operand_b.exponent});
  assign exponent_c = signed'({1'b0, operand_c.exponent});
  
  
  assign exponent_addend = signed'(exponent_c + $signed({1'b0, ~info_c.is_normal})); 
  
  assign exponent_product = (info_a.is_zero || info_b.is_zero) 
                            ? 2 - signed'(fpnew_pkg::bias(dst_fmt_q))
                            : signed'(exponent_a + info_a.is_subnormal
                                      + exponent_b + info_b.is_subnormal
                                      - 2*signed'(fpnew_pkg::bias(src_fmt_q))
                                      + signed'(fpnew_pkg::bias(dst_fmt_q))); 
  
  assign exponent_difference = exponent_addend - exponent_product;
  
  assign tentative_exponent = (exponent_difference > 0) ? exponent_addend : exponent_product;
  
  logic [SHIFT_AMOUNT_WIDTH-1:0] addend_shamt;
  always_comb begin : addend_shift_amount
    
    if (exponent_difference <= signed'(-2 * PRECISION_BITS - 1))
      addend_shamt = 3 * PRECISION_BITS + 4;
    
    else if (exponent_difference <= signed'(PRECISION_BITS + 2))
      addend_shamt = unsigned'(signed'(PRECISION_BITS) + 3 - exponent_difference);
    
    else
      addend_shamt = 0;
  end
  
  
  
  logic [PRECISION_BITS-1:0]   mantissa_a, mantissa_b, mantissa_c;
  logic [2*PRECISION_BITS-1:0] product;             
  logic [3*PRECISION_BITS+3:0] product_shifted;     
  
  assign mantissa_a = {info_a.is_normal, operand_a.mantissa};
  assign mantissa_b = {info_b.is_normal, operand_b.mantissa};
  assign mantissa_c = {info_c.is_normal, operand_c.mantissa};
  
  assign product = mantissa_a * mantissa_b;
  
  
  
  assign product_shifted = product << 2; 
  
  
  
  logic [3*PRECISION_BITS+3:0] addend_after_shift;  
  logic [PRECISION_BITS-1:0]   addend_sticky_bits;  
  logic                        sticky_before_add;   
  logic [3*PRECISION_BITS+3:0] addend_shifted;      
  logic                        inject_carry_in;     
  
  
  
  
  
  
  
  
  assign {addend_after_shift, addend_sticky_bits} =
      (mantissa_c << (3 * PRECISION_BITS + 4)) >> addend_shamt;
  assign sticky_before_add     = (| addend_sticky_bits);
  
  assign addend_shifted = (effective_subtraction) ? ~addend_after_shift : addend_after_shift;
  assign inject_carry_in = effective_subtraction & ~sticky_before_add;
  
  
  
  logic [3*PRECISION_BITS+4:0] sum_raw;   
  logic                        sum_carry; 
  logic [3*PRECISION_BITS+3:0] sum;       
  logic                        final_sign;
  
  assign sum_raw = product_shifted + addend_shifted + inject_carry_in;
  assign sum_carry = sum_raw[3*PRECISION_BITS+4];
  
  assign sum        = (effective_subtraction && ~sum_carry) ? -sum_raw : sum_raw;
  
  assign final_sign = (effective_subtraction && (sum_carry == tentative_sign))
                      ? 1'b1
                      : (effective_subtraction ? 1'b0 : tentative_sign);
  
  
  
  
  logic                          effective_subtraction_q;
  logic signed [EXP_WIDTH-1:0]   exponent_product_q;
  logic signed [EXP_WIDTH-1:0]   exponent_difference_q;
  logic signed [EXP_WIDTH-1:0]   tentative_exponent_q;
  logic [SHIFT_AMOUNT_WIDTH-1:0] addend_shamt_q;
  logic                          sticky_before_add_q;
  logic [3*PRECISION_BITS+3:0]   sum_q;
  logic                          final_sign_q;
  fpnew_pkg::fp_format_e         dst_fmt_q2;
  fpnew_pkg::roundmode_e         rnd_mode_q;
  logic                          result_is_special_q;
  fp_t                           special_result_q;
  fpnew_pkg::status_t            special_status_q;
  
  logic                  [0:NUM_MID_REGS]                         mid_pipe_eff_sub_q;
  logic signed           [0:NUM_MID_REGS][EXP_WIDTH-1:0]          mid_pipe_exp_prod_q;
  logic signed           [0:NUM_MID_REGS][EXP_WIDTH-1:0]          mid_pipe_exp_diff_q;
  logic signed           [0:NUM_MID_REGS][EXP_WIDTH-1:0]          mid_pipe_tent_exp_q;
  logic                  [0:NUM_MID_REGS][SHIFT_AMOUNT_WIDTH-1:0] mid_pipe_add_shamt_q;
  logic                  [0:NUM_MID_REGS]                         mid_pipe_sticky_q;
  logic                  [0:NUM_MID_REGS][3*PRECISION_BITS+3:0]   mid_pipe_sum_q;
  logic                  [0:NUM_MID_REGS]                         mid_pipe_final_sign_q;
  fpnew_pkg::roundmode_e [0:NUM_MID_REGS]                         mid_pipe_rnd_mode_q;
  fpnew_pkg::fp_format_e [0:NUM_MID_REGS]                         mid_pipe_dst_fmt_q;
  logic                  [0:NUM_MID_REGS]                         mid_pipe_res_is_spec_q;
  fp_t                   [0:NUM_MID_REGS]                         mid_pipe_spec_res_q;
  fpnew_pkg::status_t    [0:NUM_MID_REGS]                         mid_pipe_spec_stat_q;
  TagType                [0:NUM_MID_REGS]                         mid_pipe_tag_q;
  AuxType                [0:NUM_MID_REGS]                         mid_pipe_aux_q;
  logic                  [0:NUM_MID_REGS]                         mid_pipe_valid_q;
  
  logic [0:NUM_MID_REGS] mid_pipe_ready;
  
  assign mid_pipe_eff_sub_q[0]     = effective_subtraction;
  assign mid_pipe_exp_prod_q[0]    = exponent_product;
  assign mid_pipe_exp_diff_q[0]    = exponent_difference;
  assign mid_pipe_tent_exp_q[0]    = tentative_exponent;
  assign mid_pipe_add_shamt_q[0]   = addend_shamt;
  assign mid_pipe_sticky_q[0]      = sticky_before_add;
  assign mid_pipe_sum_q[0]         = sum;
  assign mid_pipe_final_sign_q[0]  = final_sign;
  assign mid_pipe_rnd_mode_q[0]    = inp_pipe_rnd_mode_q[NUM_INP_REGS];
  assign mid_pipe_dst_fmt_q[0]     = dst_fmt_q;
  assign mid_pipe_res_is_spec_q[0] = result_is_special;
  assign mid_pipe_spec_res_q[0]    = special_result;
  assign mid_pipe_spec_stat_q[0]   = special_status;
  assign mid_pipe_tag_q[0]         = inp_pipe_tag_q[NUM_INP_REGS];
  assign mid_pipe_aux_q[0]         = inp_pipe_aux_q[NUM_INP_REGS];
  assign mid_pipe_valid_q[0]       = inp_pipe_valid_q[NUM_INP_REGS];
  
  assign inp_pipe_ready[NUM_INP_REGS] = mid_pipe_ready[0];
  
  for (genvar i = 0; i < NUM_MID_REGS; i++) begin : gen_inside_pipeline
    
    logic reg_ena;
    
    
    
    assign mid_pipe_ready[i] = mid_pipe_ready[i+1] | ~mid_pipe_valid_q[i+1];
    
    
                           
                         
                            
  always_ff @(posedge (clk_i) or negedge (rst_ni)) begin                 
    if (!rst_ni) begin                                                   
      mid_pipe_valid_q[i+1] <= (1'b0);                                              
    end else begin                                                         
      mid_pipe_valid_q[i+1] <= (flush_i) ? (1'b0) : (mid_pipe_ready[i]) ? (mid_pipe_valid_q[i]) : (mid_pipe_valid_q[i+1]);       
    end                                                                    
  end
    
    assign reg_ena = mid_pipe_ready[i] & mid_pipe_valid_q[i];
    
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_eff_sub_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_eff_sub_q[i+1] <= (reg_ena) ? (mid_pipe_eff_sub_q[i]) : (mid_pipe_eff_sub_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_exp_prod_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_exp_prod_q[i+1] <= (reg_ena) ? (mid_pipe_exp_prod_q[i]) : (mid_pipe_exp_prod_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_exp_diff_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_exp_diff_q[i+1] <= (reg_ena) ? (mid_pipe_exp_diff_q[i]) : (mid_pipe_exp_diff_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_tent_exp_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_tent_exp_q[i+1] <= (reg_ena) ? (mid_pipe_tent_exp_q[i]) : (mid_pipe_tent_exp_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_add_shamt_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_add_shamt_q[i+1] <= (reg_ena) ? (mid_pipe_add_shamt_q[i]) : (mid_pipe_add_shamt_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_sticky_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_sticky_q[i+1] <= (reg_ena) ? (mid_pipe_sticky_q[i]) : (mid_pipe_sticky_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_sum_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_sum_q[i+1] <= (reg_ena) ? (mid_pipe_sum_q[i]) : (mid_pipe_sum_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_final_sign_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_final_sign_q[i+1] <= (reg_ena) ? (mid_pipe_final_sign_q[i]) : (mid_pipe_final_sign_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_rnd_mode_q[i+1] <= (fpnew_pkg::RNE);                        
    end else begin                                   
      mid_pipe_rnd_mode_q[i+1] <= (reg_ena) ? (mid_pipe_rnd_mode_q[i]) : (mid_pipe_rnd_mode_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_dst_fmt_q[i+1] <= (fpnew_pkg::fp_format_e'(0));                        
    end else begin                                   
      mid_pipe_dst_fmt_q[i+1] <= (reg_ena) ? (mid_pipe_dst_fmt_q[i]) : (mid_pipe_dst_fmt_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_res_is_spec_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_res_is_spec_q[i+1] <= (reg_ena) ? (mid_pipe_res_is_spec_q[i]) : (mid_pipe_res_is_spec_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_spec_res_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_spec_res_q[i+1] <= (reg_ena) ? (mid_pipe_spec_res_q[i]) : (mid_pipe_spec_res_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_spec_stat_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_spec_stat_q[i+1] <= (reg_ena) ? (mid_pipe_spec_stat_q[i]) : (mid_pipe_spec_stat_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_tag_q[i+1] <= (TagType'('0));                        
    end else begin                                   
      mid_pipe_tag_q[i+1] <= (reg_ena) ? (mid_pipe_tag_q[i]) : (mid_pipe_tag_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_aux_q[i+1] <= (AuxType'('0));                        
    end else begin                                   
      mid_pipe_aux_q[i+1] <= (reg_ena) ? (mid_pipe_aux_q[i]) : (mid_pipe_aux_q[i+1]);               
    end                                              
  end
  end
  
  assign effective_subtraction_q = mid_pipe_eff_sub_q[NUM_MID_REGS];
  assign exponent_product_q      = mid_pipe_exp_prod_q[NUM_MID_REGS];
  assign exponent_difference_q   = mid_pipe_exp_diff_q[NUM_MID_REGS];
  assign tentative_exponent_q    = mid_pipe_tent_exp_q[NUM_MID_REGS];
  assign addend_shamt_q          = mid_pipe_add_shamt_q[NUM_MID_REGS];
  assign sticky_before_add_q     = mid_pipe_sticky_q[NUM_MID_REGS];
  assign sum_q                   = mid_pipe_sum_q[NUM_MID_REGS];
  assign final_sign_q            = mid_pipe_final_sign_q[NUM_MID_REGS];
  assign rnd_mode_q              = mid_pipe_rnd_mode_q[NUM_MID_REGS];
  assign dst_fmt_q2              = mid_pipe_dst_fmt_q[NUM_MID_REGS];
  assign result_is_special_q     = mid_pipe_res_is_spec_q[NUM_MID_REGS];
  assign special_result_q        = mid_pipe_spec_res_q[NUM_MID_REGS];
  assign special_status_q        = mid_pipe_spec_stat_q[NUM_MID_REGS];
  
  
  
  logic        [LOWER_SUM_WIDTH-1:0]  sum_lower;              
  logic        [LZC_RESULT_WIDTH-1:0] leading_zero_count;     
  logic signed [LZC_RESULT_WIDTH:0]   leading_zero_count_sgn; 
  logic                               lzc_zeroes;             
  logic        [SHIFT_AMOUNT_WIDTH-1:0] norm_shamt; 
  logic signed [EXP_WIDTH-1:0]          normalized_exponent;
  logic [3*PRECISION_BITS+4:0] sum_shifted;       
  logic [PRECISION_BITS:0]     final_mantissa;    
  logic [2*PRECISION_BITS+2:0] sum_sticky_bits;   
  logic                        sticky_after_norm; 
  logic signed [EXP_WIDTH-1:0] final_exponent;
  assign sum_lower = sum_q[LOWER_SUM_WIDTH-1:0];
  
  lzc #(
    .WIDTH ( LOWER_SUM_WIDTH ),
    .MODE  ( 1               ) 
  ) i_lzc (
    .in_i    ( sum_lower          ),
    .cnt_o   ( leading_zero_count ),
    .empty_o ( lzc_zeroes         )
  );
  assign leading_zero_count_sgn = signed'({1'b0, leading_zero_count});
  
  always_comb begin : norm_shift_amount
    
    if ((exponent_difference_q <= 0) || (effective_subtraction_q && (exponent_difference_q <= 2))) begin
      
      if ((exponent_product_q - leading_zero_count_sgn + 1 >= 0) && !lzc_zeroes) begin
        
        norm_shamt          = PRECISION_BITS + 2 + leading_zero_count;
        normalized_exponent = exponent_product_q - leading_zero_count_sgn + 1; 
      
      end else begin
        
        norm_shamt          = unsigned'(signed'(PRECISION_BITS + 2 + exponent_product_q));
        normalized_exponent = 0; 
      end
    
    end else begin
      norm_shamt          = addend_shamt_q; 
      normalized_exponent = tentative_exponent_q;
    end
  end
  
  assign sum_shifted       = sum_q << norm_shamt;
  
  
  always_comb begin : small_norm
    
    {final_mantissa, sum_sticky_bits} = sum_shifted;
    final_exponent                    = normalized_exponent;
    
    if (sum_shifted[3*PRECISION_BITS+4]) begin 
      {final_mantissa, sum_sticky_bits} = sum_shifted >> 1;
      final_exponent                    = normalized_exponent + 1;
    
    end else if (sum_shifted[3*PRECISION_BITS+3]) begin 
      
    
    end else if (normalized_exponent > 1) begin
      {final_mantissa, sum_sticky_bits} = sum_shifted << 1;
      final_exponent                    = normalized_exponent - 1;
    
    end else begin
      final_exponent = '0;
    end
  end
  
  assign sticky_after_norm = (| {sum_sticky_bits}) | sticky_before_add_q;
  
  
  
  logic                                     pre_round_sign;
  logic [SUPER_EXP_BITS+SUPER_MAN_BITS-1:0] pre_round_abs; 
  logic [1:0]                               round_sticky_bits;
  logic of_before_round, of_after_round; 
  logic uf_before_round, uf_after_round; 
  logic [NUM_FORMATS-1:0][SUPER_EXP_BITS+SUPER_MAN_BITS-1:0] fmt_pre_round_abs; 
  logic [NUM_FORMATS-1:0][1:0]                               fmt_round_sticky_bits;
  logic [NUM_FORMATS-1:0]                                    fmt_of_after_round;
  logic [NUM_FORMATS-1:0]                                    fmt_uf_after_round;
  logic                                     rounded_sign;
  logic [SUPER_EXP_BITS+SUPER_MAN_BITS-1:0] rounded_abs; 
  logic                                     result_zero;
  
  assign of_before_round = final_exponent >= 2**(fpnew_pkg::exp_bits(dst_fmt_q2))-1; 
  assign uf_before_round = final_exponent == 0;               
  
  for (genvar fmt = 0; fmt < int'(NUM_FORMATS); fmt++) begin : gen_res_assemble
    
    localparam int unsigned EXP_BITS = fpnew_pkg::exp_bits(fpnew_pkg::fp_format_e'(fmt));
    localparam int unsigned MAN_BITS = fpnew_pkg::man_bits(fpnew_pkg::fp_format_e'(fmt));
    logic [EXP_BITS-1:0] pre_round_exponent;
    logic [MAN_BITS-1:0] pre_round_mantissa;
    if (FpFmtConfig[fmt]) begin : active_format
      assign pre_round_exponent = (of_before_round) ? 2**EXP_BITS-2 : final_exponent[EXP_BITS-1:0];
      assign pre_round_mantissa = (of_before_round) ? '1 : final_mantissa[SUPER_MAN_BITS-:MAN_BITS];
      
      assign fmt_pre_round_abs[fmt] = {pre_round_exponent, pre_round_mantissa}; 
      
      assign fmt_round_sticky_bits[fmt][1] = final_mantissa[SUPER_MAN_BITS-MAN_BITS] |
                                             of_before_round;
      
      if (MAN_BITS < SUPER_MAN_BITS) begin : narrow_sticky
        assign fmt_round_sticky_bits[fmt][0] = (| final_mantissa[SUPER_MAN_BITS-MAN_BITS-1:0]) |
                                               sticky_after_norm | of_before_round;
      end else begin : normal_sticky
        assign fmt_round_sticky_bits[fmt][0] = sticky_after_norm | of_before_round;
      end
    end else begin : inactive_format
      assign fmt_pre_round_abs[fmt] = '{default: fpnew_pkg::DONT_CARE};
      assign fmt_round_sticky_bits[fmt] = '{default: fpnew_pkg::DONT_CARE};
    end
  end
  
  assign pre_round_sign     = final_sign_q;
  assign pre_round_abs      = fmt_pre_round_abs[dst_fmt_q2];
  
  assign round_sticky_bits  = fmt_round_sticky_bits[dst_fmt_q2];
  
  fpnew_rounding #(
    .AbsWidth ( SUPER_EXP_BITS + SUPER_MAN_BITS )
  ) i_fpnew_rounding (
    .abs_value_i             ( pre_round_abs           ),
    .sign_i                  ( pre_round_sign          ),
    .round_sticky_bits_i     ( round_sticky_bits       ),
    .rnd_mode_i              ( rnd_mode_q              ),
    .effective_subtraction_i ( effective_subtraction_q ),
    .abs_rounded_o           ( rounded_abs             ),
    .sign_o                  ( rounded_sign            ),
    .exact_zero_o            ( result_zero             )
  );
  logic [NUM_FORMATS-1:0][WIDTH-1:0] fmt_result;
  for (genvar fmt = 0; fmt < int'(NUM_FORMATS); fmt++) begin : gen_sign_inject
    
    localparam int unsigned FP_WIDTH = fpnew_pkg::fp_width(fpnew_pkg::fp_format_e'(fmt));
    localparam int unsigned EXP_BITS = fpnew_pkg::exp_bits(fpnew_pkg::fp_format_e'(fmt));
    localparam int unsigned MAN_BITS = fpnew_pkg::man_bits(fpnew_pkg::fp_format_e'(fmt));
    if (FpFmtConfig[fmt]) begin : active_format
      always_comb begin : post_process
        
        fmt_uf_after_round[fmt] = rounded_abs[EXP_BITS+MAN_BITS-1:MAN_BITS] == '0; 
        fmt_of_after_round[fmt] = rounded_abs[EXP_BITS+MAN_BITS-1:MAN_BITS] == '1; 
        
        fmt_result[fmt]               = '1;
        fmt_result[fmt][FP_WIDTH-1:0] = {rounded_sign, rounded_abs[EXP_BITS+MAN_BITS-1:0]};
      end
    end else begin : inactive_format
      assign fmt_uf_after_round[fmt] = fpnew_pkg::DONT_CARE;
      assign fmt_of_after_round[fmt] = fpnew_pkg::DONT_CARE;
      assign fmt_result[fmt]         = '{default: fpnew_pkg::DONT_CARE};
    end
  end
  
  assign uf_after_round = fmt_uf_after_round[dst_fmt_q2];
  assign of_after_round = fmt_of_after_round[dst_fmt_q2];
  
  
  
  logic [WIDTH-1:0]     regular_result;
  fpnew_pkg::status_t   regular_status;
  
  assign regular_result = fmt_result[dst_fmt_q2];
  assign regular_status.NV = 1'b0; 
  assign regular_status.DZ = 1'b0; 
  assign regular_status.OF = of_before_round | of_after_round;   
  assign regular_status.UF = uf_after_round & regular_status.NX; 
  assign regular_status.NX = (| round_sticky_bits) | of_before_round | of_after_round;
  
  logic [WIDTH-1:0]   result_d;
  fpnew_pkg::status_t status_d;
  
  assign result_d = result_is_special_q ? special_result_q : regular_result;
  assign status_d = result_is_special_q ? special_status_q : regular_status;
  
  
  
  
  logic               [0:NUM_OUT_REGS][WIDTH-1:0] out_pipe_result_q;
  fpnew_pkg::status_t [0:NUM_OUT_REGS]            out_pipe_status_q;
  TagType             [0:NUM_OUT_REGS]            out_pipe_tag_q;
  AuxType             [0:NUM_OUT_REGS]            out_pipe_aux_q;
  logic               [0:NUM_OUT_REGS]            out_pipe_valid_q;
  
  logic [0:NUM_OUT_REGS] out_pipe_ready;
  
  assign out_pipe_result_q[0] = result_d;
  assign out_pipe_status_q[0] = status_d;
  assign out_pipe_tag_q[0]    = mid_pipe_tag_q[NUM_MID_REGS];
  assign out_pipe_aux_q[0]    = mid_pipe_aux_q[NUM_MID_REGS];
  assign out_pipe_valid_q[0]  = mid_pipe_valid_q[NUM_MID_REGS];
  
  assign mid_pipe_ready[NUM_MID_REGS] = out_pipe_ready[0];
  
  for (genvar i = 0; i < NUM_OUT_REGS; i++) begin : gen_output_pipeline
    
    logic reg_ena;
    
    
    
    assign out_pipe_ready[i] = out_pipe_ready[i+1] | ~out_pipe_valid_q[i+1];
    
    
                           
                         
                            
  always_ff @(posedge (clk_i) or negedge (rst_ni)) begin                 
    if (!rst_ni) begin                                                   
      out_pipe_valid_q[i+1] <= (1'b0);                                              
    end else begin                                                         
      out_pipe_valid_q[i+1] <= (flush_i) ? (1'b0) : (out_pipe_ready[i]) ? (out_pipe_valid_q[i]) : (out_pipe_valid_q[i+1]);       
    end                                                                    
  end
    
    assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
    
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_result_q[i+1] <= ('0);                        
    end else begin                                   
      out_pipe_result_q[i+1] <= (reg_ena) ? (out_pipe_result_q[i]) : (out_pipe_result_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_status_q[i+1] <= ('0);                        
    end else begin                                   
      out_pipe_status_q[i+1] <= (reg_ena) ? (out_pipe_status_q[i]) : (out_pipe_status_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_tag_q[i+1] <= (TagType'('0));                        
    end else begin                                   
      out_pipe_tag_q[i+1] <= (reg_ena) ? (out_pipe_tag_q[i]) : (out_pipe_tag_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_aux_q[i+1] <= (AuxType'('0));                        
    end else begin                                   
      out_pipe_aux_q[i+1] <= (reg_ena) ? (out_pipe_aux_q[i]) : (out_pipe_aux_q[i+1]);               
    end                                              
  end
  end
  
  assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
  
  assign result_o        = out_pipe_result_q[NUM_OUT_REGS];
  assign status_o        = out_pipe_status_q[NUM_OUT_REGS];
  assign extension_bit_o = 1'b1; 
  assign tag_o           = out_pipe_tag_q[NUM_OUT_REGS];
  assign aux_o           = out_pipe_aux_q[NUM_OUT_REGS];
  assign out_valid_o     = out_pipe_valid_q[NUM_OUT_REGS];
  assign busy_o          = (| {inp_pipe_valid_q, mid_pipe_valid_q, out_pipe_valid_q});
endmodule
                                      
module fpnew_fma #(
  parameter fpnew_pkg::fp_format_e   FpFormat    = fpnew_pkg::fp_format_e'(0),
  parameter int unsigned             NumPipeRegs = 0,
  parameter fpnew_pkg::pipe_config_t PipeConfig  = fpnew_pkg::BEFORE,
  parameter type                     TagType     = logic,
  parameter type                     AuxType     = logic,
  localparam int unsigned WIDTH = fpnew_pkg::fp_width(FpFormat) 
) (
  input logic                      clk_i,
  input logic                      rst_ni,
  
  input logic [2:0][WIDTH-1:0]     operands_i, 
  input logic [2:0]                is_boxed_i, 
  input fpnew_pkg::roundmode_e     rnd_mode_i,
  input fpnew_pkg::operation_e     op_i,
  input logic                      op_mod_i,
  input TagType                    tag_i,
  input AuxType                    aux_i,
  
  input  logic                     in_valid_i,
  output logic                     in_ready_o,
  input  logic                     flush_i,
  
  output logic [WIDTH-1:0]         result_o,
  output fpnew_pkg::status_t       status_o,
  output logic                     extension_bit_o,
  output TagType                   tag_o,
  output AuxType                   aux_o,
  
  output logic                     out_valid_o,
  input  logic                     out_ready_i,
  
  output logic                     busy_o
);
  
  
  
  localparam int unsigned EXP_BITS = fpnew_pkg::exp_bits(FpFormat);
  localparam int unsigned MAN_BITS = fpnew_pkg::man_bits(FpFormat);
  localparam int unsigned BIAS     = fpnew_pkg::bias(FpFormat);
  
  localparam int unsigned PRECISION_BITS = MAN_BITS + 1;
  
  localparam int unsigned LOWER_SUM_WIDTH  = 2 * PRECISION_BITS + 3;
  localparam int unsigned LZC_RESULT_WIDTH = $clog2(LOWER_SUM_WIDTH);
  
  
  
  localparam int unsigned EXP_WIDTH = unsigned'(fpnew_pkg::maximum(EXP_BITS + 2, LZC_RESULT_WIDTH));
  
  localparam int unsigned SHIFT_AMOUNT_WIDTH = $clog2(3 * PRECISION_BITS + 3);
  
  localparam NUM_INP_REGS = PipeConfig == fpnew_pkg::BEFORE
                            ? NumPipeRegs
                            : (PipeConfig == fpnew_pkg::DISTRIBUTED
                               ? ((NumPipeRegs + 1) / 3) 
                               : 0); 
  localparam NUM_MID_REGS = PipeConfig == fpnew_pkg::INSIDE
                          ? NumPipeRegs
                          : (PipeConfig == fpnew_pkg::DISTRIBUTED
                             ? ((NumPipeRegs + 2) / 3) 
                             : 0); 
  localparam NUM_OUT_REGS = PipeConfig == fpnew_pkg::AFTER
                            ? NumPipeRegs
                            : (PipeConfig == fpnew_pkg::DISTRIBUTED
                               ? (NumPipeRegs / 3) 
                               : 0); 
  
  
  
  typedef struct packed {
    logic                sign;
    logic [EXP_BITS-1:0] exponent;
    logic [MAN_BITS-1:0] mantissa;
  } fp_t;
  
  
  
  
  logic                  [0:NUM_INP_REGS][2:0][WIDTH-1:0] inp_pipe_operands_q;
  logic                  [0:NUM_INP_REGS][2:0]            inp_pipe_is_boxed_q;
  fpnew_pkg::roundmode_e [0:NUM_INP_REGS]                 inp_pipe_rnd_mode_q;
  fpnew_pkg::operation_e [0:NUM_INP_REGS]                 inp_pipe_op_q;
  logic                  [0:NUM_INP_REGS]                 inp_pipe_op_mod_q;
  TagType                [0:NUM_INP_REGS]                 inp_pipe_tag_q;
  AuxType                [0:NUM_INP_REGS]                 inp_pipe_aux_q;
  logic                  [0:NUM_INP_REGS]                 inp_pipe_valid_q;
  
  logic [0:NUM_INP_REGS] inp_pipe_ready;
  
  assign inp_pipe_operands_q[0] = operands_i;
  assign inp_pipe_is_boxed_q[0] = is_boxed_i;
  assign inp_pipe_rnd_mode_q[0] = rnd_mode_i;
  assign inp_pipe_op_q[0]       = op_i;
  assign inp_pipe_op_mod_q[0]   = op_mod_i;
  assign inp_pipe_tag_q[0]      = tag_i;
  assign inp_pipe_aux_q[0]      = aux_i;
  assign inp_pipe_valid_q[0]    = in_valid_i;
  
  assign in_ready_o = inp_pipe_ready[0];
  
  for (genvar i = 0; i < NUM_INP_REGS; i++) begin : gen_input_pipeline
    
    logic reg_ena;
    
    
    
    assign inp_pipe_ready[i] = inp_pipe_ready[i+1] | ~inp_pipe_valid_q[i+1];
    
    
                           
                         
                            
  always_ff @(posedge (clk_i) or negedge (rst_ni)) begin                 
    if (!rst_ni) begin                                                   
      inp_pipe_valid_q[i+1] <= (1'b0);                                              
    end else begin                                                         
      inp_pipe_valid_q[i+1] <= (flush_i) ? (1'b0) : (inp_pipe_ready[i]) ? (inp_pipe_valid_q[i]) : (inp_pipe_valid_q[i+1]);       
    end                                                                    
  end
    
    assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
    
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_operands_q[i+1] <= ('0);                        
    end else begin                                   
      inp_pipe_operands_q[i+1] <= (reg_ena) ? (inp_pipe_operands_q[i]) : (inp_pipe_operands_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_is_boxed_q[i+1] <= ('0);                        
    end else begin                                   
      inp_pipe_is_boxed_q[i+1] <= (reg_ena) ? (inp_pipe_is_boxed_q[i]) : (inp_pipe_is_boxed_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_rnd_mode_q[i+1] <= (fpnew_pkg::RNE);                        
    end else begin                                   
      inp_pipe_rnd_mode_q[i+1] <= (reg_ena) ? (inp_pipe_rnd_mode_q[i]) : (inp_pipe_rnd_mode_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_op_q[i+1] <= (fpnew_pkg::FMADD);                        
    end else begin                                   
      inp_pipe_op_q[i+1] <= (reg_ena) ? (inp_pipe_op_q[i]) : (inp_pipe_op_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_op_mod_q[i+1] <= ('0);                        
    end else begin                                   
      inp_pipe_op_mod_q[i+1] <= (reg_ena) ? (inp_pipe_op_mod_q[i]) : (inp_pipe_op_mod_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_tag_q[i+1] <= (TagType'('0));                        
    end else begin                                   
      inp_pipe_tag_q[i+1] <= (reg_ena) ? (inp_pipe_tag_q[i]) : (inp_pipe_tag_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_aux_q[i+1] <= (AuxType'('0));                        
    end else begin                                   
      inp_pipe_aux_q[i+1] <= (reg_ena) ? (inp_pipe_aux_q[i]) : (inp_pipe_aux_q[i+1]);               
    end                                              
  end
  end
  
  
  
  fpnew_pkg::fp_info_t [2:0] info_q;
  
  fpnew_classifier #(
    .FpFormat    ( FpFormat ),
    .NumOperands ( 3        )
    ) i_class_inputs (
    .operands_i ( inp_pipe_operands_q[NUM_INP_REGS] ),
    .is_boxed_i ( inp_pipe_is_boxed_q[NUM_INP_REGS] ),
    .info_o     ( info_q                            )
  );
  fp_t                 operand_a, operand_b, operand_c;
  fpnew_pkg::fp_info_t info_a,    info_b,    info_c;
  
  
  
  
  
  
  
  
  
  
  
  
  always_comb begin : op_select
    
    operand_a = inp_pipe_operands_q[NUM_INP_REGS][0];
    operand_b = inp_pipe_operands_q[NUM_INP_REGS][1];
    operand_c = inp_pipe_operands_q[NUM_INP_REGS][2];
    info_a    = info_q[0];
    info_b    = info_q[1];
    info_c    = info_q[2];
    
    operand_c.sign = operand_c.sign ^ inp_pipe_op_mod_q[NUM_INP_REGS];
    unique case (inp_pipe_op_q[NUM_INP_REGS])
      fpnew_pkg::FMADD:  ; 
      fpnew_pkg::FNMSUB: operand_a.sign = ~operand_a.sign; 
      fpnew_pkg::ADD: begin 
        operand_a = '{sign: 1'b0, exponent: BIAS, mantissa: '0};
        info_a    = '{is_normal: 1'b1, is_boxed: 1'b1, default: 1'b0}; 
      end
      fpnew_pkg::MUL: begin 
        operand_c = '{sign: 1'b1, exponent: '0, mantissa: '0};
        info_c    = '{is_zero: 1'b1, is_boxed: 1'b1, default: 1'b0}; 
      end
      default: begin 
        operand_a  = '{default: fpnew_pkg::DONT_CARE};
        operand_b  = '{default: fpnew_pkg::DONT_CARE};
        operand_c  = '{default: fpnew_pkg::DONT_CARE};
        info_a     = '{default: fpnew_pkg::DONT_CARE};
        info_b     = '{default: fpnew_pkg::DONT_CARE};
        info_c     = '{default: fpnew_pkg::DONT_CARE};
      end
    endcase
  end
  
  
  
  logic any_operand_inf;
  logic any_operand_nan;
  logic signalling_nan;
  logic effective_subtraction;
  logic tentative_sign;
  
  assign any_operand_inf = (| {info_a.is_inf,        info_b.is_inf,        info_c.is_inf});
  assign any_operand_nan = (| {info_a.is_nan,        info_b.is_nan,        info_c.is_nan});
  assign signalling_nan  = (| {info_a.is_signalling, info_b.is_signalling, info_c.is_signalling});
  
  assign effective_subtraction = operand_a.sign ^ operand_b.sign ^ operand_c.sign;
  
  assign tentative_sign = operand_a.sign ^ operand_b.sign;
  
  
  
  fp_t                special_result;
  fpnew_pkg::status_t special_status;
  logic               result_is_special;
  always_comb begin : special_cases
    
    special_result    = '{sign: 1'b0, exponent: '1, mantissa: 2**(MAN_BITS-1)}; 
    special_status    = '0;
    result_is_special = 1'b0;
    
    
    
    
    if ((info_a.is_inf && info_b.is_zero) || (info_a.is_zero && info_b.is_inf)) begin
      result_is_special = 1'b1; 
      special_status.NV = 1'b1; 
    
    end else if (any_operand_nan) begin
      result_is_special = 1'b1;           
      special_status.NV = signalling_nan; 
    
    end else if (any_operand_inf) begin
      result_is_special = 1'b1; 
      
      if ((info_a.is_inf || info_b.is_inf) && info_c.is_inf && effective_subtraction)
        special_status.NV = 1'b1; 
      
      else if (info_a.is_inf || info_b.is_inf) begin
        
        special_result    = '{sign: operand_a.sign ^ operand_b.sign, exponent: '1, mantissa: '0};
      
      end else if (info_c.is_inf) begin
        
        special_result    = '{sign: operand_c.sign, exponent: '1, mantissa: '0};
      end
    end
  end
  
  
  
  logic signed [EXP_WIDTH-1:0] exponent_a, exponent_b, exponent_c;
  logic signed [EXP_WIDTH-1:0] exponent_addend, exponent_product, exponent_difference;
  logic signed [EXP_WIDTH-1:0] tentative_exponent;
  
  assign exponent_a = signed'({1'b0, operand_a.exponent});
  assign exponent_b = signed'({1'b0, operand_b.exponent});
  assign exponent_c = signed'({1'b0, operand_c.exponent});
  
  
  assign exponent_addend = signed'(exponent_c + $signed({1'b0, ~info_c.is_normal})); 
  
  assign exponent_product = (info_a.is_zero || info_b.is_zero)
                            ? 2 - signed'(BIAS) 
                            : signed'(exponent_a + info_a.is_subnormal
                                      + exponent_b + info_b.is_subnormal
                                      - signed'(BIAS));
  
  assign exponent_difference = exponent_addend - exponent_product;
  
  assign tentative_exponent = (exponent_difference > 0) ? exponent_addend : exponent_product;
  
  logic [SHIFT_AMOUNT_WIDTH-1:0] addend_shamt;
  always_comb begin : addend_shift_amount
    
    if (exponent_difference <= signed'(-2 * PRECISION_BITS - 1))
      addend_shamt = 3 * PRECISION_BITS + 4;
    
    else if (exponent_difference <= signed'(PRECISION_BITS + 2))
      addend_shamt = unsigned'(signed'(PRECISION_BITS) + 3 - exponent_difference);
    
    else
      addend_shamt = 0;
  end
  
  
  
  logic [PRECISION_BITS-1:0]   mantissa_a, mantissa_b, mantissa_c;
  logic [2*PRECISION_BITS-1:0] product;             
  logic [3*PRECISION_BITS+3:0] product_shifted;     
  
  assign mantissa_a = {info_a.is_normal, operand_a.mantissa};
  assign mantissa_b = {info_b.is_normal, operand_b.mantissa};
  assign mantissa_c = {info_c.is_normal, operand_c.mantissa};
  
  assign product = mantissa_a * mantissa_b;
  
  
  
  assign product_shifted = product << 2; 
  
  
  
  logic [3*PRECISION_BITS+3:0] addend_after_shift;  
  logic [PRECISION_BITS-1:0]   addend_sticky_bits;  
  logic                        sticky_before_add;   
  logic [3*PRECISION_BITS+3:0] addend_shifted;      
  logic                        inject_carry_in;     
  
  
  
  
  
  
  
  
  assign {addend_after_shift, addend_sticky_bits} =
      (mantissa_c << (3 * PRECISION_BITS + 4)) >> addend_shamt;
  assign sticky_before_add     = (| addend_sticky_bits);
  
  
  assign addend_shifted  = (effective_subtraction) ? ~addend_after_shift : addend_after_shift;
  assign inject_carry_in = effective_subtraction & ~sticky_before_add;
  
  
  
  logic [3*PRECISION_BITS+4:0] sum_raw;   
  logic                        sum_carry; 
  logic [3*PRECISION_BITS+3:0] sum;       
  logic                        final_sign;
  
  assign sum_raw = product_shifted + addend_shifted + inject_carry_in;
  assign sum_carry = sum_raw[3*PRECISION_BITS+4];
  
  assign sum        = (effective_subtraction && ~sum_carry) ? -sum_raw : sum_raw;
  
  assign final_sign = (effective_subtraction && (sum_carry == tentative_sign))
                      ? 1'b1
                      : (effective_subtraction ? 1'b0 : tentative_sign);
  
  
  
  
  logic                          effective_subtraction_q;
  logic signed [EXP_WIDTH-1:0]   exponent_product_q;
  logic signed [EXP_WIDTH-1:0]   exponent_difference_q;
  logic signed [EXP_WIDTH-1:0]   tentative_exponent_q;
  logic [SHIFT_AMOUNT_WIDTH-1:0] addend_shamt_q;
  logic                          sticky_before_add_q;
  logic [3*PRECISION_BITS+3:0]   sum_q;
  logic                          final_sign_q;
  fpnew_pkg::roundmode_e         rnd_mode_q;
  logic                          result_is_special_q;
  fp_t                           special_result_q;
  fpnew_pkg::status_t            special_status_q;
  
  logic                  [0:NUM_MID_REGS]                         mid_pipe_eff_sub_q;
  logic signed           [0:NUM_MID_REGS][EXP_WIDTH-1:0]          mid_pipe_exp_prod_q;
  logic signed           [0:NUM_MID_REGS][EXP_WIDTH-1:0]          mid_pipe_exp_diff_q;
  logic signed           [0:NUM_MID_REGS][EXP_WIDTH-1:0]          mid_pipe_tent_exp_q;
  logic                  [0:NUM_MID_REGS][SHIFT_AMOUNT_WIDTH-1:0] mid_pipe_add_shamt_q;
  logic                  [0:NUM_MID_REGS]                         mid_pipe_sticky_q;
  logic                  [0:NUM_MID_REGS][3*PRECISION_BITS+3:0]   mid_pipe_sum_q;
  logic                  [0:NUM_MID_REGS]                         mid_pipe_final_sign_q;
  fpnew_pkg::roundmode_e [0:NUM_MID_REGS]                         mid_pipe_rnd_mode_q;
  logic                  [0:NUM_MID_REGS]                         mid_pipe_res_is_spec_q;
  fp_t                   [0:NUM_MID_REGS]                         mid_pipe_spec_res_q;
  fpnew_pkg::status_t    [0:NUM_MID_REGS]                         mid_pipe_spec_stat_q;
  TagType                [0:NUM_MID_REGS]                         mid_pipe_tag_q;
  AuxType                [0:NUM_MID_REGS]                         mid_pipe_aux_q;
  logic                  [0:NUM_MID_REGS]                         mid_pipe_valid_q;
  
  logic [0:NUM_MID_REGS] mid_pipe_ready;
  
  assign mid_pipe_eff_sub_q[0]     = effective_subtraction;
  assign mid_pipe_exp_prod_q[0]    = exponent_product;
  assign mid_pipe_exp_diff_q[0]    = exponent_difference;
  assign mid_pipe_tent_exp_q[0]    = tentative_exponent;
  assign mid_pipe_add_shamt_q[0]   = addend_shamt;
  assign mid_pipe_sticky_q[0]      = sticky_before_add;
  assign mid_pipe_sum_q[0]         = sum;
  assign mid_pipe_final_sign_q[0]  = final_sign;
  assign mid_pipe_rnd_mode_q[0]    = inp_pipe_rnd_mode_q[NUM_INP_REGS];
  assign mid_pipe_res_is_spec_q[0] = result_is_special;
  assign mid_pipe_spec_res_q[0]    = special_result;
  assign mid_pipe_spec_stat_q[0]   = special_status;
  assign mid_pipe_tag_q[0]         = inp_pipe_tag_q[NUM_INP_REGS];
  assign mid_pipe_aux_q[0]         = inp_pipe_aux_q[NUM_INP_REGS];
  assign mid_pipe_valid_q[0]       = inp_pipe_valid_q[NUM_INP_REGS];
  
  assign inp_pipe_ready[NUM_INP_REGS] = mid_pipe_ready[0];
  
  for (genvar i = 0; i < NUM_MID_REGS; i++) begin : gen_inside_pipeline
    
    logic reg_ena;
    
    
    
    assign mid_pipe_ready[i] = mid_pipe_ready[i+1] | ~mid_pipe_valid_q[i+1];
    
    
                           
                         
                            
  always_ff @(posedge (clk_i) or negedge (rst_ni)) begin                 
    if (!rst_ni) begin                                                   
      mid_pipe_valid_q[i+1] <= (1'b0);                                              
    end else begin                                                         
      mid_pipe_valid_q[i+1] <= (flush_i) ? (1'b0) : (mid_pipe_ready[i]) ? (mid_pipe_valid_q[i]) : (mid_pipe_valid_q[i+1]);       
    end                                                                    
  end
    
    assign reg_ena = mid_pipe_ready[i] & mid_pipe_valid_q[i];
    
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_eff_sub_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_eff_sub_q[i+1] <= (reg_ena) ? (mid_pipe_eff_sub_q[i]) : (mid_pipe_eff_sub_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_exp_prod_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_exp_prod_q[i+1] <= (reg_ena) ? (mid_pipe_exp_prod_q[i]) : (mid_pipe_exp_prod_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_exp_diff_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_exp_diff_q[i+1] <= (reg_ena) ? (mid_pipe_exp_diff_q[i]) : (mid_pipe_exp_diff_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_tent_exp_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_tent_exp_q[i+1] <= (reg_ena) ? (mid_pipe_tent_exp_q[i]) : (mid_pipe_tent_exp_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_add_shamt_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_add_shamt_q[i+1] <= (reg_ena) ? (mid_pipe_add_shamt_q[i]) : (mid_pipe_add_shamt_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_sticky_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_sticky_q[i+1] <= (reg_ena) ? (mid_pipe_sticky_q[i]) : (mid_pipe_sticky_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_sum_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_sum_q[i+1] <= (reg_ena) ? (mid_pipe_sum_q[i]) : (mid_pipe_sum_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_final_sign_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_final_sign_q[i+1] <= (reg_ena) ? (mid_pipe_final_sign_q[i]) : (mid_pipe_final_sign_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_rnd_mode_q[i+1] <= (fpnew_pkg::RNE);                        
    end else begin                                   
      mid_pipe_rnd_mode_q[i+1] <= (reg_ena) ? (mid_pipe_rnd_mode_q[i]) : (mid_pipe_rnd_mode_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_res_is_spec_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_res_is_spec_q[i+1] <= (reg_ena) ? (mid_pipe_res_is_spec_q[i]) : (mid_pipe_res_is_spec_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_spec_res_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_spec_res_q[i+1] <= (reg_ena) ? (mid_pipe_spec_res_q[i]) : (mid_pipe_spec_res_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_spec_stat_q[i+1] <= ('0);                        
    end else begin                                   
      mid_pipe_spec_stat_q[i+1] <= (reg_ena) ? (mid_pipe_spec_stat_q[i]) : (mid_pipe_spec_stat_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_tag_q[i+1] <= (TagType'('0));                        
    end else begin                                   
      mid_pipe_tag_q[i+1] <= (reg_ena) ? (mid_pipe_tag_q[i]) : (mid_pipe_tag_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      mid_pipe_aux_q[i+1] <= (AuxType'('0));                        
    end else begin                                   
      mid_pipe_aux_q[i+1] <= (reg_ena) ? (mid_pipe_aux_q[i]) : (mid_pipe_aux_q[i+1]);               
    end                                              
  end
  end
  
  assign effective_subtraction_q = mid_pipe_eff_sub_q[NUM_MID_REGS];
  assign exponent_product_q      = mid_pipe_exp_prod_q[NUM_MID_REGS];
  assign exponent_difference_q   = mid_pipe_exp_diff_q[NUM_MID_REGS];
  assign tentative_exponent_q    = mid_pipe_tent_exp_q[NUM_MID_REGS];
  assign addend_shamt_q          = mid_pipe_add_shamt_q[NUM_MID_REGS];
  assign sticky_before_add_q     = mid_pipe_sticky_q[NUM_MID_REGS];
  assign sum_q                   = mid_pipe_sum_q[NUM_MID_REGS];
  assign final_sign_q            = mid_pipe_final_sign_q[NUM_MID_REGS];
  assign rnd_mode_q              = mid_pipe_rnd_mode_q[NUM_MID_REGS];
  assign result_is_special_q     = mid_pipe_res_is_spec_q[NUM_MID_REGS];
  assign special_result_q        = mid_pipe_spec_res_q[NUM_MID_REGS];
  assign special_status_q        = mid_pipe_spec_stat_q[NUM_MID_REGS];
  
  
  
  logic        [LOWER_SUM_WIDTH-1:0]  sum_lower;              
  logic        [LZC_RESULT_WIDTH-1:0] leading_zero_count;     
  logic signed [LZC_RESULT_WIDTH:0]   leading_zero_count_sgn; 
  logic                               lzc_zeroes;             
  logic        [SHIFT_AMOUNT_WIDTH-1:0] norm_shamt; 
  logic signed [EXP_WIDTH-1:0]          normalized_exponent;
  logic [3*PRECISION_BITS+4:0] sum_shifted;       
  logic [PRECISION_BITS:0]     final_mantissa;    
  logic [2*PRECISION_BITS+2:0] sum_sticky_bits;   
  logic                        sticky_after_norm; 
  logic signed [EXP_WIDTH-1:0] final_exponent;
  assign sum_lower = sum_q[LOWER_SUM_WIDTH-1:0];
  
  lzc #(
    .WIDTH ( LOWER_SUM_WIDTH ),
    .MODE  ( 1               ) 
  ) i_lzc (
    .in_i    ( sum_lower          ),
    .cnt_o   ( leading_zero_count ),
    .empty_o ( lzc_zeroes         )
  );
  assign leading_zero_count_sgn = signed'({1'b0, leading_zero_count});
  
  always_comb begin : norm_shift_amount
    
    if ((exponent_difference_q <= 0) || (effective_subtraction_q && (exponent_difference_q <= 2))) begin
      
      if ((exponent_product_q - leading_zero_count_sgn + 1 >= 0) && !lzc_zeroes) begin
        
        norm_shamt          = PRECISION_BITS + 2 + leading_zero_count;
        normalized_exponent = exponent_product_q - leading_zero_count_sgn + 1; 
      
      end else begin
        
        norm_shamt          = unsigned'(signed'(PRECISION_BITS) + 2 + exponent_product_q);
        normalized_exponent = 0; 
      end
    
    end else begin
      norm_shamt          = addend_shamt_q; 
      normalized_exponent = tentative_exponent_q;
    end
  end
  
  assign sum_shifted       = sum_q << norm_shamt;
  
  
  always_comb begin : small_norm
    
    {final_mantissa, sum_sticky_bits} = sum_shifted;
    final_exponent                    = normalized_exponent;
    
    if (sum_shifted[3*PRECISION_BITS+4]) begin 
      {final_mantissa, sum_sticky_bits} = sum_shifted >> 1;
      final_exponent                    = normalized_exponent + 1;
    
    end else if (sum_shifted[3*PRECISION_BITS+3]) begin 
      
    
    end else if (normalized_exponent > 1) begin
      {final_mantissa, sum_sticky_bits} = sum_shifted << 1;
      final_exponent                    = normalized_exponent - 1;
    
    end else begin
      final_exponent = '0;
    end
  end
  
  assign sticky_after_norm = (| {sum_sticky_bits}) | sticky_before_add_q;
  
  
  
  logic                         pre_round_sign;
  logic [EXP_BITS-1:0]          pre_round_exponent;
  logic [MAN_BITS-1:0]          pre_round_mantissa;
  logic [EXP_BITS+MAN_BITS-1:0] pre_round_abs; 
  logic [1:0]                   round_sticky_bits;
  logic of_before_round, of_after_round; 
  logic uf_before_round, uf_after_round; 
  logic result_zero;
  logic                         rounded_sign;
  logic [EXP_BITS+MAN_BITS-1:0] rounded_abs; 
  
  assign of_before_round = final_exponent >= 2**(EXP_BITS)-1; 
  assign uf_before_round = final_exponent == 0;               
  
  assign pre_round_sign     = final_sign_q;
  assign pre_round_exponent = (of_before_round) ? 2**EXP_BITS-2 : unsigned'(final_exponent[EXP_BITS-1:0]);
  assign pre_round_mantissa = (of_before_round) ? '1 : final_mantissa[MAN_BITS:1]; 
  assign pre_round_abs      = {pre_round_exponent, pre_round_mantissa};
  
  assign round_sticky_bits  = (of_before_round) ? 2'b11 : {final_mantissa[0], sticky_after_norm};
  
  fpnew_rounding #(
    .AbsWidth ( EXP_BITS + MAN_BITS )
  ) i_fpnew_rounding (
    .abs_value_i             ( pre_round_abs           ),
    .sign_i                  ( pre_round_sign          ),
    .round_sticky_bits_i     ( round_sticky_bits       ),
    .rnd_mode_i              ( rnd_mode_q              ),
    .effective_subtraction_i ( effective_subtraction_q ),
    .abs_rounded_o           ( rounded_abs             ),
    .sign_o                  ( rounded_sign            ),
    .exact_zero_o            ( result_zero             )
  );
  
  assign uf_after_round = rounded_abs[EXP_BITS+MAN_BITS-1:MAN_BITS] == '0; 
  assign of_after_round = rounded_abs[EXP_BITS+MAN_BITS-1:MAN_BITS] == '1; 
  
  
  
  logic [WIDTH-1:0]     regular_result;
  fpnew_pkg::status_t   regular_status;
  
  assign regular_result    = {rounded_sign, rounded_abs};
  assign regular_status.NV = 1'b0; 
  assign regular_status.DZ = 1'b0; 
  assign regular_status.OF = of_before_round | of_after_round;   
  assign regular_status.UF = uf_after_round & regular_status.NX; 
  assign regular_status.NX = (| round_sticky_bits) | of_before_round | of_after_round;
  
  fp_t                result_d;
  fpnew_pkg::status_t status_d;
  
  assign result_d = result_is_special_q ? special_result_q : regular_result;
  assign status_d = result_is_special_q ? special_status_q : regular_status;
  
  
  
  
  fp_t                [0:NUM_OUT_REGS] out_pipe_result_q;
  fpnew_pkg::status_t [0:NUM_OUT_REGS] out_pipe_status_q;
  TagType             [0:NUM_OUT_REGS] out_pipe_tag_q;
  AuxType             [0:NUM_OUT_REGS] out_pipe_aux_q;
  logic               [0:NUM_OUT_REGS] out_pipe_valid_q;
  
  logic [0:NUM_OUT_REGS] out_pipe_ready;
  
  assign out_pipe_result_q[0] = result_d;
  assign out_pipe_status_q[0] = status_d;
  assign out_pipe_tag_q[0]    = mid_pipe_tag_q[NUM_MID_REGS];
  assign out_pipe_aux_q[0]    = mid_pipe_aux_q[NUM_MID_REGS];
  assign out_pipe_valid_q[0]  = mid_pipe_valid_q[NUM_MID_REGS];
  
  assign mid_pipe_ready[NUM_MID_REGS] = out_pipe_ready[0];
  
  for (genvar i = 0; i < NUM_OUT_REGS; i++) begin : gen_output_pipeline
    
    logic reg_ena;
    
    
    
    assign out_pipe_ready[i] = out_pipe_ready[i+1] | ~out_pipe_valid_q[i+1];
    
    
                           
                         
                            
  always_ff @(posedge (clk_i) or negedge (rst_ni)) begin                 
    if (!rst_ni) begin                                                   
      out_pipe_valid_q[i+1] <= (1'b0);                                              
    end else begin                                                         
      out_pipe_valid_q[i+1] <= (flush_i) ? (1'b0) : (out_pipe_ready[i]) ? (out_pipe_valid_q[i]) : (out_pipe_valid_q[i+1]);       
    end                                                                    
  end
    
    assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
    
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_result_q[i+1] <= ('0);                        
    end else begin                                   
      out_pipe_result_q[i+1] <= (reg_ena) ? (out_pipe_result_q[i]) : (out_pipe_result_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_status_q[i+1] <= ('0);                        
    end else begin                                   
      out_pipe_status_q[i+1] <= (reg_ena) ? (out_pipe_status_q[i]) : (out_pipe_status_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_tag_q[i+1] <= (TagType'('0));                        
    end else begin                                   
      out_pipe_tag_q[i+1] <= (reg_ena) ? (out_pipe_tag_q[i]) : (out_pipe_tag_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_aux_q[i+1] <= (AuxType'('0));                        
    end else begin                                   
      out_pipe_aux_q[i+1] <= (reg_ena) ? (out_pipe_aux_q[i]) : (out_pipe_aux_q[i+1]);               
    end                                              
  end
  end
  
  assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
  
  assign result_o        = out_pipe_result_q[NUM_OUT_REGS];
  assign status_o        = out_pipe_status_q[NUM_OUT_REGS];
  assign extension_bit_o = 1'b1; 
  assign tag_o           = out_pipe_tag_q[NUM_OUT_REGS];
  assign aux_o           = out_pipe_aux_q[NUM_OUT_REGS];
  assign out_valid_o     = out_pipe_valid_q[NUM_OUT_REGS];
  assign busy_o          = (| {inp_pipe_valid_q, mid_pipe_valid_q, out_pipe_valid_q});
endmodule
                                      
module fpnew_noncomp #(
  parameter fpnew_pkg::fp_format_e   FpFormat    = fpnew_pkg::fp_format_e'(0),
  parameter int unsigned             NumPipeRegs = 0,
  parameter fpnew_pkg::pipe_config_t PipeConfig  = fpnew_pkg::BEFORE,
  parameter type                     TagType     = logic,
  parameter type                     AuxType     = logic,
  localparam int unsigned WIDTH = fpnew_pkg::fp_width(FpFormat) 
) (
  input logic                  clk_i,
  input logic                  rst_ni,
  
  input logic [1:0][WIDTH-1:0]     operands_i, 
  input logic [1:0]                is_boxed_i, 
  input fpnew_pkg::roundmode_e     rnd_mode_i,
  input fpnew_pkg::operation_e     op_i,
  input logic                      op_mod_i,
  input TagType                    tag_i,
  input AuxType                    aux_i,
  
  input  logic                     in_valid_i,
  output logic                     in_ready_o,
  input  logic                     flush_i,
  
  output logic [WIDTH-1:0]         result_o,
  output fpnew_pkg::status_t       status_o,
  output logic                     extension_bit_o,
  output fpnew_pkg::classmask_e    class_mask_o,
  output logic                     is_class_o,
  output TagType                   tag_o,
  output AuxType                   aux_o,
  
  output logic                     out_valid_o,
  input  logic                     out_ready_i,
  
  output logic                     busy_o
);
  
  
  
  localparam int unsigned EXP_BITS = fpnew_pkg::exp_bits(FpFormat);
  localparam int unsigned MAN_BITS = fpnew_pkg::man_bits(FpFormat);
  
  localparam NUM_INP_REGS = (PipeConfig == fpnew_pkg::BEFORE || PipeConfig == fpnew_pkg::INSIDE)
                            ? NumPipeRegs
                            : (PipeConfig == fpnew_pkg::DISTRIBUTED
                               ? ((NumPipeRegs + 1) / 2) 
                               : 0); 
  localparam NUM_OUT_REGS = PipeConfig == fpnew_pkg::AFTER
                            ? NumPipeRegs
                            : (PipeConfig == fpnew_pkg::DISTRIBUTED
                               ? (NumPipeRegs / 2) 
                               : 0); 
  
  
  
  typedef struct packed {
    logic                sign;
    logic [EXP_BITS-1:0] exponent;
    logic [MAN_BITS-1:0] mantissa;
  } fp_t;
  
  
  
  
  logic                  [0:NUM_INP_REGS][1:0][WIDTH-1:0] inp_pipe_operands_q;
  logic                  [0:NUM_INP_REGS][1:0]            inp_pipe_is_boxed_q;
  fpnew_pkg::roundmode_e [0:NUM_INP_REGS]                 inp_pipe_rnd_mode_q;
  fpnew_pkg::operation_e [0:NUM_INP_REGS]                 inp_pipe_op_q;
  logic                  [0:NUM_INP_REGS]                 inp_pipe_op_mod_q;
  TagType                [0:NUM_INP_REGS]                 inp_pipe_tag_q;
  AuxType                [0:NUM_INP_REGS]                 inp_pipe_aux_q;
  logic                  [0:NUM_INP_REGS]                 inp_pipe_valid_q;
  
  logic [0:NUM_INP_REGS] inp_pipe_ready;
  
  assign inp_pipe_operands_q[0] = operands_i;
  assign inp_pipe_is_boxed_q[0] = is_boxed_i;
  assign inp_pipe_rnd_mode_q[0] = rnd_mode_i;
  assign inp_pipe_op_q[0]       = op_i;
  assign inp_pipe_op_mod_q[0]   = op_mod_i;
  assign inp_pipe_tag_q[0]      = tag_i;
  assign inp_pipe_aux_q[0]      = aux_i;
  assign inp_pipe_valid_q[0]    = in_valid_i;
  
  assign in_ready_o = inp_pipe_ready[0];
  
  for (genvar i = 0; i < NUM_INP_REGS; i++) begin : gen_input_pipeline
    
    logic reg_ena;
    
    
    
    assign inp_pipe_ready[i] = inp_pipe_ready[i+1] | ~inp_pipe_valid_q[i+1];
    
    
                           
                         
                            
  always_ff @(posedge (clk_i) or negedge (rst_ni)) begin                 
    if (!rst_ni) begin                                                   
      inp_pipe_valid_q[i+1] <= (1'b0);                                              
    end else begin                                                         
      inp_pipe_valid_q[i+1] <= (flush_i) ? (1'b0) : (inp_pipe_ready[i]) ? (inp_pipe_valid_q[i]) : (inp_pipe_valid_q[i+1]);       
    end                                                                    
  end
    
    assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
    
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_operands_q[i+1] <= ('0);                        
    end else begin                                   
      inp_pipe_operands_q[i+1] <= (reg_ena) ? (inp_pipe_operands_q[i]) : (inp_pipe_operands_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_is_boxed_q[i+1] <= ('0);                        
    end else begin                                   
      inp_pipe_is_boxed_q[i+1] <= (reg_ena) ? (inp_pipe_is_boxed_q[i]) : (inp_pipe_is_boxed_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_rnd_mode_q[i+1] <= (fpnew_pkg::RNE);                        
    end else begin                                   
      inp_pipe_rnd_mode_q[i+1] <= (reg_ena) ? (inp_pipe_rnd_mode_q[i]) : (inp_pipe_rnd_mode_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_op_q[i+1] <= (fpnew_pkg::FMADD);                        
    end else begin                                   
      inp_pipe_op_q[i+1] <= (reg_ena) ? (inp_pipe_op_q[i]) : (inp_pipe_op_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_op_mod_q[i+1] <= ('0);                        
    end else begin                                   
      inp_pipe_op_mod_q[i+1] <= (reg_ena) ? (inp_pipe_op_mod_q[i]) : (inp_pipe_op_mod_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_tag_q[i+1] <= (TagType'('0));                        
    end else begin                                   
      inp_pipe_tag_q[i+1] <= (reg_ena) ? (inp_pipe_tag_q[i]) : (inp_pipe_tag_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      inp_pipe_aux_q[i+1] <= (AuxType'('0));                        
    end else begin                                   
      inp_pipe_aux_q[i+1] <= (reg_ena) ? (inp_pipe_aux_q[i]) : (inp_pipe_aux_q[i+1]);               
    end                                              
  end
  end
  
  
  
  fpnew_pkg::fp_info_t [1:0] info_q;
  
  fpnew_classifier #(
    .FpFormat    ( FpFormat ),
    .NumOperands ( 2        )
    ) i_class_a (
    .operands_i ( inp_pipe_operands_q[NUM_INP_REGS] ),
    .is_boxed_i ( inp_pipe_is_boxed_q[NUM_INP_REGS] ),
    .info_o     ( info_q                            )
  );
  fp_t                 operand_a, operand_b;
  fpnew_pkg::fp_info_t info_a,    info_b;
  
  assign operand_a = inp_pipe_operands_q[NUM_INP_REGS][0];
  assign operand_b = inp_pipe_operands_q[NUM_INP_REGS][1];
  assign info_a    = info_q[0];
  assign info_b    = info_q[1];
  logic any_operand_inf;
  logic any_operand_nan;
  logic signalling_nan;
  
  assign any_operand_inf = (| {info_a.is_inf,        info_b.is_inf});
  assign any_operand_nan = (| {info_a.is_nan,        info_b.is_nan});
  assign signalling_nan  = (| {info_a.is_signalling, info_b.is_signalling});
  logic operands_equal, operand_a_smaller;
  
  assign operands_equal    = (operand_a == operand_b) || (info_a.is_zero && info_b.is_zero);
  
  assign operand_a_smaller = (operand_a < operand_b) ^ (operand_a.sign || operand_b.sign);
  
  
  
  fp_t                sgnj_result;
  fpnew_pkg::status_t sgnj_status;
  logic               sgnj_extension_bit;
  
  
  always_comb begin : sign_injections
    logic sign_a, sign_b; 
    
    sgnj_result = operand_a; 
    
    if (!info_a.is_boxed) sgnj_result = '{sign: 1'b0, exponent: '1, mantissa: 2**(MAN_BITS-1)};
    
    sign_a = operand_a.sign & info_a.is_boxed;
    sign_b = operand_b.sign & info_b.is_boxed;
    
    unique case (inp_pipe_rnd_mode_q[NUM_INP_REGS])
      fpnew_pkg::RNE: sgnj_result.sign = sign_b;          
      fpnew_pkg::RTZ: sgnj_result.sign = ~sign_b;         
      fpnew_pkg::RDN: sgnj_result.sign = sign_a ^ sign_b; 
      fpnew_pkg::RUP: sgnj_result      = operand_a;       
      default: sgnj_result = '{default: fpnew_pkg::DONT_CARE}; 
    endcase
  end
  assign sgnj_status = '0;        
  
  assign sgnj_extension_bit = inp_pipe_op_mod_q[NUM_INP_REGS] ? sgnj_result.sign : 1'b1;
  
  
  
  fp_t                minmax_result;
  fpnew_pkg::status_t minmax_status;
  logic               minmax_extension_bit;
  
  
  always_comb begin : min_max
    
    minmax_status = '0;
    
    minmax_status.NV = signalling_nan;
    
    if (info_a.is_nan && info_b.is_nan)
      minmax_result = '{sign: 1'b0, exponent: '1, mantissa: 2**(MAN_BITS-1)}; 
    
    else if (info_a.is_nan) minmax_result = operand_b;
    else if (info_b.is_nan) minmax_result = operand_a;
    
    else begin
      unique case (inp_pipe_rnd_mode_q[NUM_INP_REGS])
        fpnew_pkg::RNE: minmax_result = operand_a_smaller ? operand_a : operand_b; 
        fpnew_pkg::RTZ: minmax_result = operand_a_smaller ? operand_b : operand_a; 
        default: minmax_result = '{default: fpnew_pkg::DONT_CARE}; 
      endcase
    end
  end
  assign minmax_extension_bit = 1'b1; 
  
  
  
  fp_t                cmp_result;
  fpnew_pkg::status_t cmp_status;
  logic               cmp_extension_bit;
  
  
  
  always_comb begin : comparisons
    
    cmp_result = '0; 
    cmp_status = '0; 
    
    if (signalling_nan) cmp_status.NV = 1'b1; 
    
    else begin
      unique case (inp_pipe_rnd_mode_q[NUM_INP_REGS])
        fpnew_pkg::RNE: begin 
          if (any_operand_nan) cmp_status.NV = 1'b1; 
          else cmp_result = (operand_a_smaller | operands_equal) ^ inp_pipe_op_mod_q[NUM_INP_REGS];
        end
        fpnew_pkg::RTZ: begin 
          if (any_operand_nan) cmp_status.NV = 1'b1; 
          else cmp_result = (operand_a_smaller & ~operands_equal) ^ inp_pipe_op_mod_q[NUM_INP_REGS];
        end
        fpnew_pkg::RDN: begin 
          if (any_operand_nan) cmp_result = inp_pipe_op_mod_q[NUM_INP_REGS]; 
          else cmp_result = operands_equal ^ inp_pipe_op_mod_q[NUM_INP_REGS];
        end
        default: cmp_result = '{default: fpnew_pkg::DONT_CARE}; 
      endcase
    end
  end
  assign cmp_extension_bit = 1'b0; 
  
  
  
  fpnew_pkg::status_t    class_status;
  logic                  class_extension_bit;
  fpnew_pkg::classmask_e class_mask_d; 
  
  always_comb begin : classify
    if (info_a.is_normal) begin
      class_mask_d = operand_a.sign       ? fpnew_pkg::NEGNORM    : fpnew_pkg::POSNORM;
    end else if (info_a.is_subnormal) begin
      class_mask_d = operand_a.sign       ? fpnew_pkg::NEGSUBNORM : fpnew_pkg::POSSUBNORM;
    end else if (info_a.is_zero) begin
      class_mask_d = operand_a.sign       ? fpnew_pkg::NEGZERO    : fpnew_pkg::POSZERO;
    end else if (info_a.is_inf) begin
      class_mask_d = operand_a.sign       ? fpnew_pkg::NEGINF     : fpnew_pkg::POSINF;
    end else if (info_a.is_nan) begin
      class_mask_d = info_a.is_signalling ? fpnew_pkg::SNAN       : fpnew_pkg::QNAN;
    end else begin
      class_mask_d = fpnew_pkg::QNAN; 
    end
  end
  assign class_status        = '0;   
  assign class_extension_bit = 1'b0; 
  
  
  
  fp_t                   result_d;
  fpnew_pkg::status_t    status_d;
  logic                  extension_bit_d;
  logic                  is_class_d;
  
  always_comb begin : select_result
    unique case (inp_pipe_op_q[NUM_INP_REGS])
      fpnew_pkg::SGNJ: begin
        result_d        = sgnj_result;
        status_d        = sgnj_status;
        extension_bit_d = sgnj_extension_bit;
      end
      fpnew_pkg::MINMAX: begin
        result_d        = minmax_result;
        status_d        = minmax_status;
        extension_bit_d = minmax_extension_bit;
      end
      fpnew_pkg::CMP: begin
        result_d        = cmp_result;
        status_d        = cmp_status;
        extension_bit_d = cmp_extension_bit;
      end
      fpnew_pkg::CLASSIFY: begin
        result_d        = '{default: fpnew_pkg::DONT_CARE}; 
        status_d        = class_status;
        extension_bit_d = class_extension_bit;
      end
      default: begin
        result_d        = '{default: fpnew_pkg::DONT_CARE}; 
        status_d        = '{default: fpnew_pkg::DONT_CARE}; 
        extension_bit_d = fpnew_pkg::DONT_CARE;             
      end
    endcase
  end
  assign is_class_d = (inp_pipe_op_q[NUM_INP_REGS] == fpnew_pkg::CLASSIFY);
  
  
  
  
  fp_t                   [0:NUM_OUT_REGS] out_pipe_result_q;
  fpnew_pkg::status_t    [0:NUM_OUT_REGS] out_pipe_status_q;
  logic                  [0:NUM_OUT_REGS] out_pipe_extension_bit_q;
  fpnew_pkg::classmask_e [0:NUM_OUT_REGS] out_pipe_class_mask_q;
  logic                  [0:NUM_OUT_REGS] out_pipe_is_class_q;
  TagType                [0:NUM_OUT_REGS] out_pipe_tag_q;
  AuxType                [0:NUM_OUT_REGS] out_pipe_aux_q;
  logic                  [0:NUM_OUT_REGS] out_pipe_valid_q;
  
  logic [0:NUM_OUT_REGS] out_pipe_ready;
  
  assign out_pipe_result_q[0]        = result_d;
  assign out_pipe_status_q[0]        = status_d;
  assign out_pipe_extension_bit_q[0] = extension_bit_d;
  assign out_pipe_class_mask_q[0]    = class_mask_d;
  assign out_pipe_is_class_q[0]      = is_class_d;
  assign out_pipe_tag_q[0]           = inp_pipe_tag_q[NUM_INP_REGS];
  assign out_pipe_aux_q[0]           = inp_pipe_aux_q[NUM_INP_REGS];
  assign out_pipe_valid_q[0]         = inp_pipe_valid_q[NUM_INP_REGS];
  
  assign inp_pipe_ready[NUM_INP_REGS] = out_pipe_ready[0];
  
  for (genvar i = 0; i < NUM_OUT_REGS; i++) begin : gen_output_pipeline
    
    logic reg_ena;
    
    
    
    assign out_pipe_ready[i] = out_pipe_ready[i+1] | ~out_pipe_valid_q[i+1];
    
    
                           
                         
                            
  always_ff @(posedge (clk_i) or negedge (rst_ni)) begin                 
    if (!rst_ni) begin                                                   
      out_pipe_valid_q[i+1] <= (1'b0);                                              
    end else begin                                                         
      out_pipe_valid_q[i+1] <= (flush_i) ? (1'b0) : (out_pipe_ready[i]) ? (out_pipe_valid_q[i]) : (out_pipe_valid_q[i+1]);       
    end                                                                    
  end
    
    assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
    
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_result_q[i+1] <= ('0);                        
    end else begin                                   
      out_pipe_result_q[i+1] <= (reg_ena) ? (out_pipe_result_q[i]) : (out_pipe_result_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_status_q[i+1] <= ('0);                        
    end else begin                                   
      out_pipe_status_q[i+1] <= (reg_ena) ? (out_pipe_status_q[i]) : (out_pipe_status_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_extension_bit_q[i+1] <= ('0);                        
    end else begin                                   
      out_pipe_extension_bit_q[i+1] <= (reg_ena) ? (out_pipe_extension_bit_q[i]) : (out_pipe_extension_bit_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_class_mask_q[i+1] <= (fpnew_pkg::QNAN);                        
    end else begin                                   
      out_pipe_class_mask_q[i+1] <= (reg_ena) ? (out_pipe_class_mask_q[i]) : (out_pipe_class_mask_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_is_class_q[i+1] <= ('0);                        
    end else begin                                   
      out_pipe_is_class_q[i+1] <= (reg_ena) ? (out_pipe_is_class_q[i]) : (out_pipe_is_class_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_tag_q[i+1] <= (TagType'('0));                        
    end else begin                                   
      out_pipe_tag_q[i+1] <= (reg_ena) ? (out_pipe_tag_q[i]) : (out_pipe_tag_q[i+1]);               
    end                                              
  end
    
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      out_pipe_aux_q[i+1] <= (AuxType'('0));                        
    end else begin                                   
      out_pipe_aux_q[i+1] <= (reg_ena) ? (out_pipe_aux_q[i]) : (out_pipe_aux_q[i+1]);               
    end                                              
  end
  end
  
  assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
  
  assign result_o        = out_pipe_result_q[NUM_OUT_REGS];
  assign status_o        = out_pipe_status_q[NUM_OUT_REGS];
  assign extension_bit_o = out_pipe_extension_bit_q[NUM_OUT_REGS];
  assign class_mask_o    = out_pipe_class_mask_q[NUM_OUT_REGS];
  assign is_class_o      = out_pipe_is_class_q[NUM_OUT_REGS];
  assign tag_o           = out_pipe_tag_q[NUM_OUT_REGS];
  assign aux_o           = out_pipe_aux_q[NUM_OUT_REGS];
  assign out_valid_o     = out_pipe_valid_q[NUM_OUT_REGS];
  assign busy_o          = (| {inp_pipe_valid_q, out_pipe_valid_q});
endmodule
module fpnew_opgroup_block #(
  parameter fpnew_pkg::opgroup_e        OpGroup       = fpnew_pkg::ADDMUL,
  
  parameter int unsigned                Width         = 32,
  parameter logic                       EnableVectors = 1'b1,
  parameter fpnew_pkg::fmt_logic_t      FpFmtMask     = '1,
  parameter fpnew_pkg::ifmt_logic_t     IntFmtMask    = '1,
  parameter fpnew_pkg::fmt_unsigned_t   FmtPipeRegs   = '{default: 0},
  parameter fpnew_pkg::fmt_unit_types_t FmtUnitTypes  = '{default: fpnew_pkg::PARALLEL},
  parameter fpnew_pkg::pipe_config_t    PipeConfig    = fpnew_pkg::BEFORE,
  parameter type                        TagType       = logic,
  
  localparam int unsigned NUM_FORMATS  = fpnew_pkg::NUM_FP_FORMATS,
  localparam int unsigned NUM_OPERANDS = fpnew_pkg::num_operands(OpGroup)
) (
  input logic                                     clk_i,
  input logic                                     rst_ni,
  
  input logic [NUM_OPERANDS-1:0][Width-1:0]       operands_i,
  input logic [NUM_FORMATS-1:0][NUM_OPERANDS-1:0] is_boxed_i,
  input fpnew_pkg::roundmode_e                    rnd_mode_i,
  input fpnew_pkg::operation_e                    op_i,
  input logic                                     op_mod_i,
  input fpnew_pkg::fp_format_e                    src_fmt_i,
  input fpnew_pkg::fp_format_e                    dst_fmt_i,
  input fpnew_pkg::int_format_e                   int_fmt_i,
  input logic                                     vectorial_op_i,
  input TagType                                   tag_i,
  
  input  logic                                    in_valid_i,
  output logic                                    in_ready_o,
  input  logic                                    flush_i,
  
  output logic [Width-1:0]                        result_o,
  output fpnew_pkg::status_t                      status_o,
  output logic                                    extension_bit_o,
  output TagType                                  tag_o,
  
  output logic                                    out_valid_o,
  input  logic                                    out_ready_i,
  
  output logic                                    busy_o
);
  
  
  
  typedef struct packed {
    logic [Width-1:0]   result;
    fpnew_pkg::status_t status;
    logic               ext_bit;
    TagType             tag;
  } output_t;
  
  logic [NUM_FORMATS-1:0] fmt_in_ready, fmt_out_valid, fmt_out_ready, fmt_busy;
  output_t [NUM_FORMATS-1:0] fmt_outputs;
  
  
  
  assign in_ready_o = in_valid_i & fmt_in_ready[dst_fmt_i]; 
  
  
  
  for (genvar fmt = 0; fmt < int'(NUM_FORMATS); fmt++) begin : gen_parallel_slices
    
    localparam logic ANY_MERGED = fpnew_pkg::any_enabled_multi(FmtUnitTypes, FpFmtMask);
    localparam logic IS_FIRST_MERGED =
        fpnew_pkg::is_first_enabled_multi(fpnew_pkg::fp_format_e'(fmt), FmtUnitTypes, FpFmtMask);
    
    if (FpFmtMask[fmt] && (FmtUnitTypes[fmt] == fpnew_pkg::PARALLEL)) begin : active_format
      logic in_valid;
      assign in_valid = in_valid_i & (dst_fmt_i == fmt); 
      fpnew_opgroup_fmt_slice #(
        .OpGroup       ( OpGroup                      ),
        .FpFormat      ( fpnew_pkg::fp_format_e'(fmt) ),
        .Width         ( Width                        ),
        .EnableVectors ( EnableVectors                ),
        .NumPipeRegs   ( FmtPipeRegs[fmt]             ),
        .PipeConfig    ( PipeConfig                   ),
        .TagType       ( TagType                      )
      ) i_fmt_slice (
        .clk_i,
        .rst_ni,
        .operands_i     ( operands_i               ),
        .is_boxed_i     ( is_boxed_i[fmt]          ),
        .rnd_mode_i,
        .op_i,
        .op_mod_i,
        .vectorial_op_i,
        .tag_i,
        .in_valid_i     ( in_valid                 ),
        .in_ready_o     ( fmt_in_ready[fmt]        ),
        .flush_i,
        .result_o       ( fmt_outputs[fmt].result  ),
        .status_o       ( fmt_outputs[fmt].status  ),
        .extension_bit_o( fmt_outputs[fmt].ext_bit ),
        .tag_o          ( fmt_outputs[fmt].tag     ),
        .out_valid_o    ( fmt_out_valid[fmt]       ),
        .out_ready_i    ( fmt_out_ready[fmt]       ),
        .busy_o         ( fmt_busy[fmt]            )
      );
    
    end else if (FpFmtMask[fmt] && ANY_MERGED && !IS_FIRST_MERGED) begin : merged_unused
      
      assign fmt_in_ready[fmt]  = fmt_in_ready[fpnew_pkg::get_first_enabled_multi(FmtUnitTypes,
                                                                                  FpFmtMask)];
      assign fmt_out_valid[fmt] = 1'b0; 
      assign fmt_busy[fmt]      = 1'b0; 
      
      assign fmt_outputs[fmt].result  = '{default: fpnew_pkg::DONT_CARE};
      assign fmt_outputs[fmt].status  = '{default: fpnew_pkg::DONT_CARE};
      assign fmt_outputs[fmt].ext_bit = fpnew_pkg::DONT_CARE;
      assign fmt_outputs[fmt].tag     = TagType'(fpnew_pkg::DONT_CARE);
    
    end else if (!FpFmtMask[fmt] || (FmtUnitTypes[fmt] == fpnew_pkg::DISABLED)) begin : disable_fmt
      assign fmt_in_ready[fmt]  = 1'b0; 
      assign fmt_out_valid[fmt] = 1'b0; 
      assign fmt_busy[fmt]      = 1'b0; 
      
      assign fmt_outputs[fmt].result  = '{default: fpnew_pkg::DONT_CARE};
      assign fmt_outputs[fmt].status  = '{default: fpnew_pkg::DONT_CARE};
      assign fmt_outputs[fmt].ext_bit = fpnew_pkg::DONT_CARE;
      assign fmt_outputs[fmt].tag     = TagType'(fpnew_pkg::DONT_CARE);
    end
  end
  
  
  
  if (fpnew_pkg::any_enabled_multi(FmtUnitTypes, FpFmtMask)) begin : gen_merged_slice
    localparam FMT = fpnew_pkg::get_first_enabled_multi(FmtUnitTypes, FpFmtMask);
    localparam REG = fpnew_pkg::get_num_regs_multi(FmtPipeRegs, FmtUnitTypes, FpFmtMask);
    logic in_valid;
    assign in_valid = in_valid_i & (FmtUnitTypes[dst_fmt_i] == fpnew_pkg::MERGED);
    fpnew_opgroup_multifmt_slice #(
      .OpGroup       ( OpGroup          ),
      .Width         ( Width            ),
      .FpFmtConfig   ( FpFmtMask        ),
      .IntFmtConfig  ( IntFmtMask       ),
      .EnableVectors ( EnableVectors    ),
      .NumPipeRegs   ( REG              ),
      .PipeConfig    ( PipeConfig       ),
      .TagType       ( TagType          )
    ) i_multifmt_slice (
      .clk_i,
      .rst_ni,
      .operands_i,
      .is_boxed_i,
      .rnd_mode_i,
      .op_i,
      .op_mod_i,
      .src_fmt_i,
      .dst_fmt_i,
      .int_fmt_i,
      .vectorial_op_i,
      .tag_i,
      .in_valid_i      ( in_valid                 ),
      .in_ready_o      ( fmt_in_ready[FMT]        ),
      .flush_i,
      .result_o        ( fmt_outputs[FMT].result  ),
      .status_o        ( fmt_outputs[FMT].status  ),
      .extension_bit_o ( fmt_outputs[FMT].ext_bit ),
      .tag_o           ( fmt_outputs[FMT].tag     ),
      .out_valid_o     ( fmt_out_valid[FMT]       ),
      .out_ready_i     ( fmt_out_ready[FMT]       ),
      .busy_o          ( fmt_busy[FMT]            )
    );
  end
  
  
  
  output_t arbiter_output;
  
  rr_arb_tree #(
    .NumIn     ( NUM_FORMATS ),
    .DataType  ( output_t    ),
    .AxiVldRdy ( 1'b1        )
  ) i_arbiter (
    .clk_i,
    .rst_ni,
    .flush_i,
    .rr_i   ( '0             ),
    .req_i  ( fmt_out_valid  ),
    .gnt_o  ( fmt_out_ready  ),
    .data_i ( fmt_outputs    ),
    .gnt_i  ( out_ready_i    ),
    .req_o  ( out_valid_o    ),
    .data_o ( arbiter_output ),
    .idx_o  (    )
  );
  
  assign result_o        = arbiter_output.result;
  assign status_o        = arbiter_output.status;
  assign extension_bit_o = arbiter_output.ext_bit;
  assign tag_o           = arbiter_output.tag;
  assign busy_o = (| fmt_busy);
endmodule
module fpnew_opgroup_fmt_slice #(
  parameter fpnew_pkg::opgroup_e     OpGroup       = fpnew_pkg::ADDMUL,
  parameter fpnew_pkg::fp_format_e   FpFormat      = fpnew_pkg::fp_format_e'(0),
  
  parameter int unsigned             Width         = 32,
  parameter logic                    EnableVectors = 1'b1,
  parameter int unsigned             NumPipeRegs   = 0,
  parameter fpnew_pkg::pipe_config_t PipeConfig    = fpnew_pkg::BEFORE,
  parameter type                     TagType       = logic,
  
  localparam int unsigned NUM_OPERANDS = fpnew_pkg::num_operands(OpGroup)
) (
  input logic                               clk_i,
  input logic                               rst_ni,
  
  input logic [NUM_OPERANDS-1:0][Width-1:0] operands_i,
  input logic [NUM_OPERANDS-1:0]            is_boxed_i,
  input fpnew_pkg::roundmode_e              rnd_mode_i,
  input fpnew_pkg::operation_e              op_i,
  input logic                               op_mod_i,
  input logic                               vectorial_op_i,
  input TagType                             tag_i,
  
  input  logic                              in_valid_i,
  output logic                              in_ready_o,
  input  logic                              flush_i,
  
  output logic [Width-1:0]                  result_o,
  output fpnew_pkg::status_t                status_o,
  output logic                              extension_bit_o,
  output TagType                            tag_o,
  
  output logic                              out_valid_o,
  input  logic                              out_ready_i,
  
  output logic                              busy_o
);
  localparam int unsigned FP_WIDTH  = fpnew_pkg::fp_width(FpFormat);
  localparam int unsigned NUM_LANES = fpnew_pkg::num_lanes(Width, FpFormat, EnableVectors);
  logic [NUM_LANES-1:0] lane_in_ready, lane_out_valid; 
  logic                 vectorial_op;
  logic [NUM_LANES*FP_WIDTH-1:0] slice_result;
  logic [Width-1:0]              slice_regular_result, slice_class_result, slice_vec_class_result;
  fpnew_pkg::status_t    [NUM_LANES-1:0] lane_status;
  logic                  [NUM_LANES-1:0] lane_ext_bit; 
  fpnew_pkg::classmask_e [NUM_LANES-1:0] lane_class_mask;
  TagType                [NUM_LANES-1:0] lane_tags; 
  logic                  [NUM_LANES-1:0] lane_vectorial, lane_busy, lane_is_class; 
  logic result_is_vector, result_is_class;
  
  
  
  assign in_ready_o   = lane_in_ready[0]; 
  assign vectorial_op = vectorial_op_i & EnableVectors; 
  
  
  
  for (genvar lane = 0; lane < int'(NUM_LANES); lane++) begin : gen_num_lanes
    logic [FP_WIDTH-1:0] local_result; 
    logic                local_sign;
    
    if ((lane == 0) || EnableVectors) begin : active_lane
      logic in_valid, out_valid, out_ready; 
      logic [NUM_OPERANDS-1:0][FP_WIDTH-1:0] local_operands; 
      logic [FP_WIDTH-1:0]                   op_result;      
      fpnew_pkg::status_t                    op_status;
      assign in_valid = in_valid_i & ((lane == 0) | vectorial_op); 
      
      always_comb begin : prepare_input
        for (int i = 0; i < int'(NUM_OPERANDS); i++) begin
          local_operands[i] = operands_i[i][(unsigned'(lane)+1)*FP_WIDTH-1:unsigned'(lane)*FP_WIDTH];
        end
      end
      
      if (OpGroup == fpnew_pkg::ADDMUL) begin : lane_instance
        fpnew_fma #(
          .FpFormat    ( FpFormat    ),
          .NumPipeRegs ( NumPipeRegs ),
          .PipeConfig  ( PipeConfig  ),
          .TagType     ( TagType     ),
          .AuxType     ( logic       )
        ) i_fma (
          .clk_i,
          .rst_ni,
          .operands_i      ( local_operands               ),
          .is_boxed_i      ( is_boxed_i[NUM_OPERANDS-1:0] ),
          .rnd_mode_i,
          .op_i,
          .op_mod_i,
          .tag_i,
          .aux_i           ( vectorial_op         ), 
          .in_valid_i      ( in_valid             ),
          .in_ready_o      ( lane_in_ready[lane]  ),
          .flush_i,
          .result_o        ( op_result            ),
          .status_o        ( op_status            ),
          .extension_bit_o ( lane_ext_bit[lane]   ),
          .tag_o           ( lane_tags[lane]      ),
          .aux_o           ( lane_vectorial[lane] ),
          .out_valid_o     ( out_valid            ),
          .out_ready_i     ( out_ready            ),
          .busy_o          ( lane_busy[lane]      )
        );
        assign lane_is_class[lane]   = 1'b0;
        assign lane_class_mask[lane] = fpnew_pkg::NEGINF;
      end else if (OpGroup == fpnew_pkg::DIVSQRT) begin : lane_instance
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
      end else if (OpGroup == fpnew_pkg::NONCOMP) begin : lane_instance
        fpnew_noncomp #(
          .FpFormat   (FpFormat),
          .NumPipeRegs(NumPipeRegs),
          .PipeConfig (PipeConfig),
          .TagType    (TagType),
          .AuxType    (logic)
        ) i_noncomp (
          .clk_i,
          .rst_ni,
          .operands_i      ( local_operands               ),
          .is_boxed_i      ( is_boxed_i[NUM_OPERANDS-1:0] ),
          .rnd_mode_i,
          .op_i,
          .op_mod_i,
          .tag_i,
          .aux_i           ( vectorial_op          ), 
          .in_valid_i      ( in_valid              ),
          .in_ready_o      ( lane_in_ready[lane]   ),
          .flush_i,
          .result_o        ( op_result             ),
          .status_o        ( op_status             ),
          .extension_bit_o ( lane_ext_bit[lane]    ),
          .class_mask_o    ( lane_class_mask[lane] ),
          .is_class_o      ( lane_is_class[lane]   ),
          .tag_o           ( lane_tags[lane]       ),
          .aux_o           ( lane_vectorial[lane]  ),
          .out_valid_o     ( out_valid             ),
          .out_ready_i     ( out_ready             ),
          .busy_o          ( lane_busy[lane]       )
        );
      end 
      
      assign out_ready            = out_ready_i & ((lane == 0) | result_is_vector);
      assign lane_out_valid[lane] = out_valid   & ((lane == 0) | result_is_vector);
      
      assign local_result      = lane_out_valid[lane] ? op_result : '{default: lane_ext_bit[0]};
      assign lane_status[lane] = lane_out_valid[lane] ? op_status : '0;
    
    end else begin
      assign lane_out_valid[lane] = 1'b0; 
      assign lane_in_ready[lane]  = 1'b0; 
      assign local_result         = '{default: lane_ext_bit[0]}; 
      assign lane_status[lane]    = '0;
      assign lane_busy[lane]      = 1'b0;
      assign lane_is_class[lane]  = 1'b0;
    end
    
    assign slice_result[(unsigned'(lane)+1)*FP_WIDTH-1:unsigned'(lane)*FP_WIDTH] = local_result;
    
    if ((lane+1)*8 <= Width) begin : vectorial_class 
      assign local_sign = (lane_class_mask[lane] == fpnew_pkg::NEGINF ||
                           lane_class_mask[lane] == fpnew_pkg::NEGNORM ||
                           lane_class_mask[lane] == fpnew_pkg::NEGSUBNORM ||
                           lane_class_mask[lane] == fpnew_pkg::NEGZERO);
      
      assign slice_vec_class_result[(lane+1)*8-1:lane*8] = {
        local_sign,  
        ~local_sign, 
        lane_class_mask[lane] == fpnew_pkg::QNAN, 
        lane_class_mask[lane] == fpnew_pkg::SNAN, 
        lane_class_mask[lane] == fpnew_pkg::POSZERO
            || lane_class_mask[lane] == fpnew_pkg::NEGZERO, 
        lane_class_mask[lane] == fpnew_pkg::POSSUBNORM
            || lane_class_mask[lane] == fpnew_pkg::NEGSUBNORM, 
        lane_class_mask[lane] == fpnew_pkg::POSNORM
            || lane_class_mask[lane] == fpnew_pkg::NEGNORM, 
        lane_class_mask[lane] == fpnew_pkg::POSINF
            || lane_class_mask[lane] == fpnew_pkg::NEGINF 
      };
    end
  end
  
  
  
  assign result_is_vector = lane_vectorial[0];
  assign result_is_class  = lane_is_class[0];
  assign slice_regular_result = $signed({extension_bit_o, slice_result});
  localparam int unsigned CLASS_VEC_BITS = (NUM_LANES*8 > Width) ? 8 * (Width / 8) : NUM_LANES*8;
  
  if (CLASS_VEC_BITS < Width) begin : pad_vectorial_class
    assign slice_vec_class_result[Width-1:CLASS_VEC_BITS] = '0;
  end
  
  assign slice_class_result = result_is_vector ? slice_vec_class_result : lane_class_mask[0];
  
  assign result_o = result_is_class ? slice_class_result : slice_regular_result;
  assign extension_bit_o                              = lane_ext_bit[0]; 
  assign tag_o                                        = lane_tags[0];    
  assign busy_o                                       = (| lane_busy);
  assign out_valid_o                                  = lane_out_valid[0]; 
  
  always_comb begin : output_processing
    
    automatic fpnew_pkg::status_t temp_status;
    temp_status = '0;
    for (int i = 0; i < int'(NUM_LANES); i++)
      temp_status |= lane_status[i];
    status_o = temp_status;
  end
endmodule
                                      
module fpnew_opgroup_multifmt_slice #(
  parameter fpnew_pkg::opgroup_e     OpGroup       = fpnew_pkg::CONV,
  parameter int unsigned             Width         = 64,
  
  parameter fpnew_pkg::fmt_logic_t   FpFmtConfig   = '1,
  parameter fpnew_pkg::ifmt_logic_t  IntFmtConfig  = '1,
  parameter logic                    EnableVectors = 1'b1,
  parameter int unsigned             NumPipeRegs   = 0,
  parameter fpnew_pkg::pipe_config_t PipeConfig    = fpnew_pkg::BEFORE,
  parameter type                     TagType       = logic,
  
  localparam int unsigned NUM_OPERANDS = fpnew_pkg::num_operands(OpGroup),
  localparam int unsigned NUM_FORMATS  = fpnew_pkg::NUM_FP_FORMATS
) (
  input logic                                     clk_i,
  input logic                                     rst_ni,
  
  input logic [NUM_OPERANDS-1:0][Width-1:0]       operands_i,
  input logic [NUM_FORMATS-1:0][NUM_OPERANDS-1:0] is_boxed_i,
  input fpnew_pkg::roundmode_e                    rnd_mode_i,
  input fpnew_pkg::operation_e                    op_i,
  input logic                                     op_mod_i,
  input fpnew_pkg::fp_format_e                    src_fmt_i,
  input fpnew_pkg::fp_format_e                    dst_fmt_i,
  input fpnew_pkg::int_format_e                   int_fmt_i,
  input logic                                     vectorial_op_i,
  input TagType                                   tag_i,
  
  input  logic                                    in_valid_i,
  output logic                                    in_ready_o,
  input  logic                                    flush_i,
  
  output logic [Width-1:0]                        result_o,
  output fpnew_pkg::status_t                      status_o,
  output logic                                    extension_bit_o,
  output TagType                                  tag_o,
  
  output logic                                    out_valid_o,
  input  logic                                    out_ready_i,
  
  output logic                                    busy_o
);
  localparam int unsigned MAX_FP_WIDTH   = fpnew_pkg::max_fp_width(FpFmtConfig);
  localparam int unsigned MAX_INT_WIDTH  = fpnew_pkg::max_int_width(IntFmtConfig);
  localparam int unsigned NUM_LANES = fpnew_pkg::max_num_lanes(Width, FpFmtConfig, 1'b1);
  localparam int unsigned NUM_INT_FORMATS = fpnew_pkg::NUM_INT_FORMATS;
  
  localparam int unsigned FMT_BITS =
      fpnew_pkg::maximum($clog2(NUM_FORMATS), $clog2(NUM_INT_FORMATS));
  localparam int unsigned AUX_BITS = FMT_BITS + 2; 
  logic [NUM_LANES-1:0] lane_in_ready, lane_out_valid; 
  logic                 vectorial_op;
  logic [FMT_BITS-1:0]  dst_fmt; 
  logic [AUX_BITS-1:0]  aux_data;
  
  logic       dst_fmt_is_int, dst_is_cpk;
  logic [1:0] dst_vec_op; 
  logic [2:0] target_aux_d, target_aux_q;
  logic       is_up_cast, is_down_cast;
  logic [NUM_FORMATS-1:0][Width-1:0]     fmt_slice_result;
  logic [NUM_INT_FORMATS-1:0][Width-1:0] ifmt_slice_result;
  logic [Width-1:0]                      conv_slice_result;
  logic [Width-1:0] conv_target_d, conv_target_q; 
  fpnew_pkg::status_t [NUM_LANES-1:0]   lane_status;
  logic   [NUM_LANES-1:0]               lane_ext_bit; 
  TagType [NUM_LANES-1:0]               lane_tags; 
  logic   [NUM_LANES-1:0][AUX_BITS-1:0] lane_aux; 
  logic   [NUM_LANES-1:0]               lane_busy; 
  logic                result_is_vector;
  logic [FMT_BITS-1:0] result_fmt;
  logic                result_fmt_is_int, result_is_cpk;
  logic [1:0]          result_vec_op; 
  
  
  
  assign in_ready_o   = lane_in_ready[0]; 
  assign vectorial_op = vectorial_op_i & EnableVectors; 
  
  assign dst_fmt_is_int = (OpGroup == fpnew_pkg::CONV) & (op_i == fpnew_pkg::F2I);
  assign dst_is_cpk     = (OpGroup == fpnew_pkg::CONV) & (op_i == fpnew_pkg::CPKAB ||
                                                          op_i == fpnew_pkg::CPKCD);
  assign dst_vec_op     = (OpGroup == fpnew_pkg::CONV) & {(op_i == fpnew_pkg::CPKCD), op_mod_i};
  assign is_up_cast   = (fpnew_pkg::fp_width(dst_fmt_i) > fpnew_pkg::fp_width(src_fmt_i));
  assign is_down_cast = (fpnew_pkg::fp_width(dst_fmt_i) < fpnew_pkg::fp_width(src_fmt_i));
  
  assign dst_fmt    = dst_fmt_is_int ? int_fmt_i : dst_fmt_i;
  
  assign aux_data      = {dst_fmt_is_int, vectorial_op, dst_fmt};
  assign target_aux_d  = {dst_vec_op, dst_is_cpk};
  
  if (OpGroup == fpnew_pkg::CONV) begin : conv_target
    assign conv_target_d = dst_is_cpk ? operands_i[2] : operands_i[1];
  end
  
  logic [NUM_FORMATS-1:0]      is_boxed_1op;
  logic [NUM_FORMATS-1:0][1:0] is_boxed_2op;
  always_comb begin : boxed_2op
    for (int fmt = 0; fmt < NUM_FORMATS; fmt++) begin
      is_boxed_1op[fmt] = is_boxed_i[fmt][0];
      is_boxed_2op[fmt] = is_boxed_i[fmt][1:0];
    end
  end
  
  
  
  for (genvar lane = 0; lane < int'(NUM_LANES); lane++) begin : gen_num_lanes
    localparam int unsigned LANE = unsigned'(lane); 
    
    localparam fpnew_pkg::fmt_logic_t ACTIVE_FORMATS =
        fpnew_pkg::get_lane_formats(Width, FpFmtConfig, LANE);
    localparam fpnew_pkg::ifmt_logic_t ACTIVE_INT_FORMATS =
        fpnew_pkg::get_lane_int_formats(Width, FpFmtConfig, IntFmtConfig, LANE);
    localparam int unsigned MAX_WIDTH = fpnew_pkg::max_fp_width(ACTIVE_FORMATS);
    
    localparam fpnew_pkg::fmt_logic_t CONV_FORMATS =
        fpnew_pkg::get_conv_lane_formats(Width, FpFmtConfig, LANE);
    localparam fpnew_pkg::ifmt_logic_t CONV_INT_FORMATS =
        fpnew_pkg::get_conv_lane_int_formats(Width, FpFmtConfig, IntFmtConfig, LANE);
    localparam int unsigned CONV_WIDTH = fpnew_pkg::max_fp_width(CONV_FORMATS);
    
    localparam fpnew_pkg::fmt_logic_t LANE_FORMATS = (OpGroup == fpnew_pkg::CONV)
                                                     ? CONV_FORMATS : ACTIVE_FORMATS;
    localparam int unsigned LANE_WIDTH = (OpGroup == fpnew_pkg::CONV) ? CONV_WIDTH : MAX_WIDTH;
    logic [LANE_WIDTH-1:0] local_result; 
    
    if ((lane == 0) || EnableVectors) begin : active_lane
      logic in_valid, out_valid, out_ready; 
      logic [NUM_OPERANDS-1:0][LANE_WIDTH-1:0] local_operands;  
      logic [LANE_WIDTH-1:0]                   op_result;       
      fpnew_pkg::status_t                      op_status;
      assign in_valid = in_valid_i & ((lane == 0) | vectorial_op); 
      
      always_comb begin : prepare_input
        for (int unsigned i = 0; i < NUM_OPERANDS; i++) begin
          local_operands[i] = operands_i[i] >> LANE*fpnew_pkg::fp_width(src_fmt_i);
        end
        
        if (OpGroup == fpnew_pkg::CONV) begin
          
          if (op_i == fpnew_pkg::I2F) begin
            local_operands[0] = operands_i[0] >> LANE*fpnew_pkg::int_width(int_fmt_i);
          
          end else if (op_i == fpnew_pkg::F2F) begin
            if (vectorial_op && op_mod_i && is_up_cast) begin 
              local_operands[0] = operands_i[0] >> LANE*fpnew_pkg::fp_width(src_fmt_i) +
                                                   MAX_FP_WIDTH/2;
            end
          
          end else if (dst_is_cpk) begin
            if (lane == 1) begin
              local_operands[0] = operands_i[1][LANE_WIDTH-1:0]; 
            end
          end
        end
      end
      
      if (OpGroup == fpnew_pkg::ADDMUL) begin : lane_instance
        fpnew_fma_multi #(
          .FpFmtConfig ( LANE_FORMATS         ),
          .NumPipeRegs ( NumPipeRegs          ),
          .PipeConfig  ( PipeConfig           ),
          .TagType     ( TagType              ),
          .AuxType     ( logic [AUX_BITS-1:0] )
        ) i_fpnew_fma_multi (
          .clk_i,
          .rst_ni,
          .operands_i      ( local_operands  ),
          .is_boxed_i,
          .rnd_mode_i,
          .op_i,
          .op_mod_i,
          .src_fmt_i,
          .dst_fmt_i,
          .tag_i,
          .aux_i           ( aux_data            ),
          .in_valid_i      ( in_valid            ),
          .in_ready_o      ( lane_in_ready[lane] ),
          .flush_i,
          .result_o        ( op_result           ),
          .status_o        ( op_status           ),
          .extension_bit_o ( lane_ext_bit[lane]  ),
          .tag_o           ( lane_tags[lane]     ),
          .aux_o           ( lane_aux[lane]      ),
          .out_valid_o     ( out_valid           ),
          .out_ready_i     ( out_ready           ),
          .busy_o          ( lane_busy[lane]     )
        );
      end else if (OpGroup == fpnew_pkg::DIVSQRT) begin : lane_instance
        fpnew_divsqrt_multi #(
          .FpFmtConfig ( LANE_FORMATS         ),
          .NumPipeRegs ( NumPipeRegs          ),
          .PipeConfig  ( PipeConfig           ),
          .TagType     ( TagType              ),
          .AuxType     ( logic [AUX_BITS-1:0] )
        ) i_fpnew_divsqrt_multi (
          .clk_i,
          .rst_ni,
          .operands_i      ( local_operands[1:0] ), 
          .is_boxed_i      ( is_boxed_2op        ), 
          .rnd_mode_i,
          .op_i,
          .dst_fmt_i,
          .tag_i,
          .aux_i           ( aux_data            ),
          .in_valid_i      ( in_valid            ),
          .in_ready_o      ( lane_in_ready[lane] ),
          .flush_i,
          .result_o        ( op_result           ),
          .status_o        ( op_status           ),
          .extension_bit_o ( lane_ext_bit[lane]  ),
          .tag_o           ( lane_tags[lane]     ),
          .aux_o           ( lane_aux[lane]      ),
          .out_valid_o     ( out_valid           ),
          .out_ready_i     ( out_ready           ),
          .busy_o          ( lane_busy[lane]     )
        );
      end else if (OpGroup == fpnew_pkg::NONCOMP) begin : lane_instance
      end else if (OpGroup == fpnew_pkg::CONV) begin : lane_instance
        fpnew_cast_multi #(
          .FpFmtConfig  ( LANE_FORMATS         ),
          .IntFmtConfig ( CONV_INT_FORMATS     ),
          .NumPipeRegs  ( NumPipeRegs          ),
          .PipeConfig   ( PipeConfig           ),
          .TagType      ( TagType              ),
          .AuxType      ( logic [AUX_BITS-1:0] )
        ) i_fpnew_cast_multi (
          .clk_i,
          .rst_ni,
          .operands_i      ( local_operands[0]   ),
          .is_boxed_i      ( is_boxed_1op        ),
          .rnd_mode_i,
          .op_i,
          .op_mod_i,
          .src_fmt_i,
          .dst_fmt_i,
          .int_fmt_i,
          .tag_i,
          .aux_i           ( aux_data            ),
          .in_valid_i      ( in_valid            ),
          .in_ready_o      ( lane_in_ready[lane] ),
          .flush_i,
          .result_o        ( op_result           ),
          .status_o        ( op_status           ),
          .extension_bit_o ( lane_ext_bit[lane]  ),
          .tag_o           ( lane_tags[lane]     ),
          .aux_o           ( lane_aux[lane]      ),
          .out_valid_o     ( out_valid           ),
          .out_ready_i     ( out_ready           ),
          .busy_o          ( lane_busy[lane]     )
        );
      end 
      
      assign out_ready            = out_ready_i & ((lane == 0) | result_is_vector);
      assign lane_out_valid[lane] = out_valid & ((lane == 0) | result_is_vector);
      
      assign local_result      = lane_out_valid[lane] ? op_result : '{default: lane_ext_bit[0]};
      assign lane_status[lane] = lane_out_valid[lane] ? op_status : '0;
    
    end else begin : inactive_lane
      assign lane_out_valid[lane] = 1'b0; 
      assign lane_in_ready[lane]  = 1'b0; 
      assign local_result         = '{default: lane_ext_bit[0]}; 
      assign lane_status[lane]    = '0;
      assign lane_busy[lane]      = 1'b0;
    end
    
    for (genvar fmt = 0; fmt < NUM_FORMATS; fmt++) begin : pack_fp_result
      
      localparam int unsigned FP_WIDTH = fpnew_pkg::fp_width(fpnew_pkg::fp_format_e'(fmt));
      
      if (ACTIVE_FORMATS[fmt])
        assign fmt_slice_result[fmt][(LANE+1)*FP_WIDTH-1:LANE*FP_WIDTH] =
            local_result[FP_WIDTH-1:0];
    end
    
    if (OpGroup == fpnew_pkg::CONV) begin : int_results_enabled
      for (genvar ifmt = 0; ifmt < NUM_INT_FORMATS; ifmt++) begin : pack_int_result
        
        localparam int unsigned INT_WIDTH = fpnew_pkg::int_width(fpnew_pkg::int_format_e'(ifmt));
        if (ACTIVE_INT_FORMATS[ifmt])
          assign ifmt_slice_result[ifmt][(LANE+1)*INT_WIDTH-1:LANE*INT_WIDTH] =
            local_result[INT_WIDTH-1:0];
      end
    end
  end
  
  for (genvar fmt = 0; fmt < NUM_FORMATS; fmt++) begin : extend_fp_result
    
    localparam int unsigned FP_WIDTH = fpnew_pkg::fp_width(fpnew_pkg::fp_format_e'(fmt));
    if (NUM_LANES*FP_WIDTH < Width)
      assign fmt_slice_result[fmt][Width-1:NUM_LANES*FP_WIDTH] = '{default: lane_ext_bit[0]};
  end
  
  for (genvar ifmt = 0; ifmt < NUM_INT_FORMATS; ifmt++) begin : int_results_disabled
    if (OpGroup != fpnew_pkg::CONV) begin : mute_int_result
      assign ifmt_slice_result[ifmt] = '0;
    end
  end
  
  if (OpGroup == fpnew_pkg::CONV) begin : target_regs
    
    logic [0:NumPipeRegs][Width-1:0] byp_pipe_target_q;
    logic [0:NumPipeRegs][2:0]       byp_pipe_aux_q;
    logic [0:NumPipeRegs]            byp_pipe_valid_q;
    
    logic [0:NumPipeRegs] byp_pipe_ready;
    
    assign byp_pipe_target_q[0]  = conv_target_d;
    assign byp_pipe_aux_q[0]     = target_aux_d;
    assign byp_pipe_valid_q[0]   = in_valid_i & vectorial_op;
    
    for (genvar i = 0; i < NumPipeRegs; i++) begin : gen_bypass_pipeline
      
      logic reg_ena;
      
      
      
      assign byp_pipe_ready[i] = byp_pipe_ready[i+1] | ~byp_pipe_valid_q[i+1];
      
      
                           
                         
                            
  always_ff @(posedge (clk_i) or negedge (rst_ni)) begin                 
    if (!rst_ni) begin                                                   
      byp_pipe_valid_q[i+1] <= (1'b0);                                              
    end else begin                                                         
      byp_pipe_valid_q[i+1] <= (flush_i) ? (1'b0) : (byp_pipe_ready[i]) ? (byp_pipe_valid_q[i]) : (byp_pipe_valid_q[i+1]);       
    end                                                                    
  end
      
      assign reg_ena = byp_pipe_ready[i] & byp_pipe_valid_q[i];
      
      
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      byp_pipe_target_q[i+1] <= ('0);                        
    end else begin                                   
      byp_pipe_target_q[i+1] <= (reg_ena) ? (byp_pipe_target_q[i]) : (byp_pipe_target_q[i+1]);               
    end                                              
  end
      
  always_ff @(posedge clk_i or negedge rst_ni) begin 
    if (!rst_ni) begin                               
      byp_pipe_aux_q[i+1] <= ('0);                        
    end else begin                                   
      byp_pipe_aux_q[i+1] <= (reg_ena) ? (byp_pipe_aux_q[i]) : (byp_pipe_aux_q[i+1]);               
    end                                              
  end
    end
    
    assign byp_pipe_ready[NumPipeRegs] = out_ready_i & result_is_vector;
    
    assign conv_target_q = byp_pipe_target_q[NumPipeRegs];
    
    assign {result_vec_op, result_is_cpk} = byp_pipe_aux_q[NumPipeRegs];
  end else begin : no_conv
    assign {result_vec_op, result_is_cpk} = '0;
  end
  
  
  
  assign {result_fmt_is_int, result_is_vector, result_fmt} = lane_aux[0];
  assign result_o = result_fmt_is_int
                    ? ifmt_slice_result[result_fmt]
                    : fmt_slice_result[result_fmt];
  assign extension_bit_o = lane_ext_bit[0]; 
  assign tag_o           = lane_tags[0];    
  assign busy_o          = (| lane_busy);
  assign out_valid_o     = lane_out_valid[0]; 
  
  always_comb begin : output_processing
    
    automatic fpnew_pkg::status_t temp_status;
    temp_status = '0;
    for (int i = 0; i < int'(NUM_LANES); i++)
      temp_status |= lane_status[i];
    status_o = temp_status;
  end
endmodule
module fpnew_rounding #(
  parameter int unsigned AbsWidth=2 
) (
  
  input logic [AbsWidth-1:0]   abs_value_i,             
  input logic                  sign_i,
  
  input logic [1:0]            round_sticky_bits_i,     
  input fpnew_pkg::roundmode_e rnd_mode_i,
  input logic                  effective_subtraction_i, 
  
  output logic [AbsWidth-1:0]  abs_rounded_o,           
  output logic                 sign_o,
  
  output logic                 exact_zero_o             
);
  logic round_up; 
  
  
  
  
  
  
  
  
  
  always_comb begin : rounding_decision
    unique case (rnd_mode_i)
      fpnew_pkg::RNE: 
        unique case (round_sticky_bits_i)
          2'b00,
          2'b01: round_up = 1'b0;           
          2'b10: round_up = abs_value_i[0]; 
          2'b11: round_up = 1'b1;           
          default: round_up = fpnew_pkg::DONT_CARE;
        endcase
      fpnew_pkg::RTZ: round_up = 1'b0; 
      fpnew_pkg::RDN: round_up = (| round_sticky_bits_i) ? sign_i  : 1'b0; 
      fpnew_pkg::RUP: round_up = (| round_sticky_bits_i) ? ~sign_i : 1'b0; 
      fpnew_pkg::RMM: round_up = round_sticky_bits_i[1]; 
      default: round_up = fpnew_pkg::DONT_CARE; 
    endcase
  end
  
  assign abs_rounded_o = abs_value_i + round_up;
  
  assign exact_zero_o = (abs_value_i == '0) && (round_sticky_bits_i == '0);
  
  
  assign sign_o = (exact_zero_o && effective_subtraction_i)
                  ? (rnd_mode_i == fpnew_pkg::RDN)
                  : sign_i;
endmodule
module fpnew_top #(
  
  parameter fpnew_pkg::fpu_features_t       Features       = fpnew_pkg::RV64D_Xsflt,
  parameter fpnew_pkg::fpu_implementation_t Implementation = fpnew_pkg::DEFAULT_NOREGS,
  parameter type                            TagType        = logic,
  
  localparam int unsigned WIDTH        = Features.Width,
  localparam int unsigned NUM_OPERANDS = 3
) (
  input logic                               clk_i,
  input logic                               rst_ni,
  
  input logic [NUM_OPERANDS-1:0][WIDTH-1:0] operands_i,
  input fpnew_pkg::roundmode_e              rnd_mode_i,
  input fpnew_pkg::operation_e              op_i,
  input logic                               op_mod_i,
  input fpnew_pkg::fp_format_e              src_fmt_i,
  input fpnew_pkg::fp_format_e              dst_fmt_i,
  input fpnew_pkg::int_format_e             int_fmt_i,
  input logic                               vectorial_op_i,
  input TagType                             tag_i,
  
  input  logic                              in_valid_i,
  output logic                              in_ready_o,
  input  logic                              flush_i,
  
  output logic [WIDTH-1:0]                  result_o,
  output fpnew_pkg::status_t                status_o,
  output TagType                            tag_o,
  
  output logic                              out_valid_o,
  input  logic                              out_ready_i,
  
  output logic                              busy_o
);
  localparam int unsigned NUM_OPGROUPS = fpnew_pkg::NUM_OPGROUPS;
  localparam int unsigned NUM_FORMATS  = fpnew_pkg::NUM_FP_FORMATS;
  
  
  
  typedef struct packed {
    logic [WIDTH-1:0]   result;
    fpnew_pkg::status_t status;
    TagType             tag;
  } output_t;
  
  logic [NUM_OPGROUPS-1:0] opgrp_in_ready, opgrp_out_valid, opgrp_out_ready, opgrp_ext, opgrp_busy;
  output_t [NUM_OPGROUPS-1:0] opgrp_outputs;
  logic [NUM_FORMATS-1:0][NUM_OPERANDS-1:0] is_boxed;
  
  
  
  assign in_ready_o = in_valid_i & opgrp_in_ready[fpnew_pkg::get_opgroup(op_i)];
  
  for (genvar fmt = 0; fmt < int'(NUM_FORMATS); fmt++) begin : gen_nanbox_check
    localparam int unsigned FP_WIDTH = fpnew_pkg::fp_width(fpnew_pkg::fp_format_e'(fmt));
    
    if (Features.EnableNanBox && (FP_WIDTH < WIDTH)) begin : check
      for (genvar op = 0; op < int'(NUM_OPERANDS); op++) begin : operands
        assign is_boxed[fmt][op] = (!vectorial_op_i)
                                   ? operands_i[op][WIDTH-1:FP_WIDTH] == '1
                                   : 1'b1;
      end
    end else begin : no_check
      assign is_boxed[fmt] = '1;
    end
  end
  
  
  
  for (genvar opgrp = 0; opgrp < int'(NUM_OPGROUPS); opgrp++) begin : gen_operation_groups
    localparam int unsigned NUM_OPS = fpnew_pkg::num_operands(fpnew_pkg::opgroup_e'(opgrp));
    logic in_valid;
    logic [NUM_FORMATS-1:0][NUM_OPS-1:0] input_boxed;
    assign in_valid = in_valid_i & (fpnew_pkg::get_opgroup(op_i) == fpnew_pkg::opgroup_e'(opgrp));
    
    always_comb begin : slice_inputs
      for (int unsigned fmt = 0; fmt < NUM_FORMATS; fmt++)
        input_boxed[fmt] = is_boxed[fmt][NUM_OPS-1:0];
    end
    fpnew_opgroup_block #(
      .OpGroup       ( fpnew_pkg::opgroup_e'(opgrp)    ),
      .Width         ( WIDTH                           ),
      .EnableVectors ( Features.EnableVectors          ),
      .FpFmtMask     ( Features.FpFmtMask              ),
      .IntFmtMask    ( Features.IntFmtMask             ),
      .FmtPipeRegs   ( Implementation.PipeRegs[opgrp]  ),
      .FmtUnitTypes  ( Implementation.UnitTypes[opgrp] ),
      .PipeConfig    ( Implementation.PipeConfig       ),
      .TagType       ( TagType                         )
    ) i_opgroup_block (
      .clk_i,
      .rst_ni,
      .operands_i      ( operands_i[NUM_OPS-1:0] ),
      .is_boxed_i      ( input_boxed             ),
      .rnd_mode_i,
      .op_i,
      .op_mod_i,
      .src_fmt_i,
      .dst_fmt_i,
      .int_fmt_i,
      .vectorial_op_i,
      .tag_i,
      .in_valid_i      ( in_valid              ),
      .in_ready_o      ( opgrp_in_ready[opgrp] ),
      .flush_i,
      .result_o        ( opgrp_outputs[opgrp].result ),
      .status_o        ( opgrp_outputs[opgrp].status ),
      .extension_bit_o ( opgrp_ext[opgrp]            ),
      .tag_o           ( opgrp_outputs[opgrp].tag    ),
      .out_valid_o     ( opgrp_out_valid[opgrp]      ),
      .out_ready_i     ( opgrp_out_ready[opgrp]      ),
      .busy_o          ( opgrp_busy[opgrp]           )
    );
  end
  
  
  
  output_t arbiter_output;
  
  rr_arb_tree #(
    .NumIn     ( NUM_OPGROUPS ),
    .DataType  ( output_t     ),
    .AxiVldRdy ( 1'b1         )
  ) i_arbiter (
    .clk_i,
    .rst_ni,
    .flush_i,
    .rr_i   ( '0             ),
    .req_i  ( opgrp_out_valid ),
    .gnt_o  ( opgrp_out_ready ),
    .data_i ( opgrp_outputs   ),
    .gnt_i  ( out_ready_i     ),
    .req_o  ( out_valid_o     ),
    .data_o ( arbiter_output  ),
    .idx_o  (     )
  );
  
  assign result_o        = arbiter_output.result;
  assign status_o        = arbiter_output.status;
  assign tag_o           = arbiter_output.tag;
  assign busy_o = (| opgrp_busy);
endmodule
package axi_pkg;
  typedef logic [1:0] burst_t;
  typedef logic [1:0] resp_t;
  typedef logic [3:0] cache_t;
  typedef logic [2:0] prot_t;
  typedef logic [3:0] qos_t;
  typedef logic [3:0] region_t;
  typedef logic [7:0] len_t;
  typedef logic [2:0] size_t;
  typedef logic [5:0] atop_t; 
  typedef logic [3:0] nsaid_t; 
  localparam BURST_FIXED = 2'b00;
  localparam BURST_INCR  = 2'b01;
  localparam BURST_WRAP  = 2'b10;
  localparam RESP_OKAY   = 2'b00;
  localparam RESP_EXOKAY = 2'b01;
  localparam RESP_SLVERR = 2'b10;
  localparam RESP_DECERR = 2'b11;
  localparam CACHE_BUFFERABLE = 4'b0001;
  localparam CACHE_MODIFIABLE = 4'b0010;
  localparam CACHE_RD_ALLOC   = 4'b0100;
  localparam CACHE_WR_ALLOC   = 4'b1000;
  
  localparam ATOP_ATOMICSWAP  = 6'b110000;
  localparam ATOP_ATOMICCMP   = 6'b110001;
  
  localparam ATOP_NONE        = 2'b00;
  localparam ATOP_ATOMICSTORE = 2'b01;
  localparam ATOP_ATOMICLOAD  = 2'b10;
  
  localparam ATOP_LITTLE_END  = 1'b0;
  localparam ATOP_BIG_END     = 1'b1;
  
  localparam ATOP_ADD   = 3'b000;
  localparam ATOP_CLR   = 3'b001;
  localparam ATOP_EOR   = 3'b010;
  localparam ATOP_SET   = 3'b011;
  localparam ATOP_SMAX  = 3'b100;
  localparam ATOP_SMIN  = 3'b101;
  localparam ATOP_UMAX  = 3'b110;
  localparam ATOP_UMIN  = 3'b111;
  
  localparam IdWidth   = 4;
  localparam UserWidth = 1;
  localparam AddrWidth = 64;
  localparam DataWidth = 64;
  localparam StrbWidth = DataWidth / 8;
  typedef logic [IdWidth-1:0]   id_t;
  typedef logic [AddrWidth-1:0] addr_t;
  typedef logic [DataWidth-1:0] data_t;
  typedef logic [StrbWidth-1:0] strb_t;
  typedef logic [UserWidth-1:0] user_t;
  
  typedef struct packed {
      id_t     id;
      addr_t   addr;
      len_t    len;
      size_t   size;
      burst_t  burst;
      logic   lock;
      cache_t  cache;
      prot_t   prot;
      qos_t    qos;
      region_t region;
      atop_t   atop;
  } aw_chan_t;
  
  typedef struct packed {
      data_t data;
      strb_t strb;
      logic  last;
  } w_chan_t;
  
  typedef struct packed {
      id_t   id;
      resp_t resp;
  } b_chan_t;
  
  typedef struct packed {
      id_t     id;
      addr_t   addr;
      len_t    len;
      size_t   size;
      burst_t  burst;
      logic    lock;
      cache_t  cache;
      prot_t   prot;
      qos_t    qos;
      region_t region;
  } ar_chan_t;
  
  typedef struct packed {
      id_t   id;
      data_t data;
      resp_t resp;
      logic  last;
  } r_chan_t;
endpackage
package ariane_soc;
  
  localparam int unsigned NumTargets = 2;
  
  localparam int unsigned NumSources = 30;
  localparam int unsigned MaxPriority = 7;
  localparam NrSlaves = 2; 
  
  localparam IdWidth   = 4;
  localparam IdWidthSlave = IdWidth + $clog2(NrSlaves);
  typedef enum int unsigned {
    DRAM     = 0,
    GPIO     = 1,
    Ethernet = 2,
    SPI      = 3,
    Timer    = 4,
    UART     = 5,
    PLIC     = 6,
    CLINT    = 7,
    ROM      = 8,
    Debug    = 9
  } axi_slaves_t;
  localparam NB_PERIPHERALS = Debug + 1;
  localparam logic[63:0] DebugLength    = 64'h1000;
  localparam logic[63:0] ROMLength      = 64'h10000;
  localparam logic[63:0] CLINTLength    = 64'hC0000;
  localparam logic[63:0] PLICLength     = 64'h3FF_FFFF;
  localparam logic[63:0] UARTLength     = 64'h1000;
  localparam logic[63:0] TimerLength    = 64'h1000;
  localparam logic[63:0] SPILength      = 64'h800000;
  localparam logic[63:0] EthernetLength = 64'h10000;
  localparam logic[63:0] GPIOLength     = 64'h1000;
  localparam logic[63:0] DRAMLength     = 64'h40000000; 
  localparam logic[63:0] SRAMLength     = 64'h1800000;  
  
  localparam bit GenProtocolChecker = 1'b0;
  typedef enum logic [63:0] {
    DebugBase    = 64'h0000_0000,
    ROMBase      = 64'h0001_0000,
    CLINTBase    = 64'h0200_0000,
    PLICBase     = 64'h0C00_0000,
    UARTBase     = 64'h1000_0000,
    TimerBase    = 64'h1800_0000,
    SPIBase      = 64'h2000_0000,
    EthernetBase = 64'h3000_0000,
    GPIOBase     = 64'h4000_0000,
    DRAMBase     = 64'h8000_0000
  } soc_bus_start_t;
  localparam NrRegion = 1;
  localparam logic [NrRegion-1:0][NB_PERIPHERALS-1:0] ValidRule = {{NrRegion * NB_PERIPHERALS}{1'b1}};
  localparam ariane_pkg::ariane_cfg_t ArianeSocCfg = '{
    RASDepth: 2,
    BTBEntries: 32,
    BHTEntries: 128,
    
    NrNonIdempotentRules:  1,
    NonIdempotentAddrBase: {64'b0},
    NonIdempotentLength:   {DRAMBase},
    NrExecuteRegionRules:  3,
    ExecuteRegionAddrBase: {DRAMBase,   ROMBase,   DebugBase},
    ExecuteRegionLength:   {DRAMLength, ROMLength, DebugLength},
    
    NrCachedRegionRules:    1,
    CachedRegionAddrBase:  {DRAMBase},
    CachedRegionLength:    {DRAMLength},
    
    Axi64BitCompliant:      1'b1,
    SwapEndianess:          1'b0,
    
    DmBaseAddress:          DebugBase,
    NrPMPEntries:           8
  };
endpackage
package ariane_axi_soc;
    
    typedef enum logic { SINGLE_REQ, CACHE_LINE_REQ } ad_req_t;
    localparam UserWidth = 1;
    localparam AddrWidth = 64;
    localparam DataWidth = 64;
    localparam StrbWidth = DataWidth / 8;
    typedef logic [ariane_soc::IdWidth-1:0]      id_t;
    typedef logic [ariane_soc::IdWidthSlave-1:0] id_slv_t;
    typedef logic [AddrWidth-1:0] addr_t;
    typedef logic [DataWidth-1:0] data_t;
    typedef logic [StrbWidth-1:0] strb_t;
    typedef logic [UserWidth-1:0] user_t;
    
    typedef struct packed {
        id_t              id;
        addr_t            addr;
        axi_pkg::len_t    len;
        axi_pkg::size_t   size;
        axi_pkg::burst_t  burst;
        logic             lock;
        axi_pkg::cache_t  cache;
        axi_pkg::prot_t   prot;
        axi_pkg::qos_t    qos;
        axi_pkg::region_t region;
        axi_pkg::atop_t   atop;
        user_t            user;
    } aw_chan_t;
    
    typedef struct packed {
        id_slv_t          id;
        addr_t            addr;
        axi_pkg::len_t    len;
        axi_pkg::size_t   size;
        axi_pkg::burst_t  burst;
        logic             lock;
        axi_pkg::cache_t  cache;
        axi_pkg::prot_t   prot;
        axi_pkg::qos_t    qos;
        axi_pkg::region_t region;
        axi_pkg::atop_t   atop;
        user_t            user;
    } aw_chan_slv_t;
    
    typedef struct packed {
        data_t data;
        strb_t strb;
        logic  last;
        user_t user;
    } w_chan_t;
    
    typedef struct packed {
        id_t            id;
        axi_pkg::resp_t resp;
        user_t          user;
    } b_chan_t;
    
    typedef struct packed {
        id_slv_t        id;
        axi_pkg::resp_t resp;
        user_t          user;
    } b_chan_slv_t;
    
    typedef struct packed {
        id_t             id;
        addr_t            addr;
        axi_pkg::len_t    len;
        axi_pkg::size_t   size;
        axi_pkg::burst_t  burst;
        logic             lock;
        axi_pkg::cache_t  cache;
        axi_pkg::prot_t   prot;
        axi_pkg::qos_t    qos;
        axi_pkg::region_t region;
        user_t            user;
    } ar_chan_t;
    
    typedef struct packed {
        id_slv_t          id;
        addr_t            addr;
        axi_pkg::len_t    len;
        axi_pkg::size_t   size;
        axi_pkg::burst_t  burst;
        logic             lock;
        axi_pkg::cache_t  cache;
        axi_pkg::prot_t   prot;
        axi_pkg::qos_t    qos;
        axi_pkg::region_t region;
        user_t            user;
    } ar_chan_slv_t;
    
    typedef struct packed {
        id_t            id;
        data_t          data;
        axi_pkg::resp_t resp;
        logic           last;
        user_t          user;
    } r_chan_t;
    
    typedef struct packed {
        id_slv_t        id;
        data_t          data;
        axi_pkg::resp_t resp;
        logic           last;
        user_t          user;
    } r_chan_slv_t;
    
    typedef struct packed {
        aw_chan_t aw;
        logic     aw_valid;
        w_chan_t  w;
        logic     w_valid;
        logic     b_ready;
        ar_chan_t ar;
        logic     ar_valid;
        logic     r_ready;
    } req_t;
    typedef struct packed {
        logic     aw_ready;
        logic     ar_ready;
        logic     w_ready;
        logic     b_valid;
        b_chan_t  b;
        logic     r_valid;
        r_chan_t  r;
    } resp_t;
    typedef struct packed {
        aw_chan_slv_t aw;
        logic         aw_valid;
        w_chan_t      w;
        logic         w_valid;
        logic         b_ready;
        ar_chan_slv_t ar;
        logic         ar_valid;
        logic         r_ready;
    } req_slv_t;
    typedef struct packed {
        logic         aw_ready;
        logic         ar_ready;
        logic         w_ready;
        logic         b_valid;
        b_chan_slv_t  b;
        logic         r_valid;
        r_chan_slv_t  r;
    } resp_slv_t;
endpackage
package ariane_axi;
    
    typedef enum logic { SINGLE_REQ, CACHE_LINE_REQ } ad_req_t;
    localparam IdWidth   = 4; 
    localparam UserWidth = 1;
    localparam AddrWidth = 64;
    localparam DataWidth = 64;
    localparam StrbWidth = DataWidth / 8;
    typedef logic   [IdWidth-1:0]   id_t;
    typedef logic [AddrWidth-1:0] addr_t;
    typedef logic [DataWidth-1:0] data_t;
    typedef logic [StrbWidth-1:0] strb_t;
    typedef logic [UserWidth-1:0] user_t;
    
    typedef struct packed {
        id_t              id;
        addr_t            addr;
        axi_pkg::len_t    len;
        axi_pkg::size_t   size;
        axi_pkg::burst_t  burst;
        logic             lock;
        axi_pkg::cache_t  cache;
        axi_pkg::prot_t   prot;
        axi_pkg::qos_t    qos;
        axi_pkg::region_t region;
        axi_pkg::atop_t   atop;
        user_t            user;
    } aw_chan_t;
    
    typedef struct packed {
        data_t data;
        strb_t strb;
        logic  last;
        user_t user;
    } w_chan_t;
    
    typedef struct packed {
        id_t            id;
        axi_pkg::resp_t resp;
        user_t          user;
    } b_chan_t;
    
    typedef struct packed {
        id_t             id;
        addr_t            addr;
        axi_pkg::len_t    len;
        axi_pkg::size_t   size;
        axi_pkg::burst_t  burst;
        logic             lock;
        axi_pkg::cache_t  cache;
        axi_pkg::prot_t   prot;
        axi_pkg::qos_t    qos;
        axi_pkg::region_t region;
        user_t            user;
    } ar_chan_t;
    
    typedef struct packed {
        id_t            id;
        data_t          data;
        axi_pkg::resp_t resp;
        logic           last;
        user_t          user;
    } r_chan_t;
    
    typedef struct packed {
        aw_chan_t aw;
        logic     aw_valid;
        w_chan_t  w;
        logic     w_valid;
        logic     b_ready;
        ar_chan_t ar;
        logic     ar_valid;
        logic     r_ready;
    } req_t;
    typedef struct packed {
        logic     aw_ready;
        logic     ar_ready;
        logic     w_ready;
        logic     b_valid;
        b_chan_t  b;
        logic     r_valid;
        r_chan_t  r;
    } resp_t;
endpackage
  
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
  
package wt_cache_pkg;
  
  
  localparam L15_SET_ASSOC           = 4;
  localparam L15_TID_WIDTH           = 1;
  localparam L15_TLB_CSM_WIDTH       = 33;
  localparam L15_WAY_WIDTH           = $clog2(L15_SET_ASSOC);
  localparam L1I_WAY_WIDTH           = $clog2(ariane_pkg::ICACHE_SET_ASSOC);
  localparam L1D_WAY_WIDTH           = $clog2(ariane_pkg::DCACHE_SET_ASSOC);
  
  localparam ADAPTER_REQ_FIFO_DEPTH  = 2;
  localparam ADAPTER_RTRN_FIFO_DEPTH = 2;
  
  localparam ICACHE_OFFSET_WIDTH     = $clog2(ariane_pkg::ICACHE_LINE_WIDTH/8);
  localparam ICACHE_NUM_WORDS        = 2**(ariane_pkg::ICACHE_INDEX_WIDTH-ICACHE_OFFSET_WIDTH);
  localparam ICACHE_CL_IDX_WIDTH     = $clog2(ICACHE_NUM_WORDS);
  localparam DCACHE_OFFSET_WIDTH     = $clog2(ariane_pkg::DCACHE_LINE_WIDTH/8);
  localparam DCACHE_NUM_WORDS        = 2**(ariane_pkg::DCACHE_INDEX_WIDTH-DCACHE_OFFSET_WIDTH);
  localparam DCACHE_CL_IDX_WIDTH     = $clog2(DCACHE_NUM_WORDS);
  localparam DCACHE_NUM_BANKS        = ariane_pkg::DCACHE_LINE_WIDTH/64;
  localparam DCACHE_NUM_BANKS_WIDTH  = $clog2(DCACHE_NUM_BANKS);
  
  localparam DCACHE_WBUF_DEPTH       = 8;
  localparam DCACHE_MAX_TX           = 2**L15_TID_WIDTH;
  localparam CACHE_ID_WIDTH          = L15_TID_WIDTH;
  typedef struct packed {
    logic [ariane_pkg::DCACHE_INDEX_WIDTH+ariane_pkg::DCACHE_TAG_WIDTH-1:0] wtag;
    logic [63:0]                                                            data;
    logic [7:0]                                                             dirty;   
    logic [7:0]                                                             valid;   
    logic [7:0]                                                             txblock; 
    logic                                                                   checked; 
    logic [ariane_pkg::DCACHE_SET_ASSOC-1:0]                                hit_oh;  
  } wbuffer_t;
  
  
  
  typedef struct packed {
    logic                                 vld;
    logic [7:0]                           be;
    logic [$clog2(DCACHE_WBUF_DEPTH)-1:0] ptr;
  } tx_stat_t;
  
  typedef enum logic [1:0] {
    DCACHE_STORE_REQ,
    DCACHE_LOAD_REQ,
    DCACHE_ATOMIC_REQ,
    DCACHE_INT_REQ
  }  dcache_out_t;
  typedef enum logic [2:0] {
    DCACHE_INV_REQ,  
    DCACHE_STORE_ACK,
    DCACHE_LOAD_ACK,
    DCACHE_ATOMIC_ACK,
    DCACHE_INT_ACK
  }  dcache_in_t;
  typedef enum logic [0:0] {
    ICACHE_INV_REQ, 
    ICACHE_IFILL_ACK
  } icache_in_t;
  
  typedef struct packed {
    logic                                            vld;         
    logic                                            all;         
    logic [ariane_pkg::ICACHE_INDEX_WIDTH-1:0]       idx;         
    logic [L15_WAY_WIDTH-1:0]                        way;         
  } icache_inval_t;
  typedef struct packed {
    logic [$clog2(ariane_pkg::ICACHE_SET_ASSOC)-1:0] way;         
    logic [riscv::PLEN-1:0]                          paddr;       
    logic                                            nc;          
    logic [CACHE_ID_WIDTH-1:0]                       tid;         
  } icache_req_t;
  typedef struct packed {
    icache_in_t                                      rtype;       
    logic [ariane_pkg::ICACHE_LINE_WIDTH-1:0]        data;        
    icache_inval_t                                   inv;         
    logic [CACHE_ID_WIDTH-1:0]                       tid;         
  } icache_rtrn_t;
  
  typedef struct packed {
    logic                                            vld;         
    logic                                            all;         
    logic [ariane_pkg::DCACHE_INDEX_WIDTH-1:0]       idx;         
    logic [L15_WAY_WIDTH-1:0]                        way;         
  } dcache_inval_t;
  typedef struct packed {
    dcache_out_t                                     rtype;       
    logic [2:0]                                      size;        
    logic [L1D_WAY_WIDTH-1:0]                        way;         
    logic [riscv::PLEN-1:0]                          paddr;       
    logic [63:0]                                     data;        
    logic                                            nc;          
    logic [CACHE_ID_WIDTH-1:0]                       tid;         
    ariane_pkg::amo_t                                amo_op;      
  } dcache_req_t;
  typedef struct packed {
    dcache_in_t                                      rtype;       
    logic [ariane_pkg::DCACHE_LINE_WIDTH-1:0]        data;        
    dcache_inval_t                                   inv;         
    logic [CACHE_ID_WIDTH-1:0]                       tid;         
  } dcache_rtrn_t;
  
  
  typedef enum logic [4:0] {
    L15_LOAD_RQ     = 5'b00000, 
    L15_IMISS_RQ    = 5'b10000, 
    L15_STORE_RQ    = 5'b00001, 
    L15_ATOMIC_RQ   = 5'b00110, 
    
    
    
    L15_STRLOAD_RQ  = 5'b00100, 
    L15_STRST_RQ    = 5'b00101, 
    L15_STQ_RQ      = 5'b00111, 
    L15_INT_RQ      = 5'b01001, 
    L15_FWD_RQ      = 5'b01101, 
    L15_FWD_RPY     = 5'b01110, 
    L15_RSVD_RQ     = 5'b11111  
  } l15_reqtypes_t;
  
  typedef enum logic [3:0] {
    L15_LOAD_RET               = 4'b0000, 
    
    L15_ST_ACK                 = 4'b0100, 
    
    L15_INT_RET                = 4'b0111, 
    L15_TEST_RET               = 4'b0101, 
    L15_FP_RET                 = 4'b1000, 
    L15_IFILL_RET              = 4'b0001, 
    L15_EVICT_REQ              = 4'b0011, 
    L15_ERR_RET                = 4'b1100, 
    L15_STRLOAD_RET            = 4'b0010, 
    L15_STRST_ACK              = 4'b0110, 
    L15_FWD_RQ_RET             = 4'b1010, 
    L15_FWD_RPY_RET            = 4'b1011, 
    L15_RSVD_RET               = 4'b1111, 
    L15_CPX_RESTYPE_ATOMIC_RES = 4'b1110  
  } l15_rtrntypes_t;
  typedef struct packed {
    logic                              l15_val;                   
    logic                              l15_req_ack;               
    l15_reqtypes_t                     l15_rqtype;                
    logic                              l15_nc;                    
    logic [2:0]                        l15_size;                  
    logic [L15_TID_WIDTH-1:0]          l15_threadid;              
    logic                              l15_prefetch;              
    logic                              l15_invalidate_cacheline;  
    logic                              l15_blockstore;            
    logic                              l15_blockinitstore;        
    logic [L15_WAY_WIDTH-1:0]          l15_l1rplway;              
    logic [39:0]                       l15_address;               
    logic [63:0]                       l15_data;                  
    logic [63:0]                       l15_data_next_entry;       
    logic [L15_TLB_CSM_WIDTH-1:0]      l15_csm_data;              
    logic [3:0]                        l15_amo_op;                
  } l15_req_t;
  typedef struct packed {
    logic                              l15_ack;                   
    logic                              l15_header_ack;            
    logic                              l15_val;                   
    l15_rtrntypes_t                    l15_returntype;            
    logic                              l15_l2miss;                
    logic [1:0]                        l15_error;                 
    logic                              l15_noncacheable;          
    logic                              l15_atomic;                
    logic [L15_TID_WIDTH-1:0]          l15_threadid;              
    logic                              l15_prefetch;              
    logic                              l15_f4b;                   
    logic [63:0]                       l15_data_0;                
    logic [63:0]                       l15_data_1;                
    logic [63:0]                       l15_data_2;                
    logic [63:0]                       l15_data_3;                
    logic                              l15_inval_icache_all_way;  
    logic                              l15_inval_dcache_all_way;  
    logic [15:4]                       l15_inval_address_15_4;    
    logic                              l15_cross_invalidate;      
    logic [L15_WAY_WIDTH-1:0]          l15_cross_invalidate_way;  
    logic                              l15_inval_dcache_inval;    
    logic                              l15_inval_icache_inval;    
    logic [L15_WAY_WIDTH-1:0]          l15_inval_way;             
    logic                              l15_blockinitstore;        
  } l15_rtrn_t;
  
  function automatic logic[63:0] swendian64(input logic[63:0] in);
    automatic logic[63:0] out;
    for(int k=0; k<64;k+=8)begin
        out[k +: 8] = in[63-k -: 8];
    end
    return out;
  endfunction
  function automatic logic [ariane_pkg::ICACHE_SET_ASSOC-1:0] icache_way_bin2oh (
    input logic [L1I_WAY_WIDTH-1:0] in
  );
    logic [ariane_pkg::ICACHE_SET_ASSOC-1:0] out;
    out     = '0;
    out[in] = 1'b1;
    return out;
  endfunction
  function automatic logic [ariane_pkg::DCACHE_SET_ASSOC-1:0] dcache_way_bin2oh (
    input logic [L1D_WAY_WIDTH-1:0] in
  );
    logic [ariane_pkg::DCACHE_SET_ASSOC-1:0] out;
    out     = '0;
    out[in] = 1'b1;
    return out;
  endfunction
  function automatic logic [DCACHE_NUM_BANKS-1:0] dcache_cl_bin2oh (
    input logic [DCACHE_NUM_BANKS_WIDTH-1:0] in
  );
    logic [DCACHE_NUM_BANKS-1:0] out;
    out     = '0;
    out[in] = 1'b1;
    return out;
  endfunction
  function automatic logic [5:0] popcnt64 (
    input logic [63:0] in
  );
    logic [5:0] cnt= 0;
    foreach (in[k]) begin
      cnt += 6'(in[k]);
    end
    return cnt;
  endfunction : popcnt64
  function automatic logic [7:0] toByteEnable8(
    input logic [2:0] offset,
    input logic [1:0] size
  );
    logic [7:0] be;
    be = '0;
    unique case(size)
      2'b00:   be[offset]       = '1; 
      2'b01:   be[offset +:2 ]  = '1; 
      2'b10:   be[offset +:4 ]  = '1; 
      default: be               = '1; 
    endcase 
    return be;
  endfunction : toByteEnable8
  
  function automatic logic [63:0] repData64(
    input logic [63:0] data,
    input logic [2:0]  offset,
    input logic [1:0]  size
  );
    logic [63:0] out;
    unique case(size)
      2'b00:   for(int k=0; k<8; k++) out[k*8  +: 8]    = data[offset*8 +: 8];  
      2'b01:   for(int k=0; k<4; k++) out[k*16 +: 16]   = data[offset*8 +: 16]; 
      2'b10:   for(int k=0; k<2; k++) out[k*32 +: 32]   = data[offset*8 +: 32]; 
      default: out   = data; 
    endcase 
    return out;
  endfunction : repData64
  
  
  
  function automatic logic [1:0] toSize64(
    input logic  [7:0] be
  );
    logic [1:0] size;
    unique case(be)
      8'b1111_1111:                                           size = 2'b11;  
      8'b0000_1111, 8'b1111_0000:                             size = 2'b10; 
      8'b1100_0000, 8'b0011_0000, 8'b0000_1100, 8'b0000_0011: size = 2'b01; 
      default:                                                size = 2'b00; 
    endcase 
    return size;
  endfunction : toSize64
  
  
  
  
  
  
  function automatic logic [riscv::PLEN-1:0] paddrSizeAlign(
    input logic [riscv::PLEN-1:0] paddr,
    input logic [2:0]  size
  );
    logic [riscv::PLEN-1:0] out;
    out = paddr;
    unique case (size)
      3'b001: out[0:0]                     = '0;
      3'b010: out[1:0]                     = '0;
      3'b011: out[2:0]                     = '0;
      3'b111: out[DCACHE_OFFSET_WIDTH-1:0] = '0;
      default: ;
    endcase
    return out;
  endfunction : paddrSizeAlign
endpackage
package std_cache_pkg;
    
    localparam DCACHE_BYTE_OFFSET = $clog2(ariane_pkg::DCACHE_LINE_WIDTH/8);
    localparam DCACHE_NUM_WORDS   = 2**(ariane_pkg::DCACHE_INDEX_WIDTH-DCACHE_BYTE_OFFSET);
    localparam DCACHE_DIRTY_WIDTH = ariane_pkg::DCACHE_SET_ASSOC*2;
    
    typedef struct packed {
        logic [1:0]      id;     
        logic            valid;
        logic            we;
        logic [55:0]     addr;
        logic [7:0][7:0] wdata;
        logic [7:0]      be;
    } mshr_t;
    typedef struct packed {
        logic         valid;
        logic [63:0]  addr;
        logic [7:0]   be;
        logic [1:0]   size;
        logic         we;
        logic [63:0]  wdata;
        logic         bypass;
    } miss_req_t;
    typedef struct packed {
        logic [ariane_pkg::DCACHE_TAG_WIDTH-1:0]  tag;    
        logic [ariane_pkg::DCACHE_LINE_WIDTH-1:0] data;   
        logic                                     valid;  
        logic                                     dirty;  
    } cache_line_t;
    
    typedef struct packed {
        logic [(ariane_pkg::DCACHE_TAG_WIDTH+7)/8-1:0]  tag;    
        logic [(ariane_pkg::DCACHE_LINE_WIDTH+7)/8-1:0] data;   
        logic [ariane_pkg::DCACHE_SET_ASSOC-1:0]        vldrty; 
    } cl_be_t;
    
    function automatic logic [$clog2(ariane_pkg::DCACHE_SET_ASSOC)-1:0] one_hot_to_bin (
        input logic [ariane_pkg::DCACHE_SET_ASSOC-1:0] in
    );
        for (int unsigned i = 0; i < ariane_pkg::DCACHE_SET_ASSOC; i++) begin
            if (in[i])
                return i;
        end
    endfunction
    
    function automatic logic [ariane_pkg::DCACHE_SET_ASSOC-1:0] get_victim_cl (
        input logic [ariane_pkg::DCACHE_SET_ASSOC-1:0] valid_dirty
    );
        
        logic [ariane_pkg::DCACHE_SET_ASSOC-1:0] oh = '0;
        for (int unsigned i = 0; i < ariane_pkg::DCACHE_SET_ASSOC; i++) begin
            if (valid_dirty[i]) begin
                oh[i] = 1'b1;
                return oh;
            end
        end
    endfunction
endpackage : std_cache_pkg
interface AXI_BUS #(
  parameter AXI_ADDR_WIDTH = -1,
  parameter AXI_DATA_WIDTH = -1,
  parameter AXI_ID_WIDTH   = -1,
  parameter AXI_USER_WIDTH = -1
);
  import axi_pkg::*;
  localparam AXI_STRB_WIDTH = AXI_DATA_WIDTH / 8;
  typedef logic [AXI_ID_WIDTH-1:0]   id_t;
  typedef logic [AXI_ADDR_WIDTH-1:0] addr_t;
  typedef logic [AXI_DATA_WIDTH-1:0] data_t;
  typedef logic [AXI_STRB_WIDTH-1:0] strb_t;
  typedef logic [AXI_USER_WIDTH-1:0] user_t;
  typedef logic [5:0] atop_t;
  id_t        aw_id;
  addr_t      aw_addr;
  logic [7:0] aw_len;
  logic [2:0] aw_size;
  burst_t     aw_burst;
  logic       aw_lock;
  cache_t     aw_cache;
  prot_t      aw_prot;
  qos_t       aw_qos;
  atop_t      aw_atop;
  region_t    aw_region;
  user_t      aw_user;
  logic       aw_valid;
  logic       aw_ready;
  data_t      w_data;
  strb_t      w_strb;
  logic       w_last;
  user_t      w_user;
  logic       w_valid;
  logic       w_ready;
  id_t        b_id;
  resp_t      b_resp;
  user_t      b_user;
  logic       b_valid;
  logic       b_ready;
  id_t        ar_id;
  addr_t      ar_addr;
  logic [7:0] ar_len;
  logic [2:0] ar_size;
  burst_t     ar_burst;
  logic       ar_lock;
  cache_t     ar_cache;
  prot_t      ar_prot;
  qos_t       ar_qos;
  region_t    ar_region;
  user_t      ar_user;
  logic       ar_valid;
  logic       ar_ready;
  id_t        r_id;
  data_t      r_data;
  resp_t      r_resp;
  logic       r_last;
  user_t      r_user;
  logic       r_valid;
  logic       r_ready;
  modport Master (
    output aw_id, aw_addr, aw_len, aw_size, aw_burst, aw_lock, aw_cache, aw_prot, aw_qos, aw_atop, aw_region, aw_user, aw_valid, input aw_ready,
    output w_data, w_strb, w_last, w_user, w_valid, input w_ready,
    input b_id, b_resp, b_user, b_valid, output b_ready,
    output ar_id, ar_addr, ar_len, ar_size, ar_burst, ar_lock, ar_cache, ar_prot, ar_qos, ar_region, ar_user, ar_valid, input ar_ready,
    input r_id, r_data, r_resp, r_last, r_user, r_valid, output r_ready
  );
  modport Slave (
    input aw_id, aw_addr, aw_len, aw_size, aw_burst, aw_lock, aw_cache, aw_prot, aw_qos, aw_atop, aw_region, aw_user, aw_valid, output aw_ready,
    input w_data, w_strb, w_last, w_user, w_valid, output w_ready,
    output b_id, b_resp, b_user, b_valid, input b_ready,
    input ar_id, ar_addr, ar_len, ar_size, ar_burst, ar_lock, ar_cache, ar_prot, ar_qos, ar_region, ar_user, ar_valid, output ar_ready,
    output r_id, r_data, r_resp, r_last, r_user, r_valid, input r_ready
  );
endinterface
interface AXI_BUS_ASYNC
#(
  parameter AXI_ADDR_WIDTH = -1,
  parameter AXI_DATA_WIDTH = -1,
  parameter AXI_ID_WIDTH   = -1,
  parameter AXI_USER_WIDTH = -1,
  parameter BUFFER_WIDTH   = -1
);
  localparam AXI_STRB_WIDTH = AXI_DATA_WIDTH / 8;
  logic [AXI_ID_WIDTH-1:0]    aw_id;
  logic [AXI_ADDR_WIDTH-1:0]  aw_addr;
  logic [7:0]                 aw_len;
  logic [2:0]                 aw_size;
  logic [1:0]                 aw_burst;
  logic                       aw_lock;
  logic [3:0]                 aw_cache;
  logic [2:0]                 aw_prot;
  logic [3:0]                 aw_qos;
  logic [5:0]                 aw_atop;
  logic [3:0]                 aw_region;
  logic [AXI_USER_WIDTH-1:0]  aw_user;
  logic [BUFFER_WIDTH-1:0]    aw_writetoken;
  logic [BUFFER_WIDTH-1:0]    aw_readpointer;
  logic [AXI_DATA_WIDTH-1:0]  w_data;
  logic [AXI_STRB_WIDTH-1:0]  w_strb;
  logic                       w_last;
  logic [AXI_USER_WIDTH-1:0]  w_user;
  logic [BUFFER_WIDTH-1:0]    w_writetoken;
  logic [BUFFER_WIDTH-1:0]    w_readpointer;
  logic [AXI_ID_WIDTH-1:0]    b_id;
  logic [1:0]                 b_resp;
  logic [AXI_USER_WIDTH-1:0]  b_user;
  logic [BUFFER_WIDTH-1:0]    b_writetoken;
  logic [BUFFER_WIDTH-1:0]    b_readpointer;
  logic [AXI_ID_WIDTH-1:0]    ar_id;
  logic [AXI_ADDR_WIDTH-1:0]  ar_addr;
  logic [7:0]                 ar_len;
  logic [2:0]                 ar_size;
  logic [1:0]                 ar_burst;
  logic                       ar_lock;
  logic [3:0]                 ar_cache;
  logic [2:0]                 ar_prot;
  logic [3:0]                 ar_qos;
  logic [3:0]                 ar_region;
  logic [AXI_USER_WIDTH-1:0]  ar_user;
  logic [BUFFER_WIDTH-1:0]    ar_writetoken;
  logic [BUFFER_WIDTH-1:0]    ar_readpointer;
  logic [AXI_ID_WIDTH-1:0]    r_id;
  logic [AXI_DATA_WIDTH-1:0]  r_data;
  logic [1:0]                 r_resp;
  logic                       r_last;
  logic [AXI_USER_WIDTH-1:0]  r_user;
  logic [BUFFER_WIDTH-1:0]    r_writetoken;
  logic [BUFFER_WIDTH-1:0]    r_readpointer;
  modport Master (
    output aw_id, aw_addr, aw_len, aw_size, aw_burst, aw_lock, aw_cache, aw_prot, aw_qos, aw_atop, aw_region, aw_user, aw_writetoken, input aw_readpointer,
    output w_data, w_strb, w_last, w_user, w_writetoken, input w_readpointer,
    input b_id, b_resp, b_user, b_writetoken, output b_readpointer,
    output ar_id, ar_addr, ar_len, ar_size, ar_burst, ar_lock, ar_cache, ar_prot, ar_qos, ar_region, ar_user, ar_writetoken, input ar_readpointer,
    input r_id, r_data, r_resp, r_last, r_user, r_writetoken, output r_readpointer
  );
  modport Slave (
    input aw_id, aw_addr, aw_len, aw_size, aw_burst, aw_lock, aw_cache, aw_prot, aw_qos, aw_atop, aw_region, aw_user, aw_writetoken, output aw_readpointer,
    input w_data, w_strb, w_last, w_user, w_writetoken, output w_readpointer,
    output b_id, b_resp, b_user, b_writetoken, input b_readpointer,
    input ar_id, ar_addr, ar_len, ar_size, ar_burst, ar_lock, ar_cache, ar_prot, ar_qos, ar_region, ar_user, ar_writetoken, output ar_readpointer,
    output r_id, r_data, r_resp, r_last, r_user, r_writetoken, input r_readpointer
  );
endinterface
interface AXI_LITE #(
  parameter AXI_ADDR_WIDTH = -1,
  parameter AXI_DATA_WIDTH = -1
);
  import axi_pkg::*;
  localparam AXI_STRB_WIDTH = AXI_DATA_WIDTH / 8;
  typedef logic [AXI_ADDR_WIDTH-1:0] addr_t;
  typedef logic [AXI_DATA_WIDTH-1:0] data_t;
  typedef logic [AXI_STRB_WIDTH-1:0] strb_t;
  
  addr_t aw_addr;
  logic  aw_valid;
  logic  aw_ready;
  data_t w_data;
  strb_t w_strb;
  logic  w_valid;
  logic  w_ready;
  resp_t b_resp;
  logic  b_valid;
  logic  b_ready;
  addr_t ar_addr;
  logic  ar_valid;
  logic  ar_ready;
  data_t r_data;
  resp_t r_resp;
  logic  r_valid;
  logic  r_ready;
  modport Master (
    output aw_addr, aw_valid, input aw_ready,
    output w_data, w_strb, w_valid, input w_ready,
    input b_resp, b_valid, output b_ready,
    output ar_addr, ar_valid, input ar_ready,
    input r_data, r_resp, r_valid, output r_ready
  );
  modport Slave (
    input aw_addr, aw_valid, output aw_ready,
    input w_data, w_strb, w_valid, output w_ready,
    output b_resp, b_valid, input b_ready,
    input ar_addr, ar_valid, output ar_ready,
    output r_data, r_resp, r_valid, input r_ready
  );
  
  modport out (
    output aw_addr, aw_valid, input aw_ready,
    output w_data, w_strb, w_valid, input w_ready,
    input b_resp, b_valid, output b_ready,
    output ar_addr, ar_valid, input ar_ready,
    input r_data, r_resp, r_valid, output r_ready
  );
  
  modport in (
    input aw_addr, aw_valid, output aw_ready,
    input w_data, w_strb, w_valid, output w_ready,
    output b_resp, b_valid, input b_ready,
    input ar_addr, ar_valid, output ar_ready,
    output r_data, r_resp, r_valid, input r_ready
  );
endinterface
interface AXI_ROUTING_RULES #(
  
  parameter int AXI_ADDR_WIDTH = -1,
  
  parameter int NUM_SLAVE  = -1,
  
  parameter int NUM_RULES  = -1
);
  struct packed {
    logic enabled;
    logic [AXI_ADDR_WIDTH-1:0] mask;
    logic [AXI_ADDR_WIDTH-1:0] base;
  } [NUM_RULES-1:0] rules [NUM_SLAVE];
  modport xbar(input rules);
  modport cfg(output rules);
endinterface
interface AXI_ARBITRATION #(
  
  parameter int NUM_REQ = -1
);
  
  logic [NUM_REQ-1:0] in_req;
  logic [NUM_REQ-1:0] in_ack;
  
  logic out_req;
  logic out_ack;
  logic [$clog2(NUM_REQ)-1:0] out_sel;
  
  modport arb(input  in_req, out_ack, output out_req, out_sel, in_ack);
  
  modport req(output in_req, out_ack, input  out_req, out_sel, in_ack);
endinterface
module sram #(
    parameter DATA_WIDTH = 64,
    parameter NUM_WORDS  = 1024,
    parameter OUT_REGS   = 0,    
    parameter DROMAJO_RAM  = 0
)(
   input  logic                          clk_i,
   input  logic                          rst_ni,
   input  logic                          req_i,
   input  logic                          we_i,
   input  logic [$clog2(NUM_WORDS)-1:0]  addr_i,
   input  logic [DATA_WIDTH-1:0]         wdata_i,
   input  logic [(DATA_WIDTH+7)/8-1:0]   be_i,
   output logic [DATA_WIDTH-1:0]         rdata_o
);
localparam DATA_WIDTH_ALIGNED = ((DATA_WIDTH+63)/64)*64;
localparam BE_WIDTH_ALIGNED   = (((DATA_WIDTH+7)/8+7)/8)*8;
logic [DATA_WIDTH_ALIGNED-1:0]  wdata_aligned;
logic [BE_WIDTH_ALIGNED-1:0]    be_aligned;
logic [DATA_WIDTH_ALIGNED-1:0]  rdata_aligned;
always_comb begin : p_align
    wdata_aligned                    ='0;
    be_aligned                       ='0;
    wdata_aligned[DATA_WIDTH-1:0]    = wdata_i;
    be_aligned[BE_WIDTH_ALIGNED-1:0] = be_i;
    rdata_o = rdata_aligned[DATA_WIDTH-1:0];
end
  for (genvar k = 0; k<(DATA_WIDTH+63)/64; k++) begin : gen_cut
    if (DROMAJO_RAM) begin : gen_dromajo
      dromajo_ram #(
        .ADDR_WIDTH($clog2(NUM_WORDS)),
        .DATA_DEPTH(NUM_WORDS),
        .OUT_REGS (0)
      ) i_ram (
          .Clk_CI    ( clk_i                     ),
          .Rst_RBI   ( rst_ni                    ),
          .CSel_SI   ( req_i                     ),
          .WrEn_SI   ( we_i                      ),
          .BEn_SI    ( be_aligned[k*8 +: 8]      ),
          .WrData_DI ( wdata_aligned[k*64 +: 64] ),
          .Addr_DI   ( addr_i                    ),
          .RdData_DO ( rdata_aligned[k*64 +: 64] )
      );
    end else begin : gen_mem
      
      SyncSpRamBeNx64 #(
        .ADDR_WIDTH($clog2(NUM_WORDS)),
        .DATA_DEPTH(NUM_WORDS),
        .OUT_REGS (0),
        
        
        .SIM_INIT (1)
      ) i_ram (
          .Clk_CI    ( clk_i                     ),
          .Rst_RBI   ( rst_ni                    ),
          .CSel_SI   ( req_i                     ),
          .WrEn_SI   ( we_i                      ),
          .BEn_SI    ( be_aligned[k*8 +: 8]      ),
          .WrData_DI ( wdata_aligned[k*64 +: 64] ),
          .Addr_DI   ( addr_i                    ),
          .RdData_DO ( rdata_aligned[k*64 +: 64] )
      );
    end
  end
endmodule : sram
module axi_master_connect (
    input  ariane_axi::req_t    axi_req_i,
    output ariane_axi::resp_t   axi_resp_o,
    AXI_BUS.Master master
);
    assign master.aw_id         = axi_req_i.aw.id;
    assign master.aw_addr       = axi_req_i.aw.addr;
    assign master.aw_len        = axi_req_i.aw.len;
    assign master.aw_size       = axi_req_i.aw.size;
    assign master.aw_burst      = axi_req_i.aw.burst;
    assign master.aw_lock       = axi_req_i.aw.lock;
    assign master.aw_cache      = axi_req_i.aw.cache;
    assign master.aw_prot       = axi_req_i.aw.prot;
    assign master.aw_qos        = axi_req_i.aw.qos;
    assign master.aw_atop       = axi_req_i.aw.atop;
    assign master.aw_region     = axi_req_i.aw.region;
    assign master.aw_user       = '0;
    assign master.aw_valid      = axi_req_i.aw_valid;
    assign axi_resp_o.aw_ready  = master.aw_ready;
    assign master.w_data        = axi_req_i.w.data;
    assign master.w_strb        = axi_req_i.w.strb;
    assign master.w_last        = axi_req_i.w.last;
    assign master.w_user        = '0;
    assign master.w_valid       = axi_req_i.w_valid;
    assign axi_resp_o.w_ready   = master.w_ready;
    assign axi_resp_o.b.id      = master.b_id;
    assign axi_resp_o.b.resp    = master.b_resp;
    assign axi_resp_o.b_valid   = master.b_valid;
    assign master.b_ready       = axi_req_i.b_ready;
    assign master.ar_id         = axi_req_i.ar.id;
    assign master.ar_addr       = axi_req_i.ar.addr;
    assign master.ar_len        = axi_req_i.ar.len;
    assign master.ar_size       = axi_req_i.ar.size;
    assign master.ar_burst      = axi_req_i.ar.burst;
    assign master.ar_lock       = axi_req_i.ar.lock;
    assign master.ar_cache      = axi_req_i.ar.cache;
    assign master.ar_prot       = axi_req_i.ar.prot;
    assign master.ar_qos        = axi_req_i.ar.qos;
    assign master.ar_region     = axi_req_i.ar.region;
    assign master.ar_user       = '0;
    assign master.ar_valid      = axi_req_i.ar_valid;
    assign axi_resp_o.ar_ready  = master.ar_ready;
    assign axi_resp_o.r.id      = master.r_id;
    assign axi_resp_o.r.data    = master.r_data;
    assign axi_resp_o.r.resp    = master.r_resp;
    assign axi_resp_o.r.last    = master.r_last;
    assign axi_resp_o.r_valid   = master.r_valid;
    assign master.r_ready       = axi_req_i.r_ready;
endmodule
module axi_master_connect_rev (
    output ariane_axi::req_t    axi_req_o,
    input  ariane_axi::resp_t   axi_resp_i,
    AXI_BUS.Slave master
);
    assign  axi_req_o.aw.atop    = '0; 
    assign  axi_req_o.aw.id      = master.aw_id;
    assign  axi_req_o.aw.addr    = master.aw_addr;
    assign  axi_req_o.aw.len     = master.aw_len;
    assign  axi_req_o.aw.size    = master.aw_size;
    assign  axi_req_o.aw.burst   = master.aw_burst;
    assign  axi_req_o.aw.lock    = master.aw_lock;
    assign  axi_req_o.aw.cache   = master.aw_cache;
    assign  axi_req_o.aw.prot    = master.aw_prot;
    assign  axi_req_o.aw.qos     = master.aw_qos;
    assign  axi_req_o.aw.region  = master.aw_region;
    
    assign  axi_req_o.aw_valid   = master.aw_valid;
    assign  master.aw_ready       = axi_resp_i.aw_ready;
    assign  axi_req_o.w.data     = master.w_data;
    assign  axi_req_o.w.strb     = master.w_strb;
    assign  axi_req_o.w.last     = master.w_last;
    
    assign  axi_req_o.w_valid    = master.w_valid;
    assign  master.w_ready        = axi_resp_i.w_ready;
    assign  master.b_id           = axi_resp_i.b.id;
    assign  master.b_resp         = axi_resp_i.b.resp;
    assign  master.b_valid        = axi_resp_i.b_valid;
    assign  axi_req_o.b_ready    = master.b_ready;
    assign  axi_req_o.ar.id      = master.ar_id;
    assign  axi_req_o.ar.addr    = master.ar_addr;
    assign  axi_req_o.ar.len     = master.ar_len;
    assign  axi_req_o.ar.size    = master.ar_size;
    assign  axi_req_o.ar.burst   = master.ar_burst;
    assign  axi_req_o.ar.lock    = master.ar_lock;
    assign  axi_req_o.ar.cache   = master.ar_cache;
    assign  axi_req_o.ar.prot    = master.ar_prot;
    assign  axi_req_o.ar.qos     = master.ar_qos;
    assign  axi_req_o.ar.region  = master.ar_region;
    
    assign  axi_req_o.ar_valid   = master.ar_valid;
    assign  master.ar_ready       = axi_resp_i.ar_ready;
    assign  master.r_id           = axi_resp_i.r.id;
    assign  master.r_data         = axi_resp_i.r.data;
    assign  master.r_resp         = axi_resp_i.r.resp;
    assign  master.r_last         = axi_resp_i.r.last;
    assign  master.r_valid        = axi_resp_i.r_valid;
    assign  axi_req_o.r_ready    = master.r_ready;
endmodule
module axi_slave_connect (
    output ariane_axi::req_t    axi_req_o,
    input  ariane_axi::resp_t   axi_resp_i,
    AXI_BUS.Slave slave
);
    assign  axi_req_o.aw.id      = slave.aw_id;
    assign  axi_req_o.aw.addr    = slave.aw_addr;
    assign  axi_req_o.aw.len     = slave.aw_len;
    assign  axi_req_o.aw.size    = slave.aw_size;
    assign  axi_req_o.aw.burst   = slave.aw_burst;
    assign  axi_req_o.aw.lock    = slave.aw_lock;
    assign  axi_req_o.aw.cache   = slave.aw_cache;
    assign  axi_req_o.aw.prot    = slave.aw_prot;
    assign  axi_req_o.aw.qos     = slave.aw_qos;
    assign  axi_req_o.aw.atop    = slave.aw_atop;
    assign  axi_req_o.aw.region  = slave.aw_region;
    
    assign  axi_req_o.aw_valid   = slave.aw_valid;
    assign  slave.aw_ready       = axi_resp_i.aw_ready;
    assign  axi_req_o.w.data     = slave.w_data;
    assign  axi_req_o.w.strb     = slave.w_strb;
    assign  axi_req_o.w.last     = slave.w_last;
    
    assign  axi_req_o.w_valid    = slave.w_valid;
    assign  slave.w_ready        = axi_resp_i.w_ready;
    assign  slave.b_id           = axi_resp_i.b.id;
    assign  slave.b_resp         = axi_resp_i.b.resp;
    assign  slave.b_valid        = axi_resp_i.b_valid;
    assign  slave.b_user         = 1'b0;
    assign  axi_req_o.b_ready    = slave.b_ready;
    assign  axi_req_o.ar.id      = slave.ar_id;
    assign  axi_req_o.ar.addr    = slave.ar_addr;
    assign  axi_req_o.ar.len     = slave.ar_len;
    assign  axi_req_o.ar.size    = slave.ar_size;
    assign  axi_req_o.ar.burst   = slave.ar_burst;
    assign  axi_req_o.ar.lock    = slave.ar_lock;
    assign  axi_req_o.ar.cache   = slave.ar_cache;
    assign  axi_req_o.ar.prot    = slave.ar_prot;
    assign  axi_req_o.ar.qos     = slave.ar_qos;
    assign  axi_req_o.ar.region  = slave.ar_region;
    
    assign  axi_req_o.ar_valid   = slave.ar_valid;
    assign  slave.ar_ready       = axi_resp_i.ar_ready;
    assign  slave.r_id           = axi_resp_i.r.id;
    assign  slave.r_data         = axi_resp_i.r.data;
    assign  slave.r_resp         = axi_resp_i.r.resp;
    assign  slave.r_last         = axi_resp_i.r.last;
    assign  slave.r_valid        = axi_resp_i.r_valid;
    assign  slave.r_user         = 1'b0;
    assign  axi_req_o.r_ready    = slave.r_ready;
endmodule
module axi_slave_connect_rev (
    input  ariane_axi::req_t    axi_req_i,
    output ariane_axi::resp_t   axi_resp_o,
    AXI_BUS.Master slave
);
    assign slave.aw_id         = axi_req_i.aw.id;
    assign slave.aw_addr       = axi_req_i.aw.addr;
    assign slave.aw_len        = axi_req_i.aw.len;
    assign slave.aw_size       = axi_req_i.aw.size;
    assign slave.aw_burst      = axi_req_i.aw.burst;
    assign slave.aw_lock       = axi_req_i.aw.lock;
    assign slave.aw_cache      = axi_req_i.aw.cache;
    assign slave.aw_prot       = axi_req_i.aw.prot;
    assign slave.aw_qos        = axi_req_i.aw.qos;
    assign slave.aw_region     = axi_req_i.aw.region;
    assign slave.aw_user       = '0;
    assign slave.aw_valid      = axi_req_i.aw_valid;
    assign axi_resp_o.aw_ready = slave.aw_ready;
    assign slave.w_data        = axi_req_i.w.data;
    assign slave.w_strb        = axi_req_i.w.strb;
    assign slave.w_last        = axi_req_i.w.last;
    assign slave.w_user        = '0;
    assign slave.w_valid       = axi_req_i.w_valid;
    assign axi_resp_o.w_ready  = slave.w_ready;
    assign axi_resp_o.b.id     = slave.b_id;
    assign axi_resp_o.b.resp   = slave.b_resp;
    assign axi_resp_o.b_valid  = slave.b_valid;
    assign slave.b_ready       = axi_req_i.b_ready;
    assign slave.ar_id         = axi_req_i.ar.id;
    assign slave.ar_addr       = axi_req_i.ar.addr;
    assign slave.ar_len        = axi_req_i.ar.len;
    assign slave.ar_size       = axi_req_i.ar.size;
    assign slave.ar_burst      = axi_req_i.ar.burst;
    assign slave.ar_lock       = axi_req_i.ar.lock;
    assign slave.ar_cache      = axi_req_i.ar.cache;
    assign slave.ar_prot       = axi_req_i.ar.prot;
    assign slave.ar_qos        = axi_req_i.ar.qos;
    assign slave.ar_region     = axi_req_i.ar.region;
    assign slave.ar_user       = '0;
    assign slave.ar_valid      = axi_req_i.ar_valid;
    assign axi_resp_o.ar_ready = slave.ar_ready;
    assign axi_resp_o.r.id     = slave.r_id;
    assign axi_resp_o.r.data   = slave.r_data;
    assign axi_resp_o.r.resp   = slave.r_resp;
    assign axi_resp_o.r.last   = slave.r_last;
    assign axi_resp_o.r_valid  = slave.r_valid;
    assign slave.r_ready       = axi_req_i.r_ready;
endmodule
  
module SyncSpRamBeNx64
#(
  parameter ADDR_WIDTH = 10,
  parameter DATA_DEPTH = 1024, 
  parameter OUT_REGS   = 0,    
  parameter SIM_INIT   = 0     
                               
                               
)(
  input  logic                  Clk_CI,
  input  logic                  Rst_RBI,
  input  logic                  CSel_SI,
  input  logic                  WrEn_SI,
  input  logic [7:0]            BEn_SI,
  input  logic [63:0]           WrData_DI,
  input  logic [ADDR_WIDTH-1:0] Addr_DI,
  output logic [63:0]           RdData_DO
);
  
  
  
  
  localparam DATA_BYTES = 8;
  logic [DATA_BYTES*8-1:0] RdData_DN;
  logic [DATA_BYTES*8-1:0] RdData_DP;
  
  
  
  
    logic [DATA_BYTES*8-1:0] Mem_DP[DATA_DEPTH-1:0];
    always_ff @(posedge Clk_CI) begin
      
      automatic logic [63:0] val;
      if(Rst_RBI == 1'b0 && SIM_INIT>0) begin
        for(int k=0; k<DATA_DEPTH;k++) begin
          if(SIM_INIT==1) val = '0;
      
      
          else val = 64'hdeadbeefdeadbeef;
          Mem_DP[k] = val;
        end
      end else
      
      if(CSel_SI) begin
        if(WrEn_SI) begin
          if(BEn_SI[0]) Mem_DP[Addr_DI][7:0]   <= WrData_DI[7:0];
          if(BEn_SI[1]) Mem_DP[Addr_DI][15:8]  <= WrData_DI[15:8];
          if(BEn_SI[2]) Mem_DP[Addr_DI][23:16] <= WrData_DI[23:16];
          if(BEn_SI[3]) Mem_DP[Addr_DI][31:24] <= WrData_DI[31:24];
          if(BEn_SI[4]) Mem_DP[Addr_DI][39:32] <= WrData_DI[39:32];
          if(BEn_SI[5]) Mem_DP[Addr_DI][47:40] <= WrData_DI[47:40];
          if(BEn_SI[6]) Mem_DP[Addr_DI][55:48] <= WrData_DI[55:48];
          if(BEn_SI[7]) Mem_DP[Addr_DI][63:56] <= WrData_DI[63:56];
        end
        RdData_DN <= Mem_DP[Addr_DI];
      end
    end
  
  
  
  
  
      
      
  
  
  
  
  
  generate
    if (OUT_REGS>0) begin : g_outreg
      always_ff @(posedge Clk_CI or negedge Rst_RBI) begin
        if(Rst_RBI == 1'b0)
        begin
          RdData_DP  <= 0;
        end
        else
        begin
          RdData_DP  <= RdData_DN;
        end
      end
    end
  endgenerate 
  
  generate
    if (OUT_REGS==0) begin : g_oureg_byp
      assign RdData_DP  = RdData_DN;
    end
  endgenerate
  assign RdData_DO = RdData_DP;
  
  
  
  
  assert property
    (@(posedge Clk_CI) (longint'(2)**longint'(ADDR_WIDTH) >= longint'(DATA_DEPTH)))
    else $error("depth out of bounds");
  
  
    
    
  
endmodule 
module dromajo_ram
#(
  parameter ADDR_WIDTH = 10,
  parameter DATA_DEPTH = 1024, 
  parameter OUT_REGS   = 0     
)(
  input  logic                  Clk_CI,
  input  logic                  Rst_RBI,
  input  logic                  CSel_SI,
  input  logic                  WrEn_SI,
  input  logic [7:0]            BEn_SI,
  input  logic [63:0]           WrData_DI,
  input  logic [ADDR_WIDTH-1:0] Addr_DI,
  output logic [63:0]           RdData_DO
);
  
  
  
  
  localparam DATA_BYTES = 8;
  logic [DATA_BYTES*8-1:0] RdData_DN;
  logic [DATA_BYTES*8-1:0] RdData_DP;
  logic [DATA_BYTES*8-1:0] Mem_DP[DATA_DEPTH-1:0];
  
  
  
  
  initial begin
    integer hex_file, num_bytes;
    longint address, value;
    string f_name;
    
    for (int k=0; k<DATA_DEPTH; k++) begin
      Mem_DP[k] = 0;
    end
    
    if ($value$plusargs("checkpoint=%s", f_name)) begin
      hex_file = $fopen({f_name,".mainram.hex"}, "r");
      while (!$feof(hex_file)) begin
        num_bytes = $fscanf(hex_file, "%d %h\n", address, value);
        
        Mem_DP[address] = value;
      end
      $display("Done syncing RAM with dromajo...\n");
    end else begin
      $display("Failed syncing RAM: provide path to a checkpoint.\n");
    end
  end
  always @(posedge Clk_CI) begin
    if(CSel_SI) begin
      if(WrEn_SI) begin
        if(BEn_SI[0]) Mem_DP[Addr_DI][7:0]   <= WrData_DI[7:0];
        if(BEn_SI[1]) Mem_DP[Addr_DI][15:8]  <= WrData_DI[15:8];
        if(BEn_SI[2]) Mem_DP[Addr_DI][23:16] <= WrData_DI[23:16];
        if(BEn_SI[3]) Mem_DP[Addr_DI][31:24] <= WrData_DI[31:24];
        if(BEn_SI[4]) Mem_DP[Addr_DI][39:32] <= WrData_DI[39:32];
        if(BEn_SI[5]) Mem_DP[Addr_DI][47:40] <= WrData_DI[47:40];
        if(BEn_SI[6]) Mem_DP[Addr_DI][55:48] <= WrData_DI[55:48];
        if(BEn_SI[7]) Mem_DP[Addr_DI][63:56] <= WrData_DI[63:56];
      end
      RdData_DN <= Mem_DP[Addr_DI];
    end
  end
  
  
  
  
  generate
    if (OUT_REGS>0) begin : g_outreg
      always_ff @(posedge Clk_CI or negedge Rst_RBI) begin
        if(Rst_RBI == 1'b0)
        begin
          RdData_DP  <= 0;
        end
        else
        begin
          RdData_DP  <= RdData_DN;
        end
      end
    end
  endgenerate 
  
  generate
    if (OUT_REGS==0) begin : g_oureg_byp
      assign RdData_DP  = RdData_DN;
    end
  endgenerate
  assign RdData_DO = RdData_DP;
  
  
  
  
  assert property
    (@(posedge Clk_CI) (longint'(2)**longint'(ADDR_WIDTH) >= longint'(DATA_DEPTH)))
    else $error("depth out of bounds");
  
endmodule 
module axi2mem #(
    parameter int unsigned AXI_ID_WIDTH      = 10,
    parameter int unsigned AXI_ADDR_WIDTH    = 64,
    parameter int unsigned AXI_DATA_WIDTH    = 64,
    parameter int unsigned AXI_USER_WIDTH    = 10
)(
    input logic                         clk_i,    
    input logic                         rst_ni,  
    AXI_BUS.Slave                       slave,
    output logic                        req_o,
    output logic                        we_o,
    output logic [AXI_ADDR_WIDTH-1:0]   addr_o,
    output logic [AXI_DATA_WIDTH/8-1:0] be_o,
    output logic [AXI_DATA_WIDTH-1:0]   data_o,
    input  logic [AXI_DATA_WIDTH-1:0]   data_i
);
    
    
    
    
    typedef enum logic [1:0] { FIXED = 2'b00, INCR = 2'b01, WRAP = 2'b10} axi_burst_t;
    localparam LOG_NR_BYTES = $clog2(AXI_DATA_WIDTH/8);
    typedef struct packed {
        logic [AXI_ID_WIDTH-1:0]   id;
        logic [AXI_ADDR_WIDTH-1:0] addr;
        logic [7:0]                len;
        logic [2:0]                size;
        axi_burst_t                burst;
    } ax_req_t;
    
    enum logic [2:0] { IDLE, READ, WRITE, SEND_B, WAIT_WVALID }  state_d, state_q;
    ax_req_t                   ax_req_d, ax_req_q;
    logic [AXI_ADDR_WIDTH-1:0] req_addr_d, req_addr_q;
    logic [7:0]                cnt_d, cnt_q;
    function automatic logic [AXI_ADDR_WIDTH-1:0] get_wrap_bounadry (input logic [AXI_ADDR_WIDTH-1:0] unaligned_address, input logic [7:0] len);
        logic [AXI_ADDR_WIDTH-1:0] warp_address = '0;
        
        if (len == 4'b1)
            warp_address[AXI_ADDR_WIDTH-1:1+LOG_NR_BYTES] = unaligned_address[AXI_ADDR_WIDTH-1:1+LOG_NR_BYTES];
        else if (len == 4'b11)
            warp_address[AXI_ADDR_WIDTH-1:2+LOG_NR_BYTES] = unaligned_address[AXI_ADDR_WIDTH-1:2+LOG_NR_BYTES];
        else if (len == 4'b111)
            warp_address[AXI_ADDR_WIDTH-1:3+LOG_NR_BYTES] = unaligned_address[AXI_ADDR_WIDTH-3:2+LOG_NR_BYTES];
        else if (len == 4'b1111)
            warp_address[AXI_ADDR_WIDTH-1:4+LOG_NR_BYTES] = unaligned_address[AXI_ADDR_WIDTH-3:4+LOG_NR_BYTES];
        return warp_address;
    endfunction
    logic [AXI_ADDR_WIDTH-1:0] aligned_address;
    logic [AXI_ADDR_WIDTH-1:0] wrap_boundary;
    logic [AXI_ADDR_WIDTH-1:0] upper_wrap_boundary;
    logic [AXI_ADDR_WIDTH-1:0] cons_addr;
    always_comb begin
        
        aligned_address = {ax_req_q.addr[AXI_ADDR_WIDTH-1:LOG_NR_BYTES], {{LOG_NR_BYTES}{1'b0}}};
        wrap_boundary = get_wrap_bounadry(ax_req_q.addr, ax_req_q.len);
        
        upper_wrap_boundary = wrap_boundary + ((ax_req_q.len + 1) << LOG_NR_BYTES);
        
        cons_addr = aligned_address + (cnt_q << LOG_NR_BYTES);
        
        
        state_d    = state_q;
        ax_req_d   = ax_req_q;
        req_addr_d = req_addr_q;
        cnt_d      = cnt_q;
        
        data_o = slave.w_data;
        be_o   = slave.w_strb;
        we_o   = 1'b0;
        req_o  = 1'b0;
        addr_o = '0;
        
        
        slave.aw_ready = 1'b0;
        slave.ar_ready = 1'b0;
        
        slave.r_valid  = 1'b0;
        slave.r_data   = data_i;
        slave.r_resp   = '0;
        slave.r_last   = '0;
        slave.r_id     = ax_req_q.id;
        slave.r_user   = '0;
        
        slave.w_ready  = 1'b0;
        
        slave.b_valid  = 1'b0;
        slave.b_resp   = 1'b0;
        slave.b_id     = 1'b0;
        slave.b_user   = 1'b0;
        case (state_q)
            IDLE: begin
                
                
                
                
                if (slave.ar_valid) begin
                    slave.ar_ready = 1'b1;
                    
                    ax_req_d       = {slave.ar_id, slave.ar_addr, slave.ar_len, slave.ar_size, slave.ar_burst};
                    state_d        = READ;
                    
                    req_o          = 1'b1;
                    addr_o         = slave.ar_addr;
                    
                    req_addr_d     = slave.ar_addr;
                    
                    cnt_d          = 1;
                
                
                
                end else if (slave.aw_valid) begin
                    slave.aw_ready = 1'b1;
                    slave.w_ready  = 1'b1;
                    addr_o         = slave.aw_addr;
                    
                    ax_req_d       = {slave.aw_id, slave.aw_addr, slave.aw_len, slave.aw_size, slave.aw_burst};
                    
                    if (slave.w_valid) begin
                        req_o          = 1'b1;
                        we_o           = 1'b1;
                        state_d        = (slave.w_last) ? SEND_B : WRITE;
                        cnt_d          = 1;
                    
                    end else
                        state_d = WAIT_WVALID;
                end
            end
            
            WAIT_WVALID: begin
                slave.w_ready = 1'b1;
                addr_o = ax_req_q.addr;
                
                if (slave.w_valid) begin
                    req_o          = 1'b1;
                    we_o           = 1'b1;
                    state_d        = (slave.w_last) ? SEND_B : WRITE;
                    cnt_d          = 1;
                end
            end
            READ: begin
                
                req_o  = 1'b1;
                addr_o = req_addr_q;
                
                slave.r_valid = 1'b1;
                slave.r_data  = data_i;
                slave.r_id    = ax_req_q.id;
                slave.r_last  = (cnt_q == ax_req_q.len + 1);
                
                if (slave.r_ready) begin
                    
                    
                    
                    
                    case (ax_req_q.burst)
                        FIXED, INCR: addr_o = cons_addr;
                        WRAP:  begin
                            
                            if (cons_addr == upper_wrap_boundary) begin
                                addr_o = wrap_boundary;
                            
                            end else if (cons_addr > upper_wrap_boundary) begin
                                addr_o = ax_req_q.addr + ((cnt_q - ax_req_q.len) << LOG_NR_BYTES);
                            
                            end else begin
                                addr_o = cons_addr;
                            end
                        end
                    endcase
                    
                    
                    if (slave.r_last) begin
                        state_d = IDLE;
                        
                        req_o = 1'b0;
                    end
                    
                    req_addr_d = addr_o;
                    
                    cnt_d = cnt_q + 1;
                    
                end
            end
            
            WRITE: begin
                slave.w_ready = 1'b1;
                
                if (slave.w_valid) begin
                    req_o         = 1'b1;
                    we_o          = 1'b1;
                    
                    
                    
                    
                    case (ax_req_q.burst)
                        FIXED, INCR: addr_o = cons_addr;
                        WRAP:  begin
                            
                            if (cons_addr == upper_wrap_boundary) begin
                                addr_o = wrap_boundary;
                            
                            end else if (cons_addr > upper_wrap_boundary) begin
                                addr_o = ax_req_q.addr + ((cnt_q - ax_req_q.len) << LOG_NR_BYTES);
                            
                            end else begin
                                addr_o = cons_addr;
                            end
                        end
                    endcase
                    
                    req_addr_d = addr_o;
                    
                    cnt_d = cnt_q + 1;
                    if (slave.w_last)
                        state_d = SEND_B;
                end
            end
            
            SEND_B: begin
                slave.b_valid = 1'b1;
                slave.b_id    = ax_req_q.id;
                if (slave.b_ready)
                    state_d = IDLE;
            end
        endcase
    end
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (~rst_ni) begin
            state_q    <= IDLE;
            ax_req_q  <= '0;
            req_addr_q <= '0;
            cnt_q      <= '0;
        end else begin
            state_q    <= state_d;
            ax_req_q   <= ax_req_d;
            req_addr_q <= req_addr_d;
            cnt_q      <= cnt_d;
        end
    end
endmodule
module pulp_clock_gating
(
    input  logic clk_i,
    input  logic en_i,
    input  logic test_en_i,
    output logic clk_o
);
    logic     clk_en;
    always_latch
    begin
      if (clk_i == 1'b0)
        clk_en <= en_i | test_en_i;
    end
    assign clk_o = clk_i & clk_en;
endmodule
module cluster_clock_inverter
  (
   input  logic clk_i,
   output logic clk_o
   );
   
   assign clk_o = ~clk_i;
   
endmodule
module pulp_clock_mux2
  (
   input  logic clk0_i,
   input  logic clk1_i,
   input  logic clk_sel_i,
   output logic clk_o
   );
   
   always_comb
     begin
	if (clk_sel_i == 1'b0)
	  clk_o = clk0_i;
	else
	  clk_o = clk1_i;
     end
   
endmodule
module pmp #(
    parameter int unsigned PLEN = 34,       
    parameter int unsigned PMP_LEN = 32,    
    parameter int unsigned NR_ENTRIES = 4
) (
    
    input logic [PLEN-1:0] addr_i,
    input riscv::pmp_access_t access_type_i,
    input riscv::priv_lvl_t priv_lvl_i,
    
    input logic [15:0][PMP_LEN-1:0] conf_addr_i,
    input riscv::pmpcfg_t [15:0] conf_i,
    
    output logic allow_o
);
    
    if (NR_ENTRIES > 0) begin : gen_pmp
        logic [NR_ENTRIES-1:0] match;
        for (genvar i = 0; i < NR_ENTRIES; i++) begin
            logic [PMP_LEN-1:0] conf_addr_prev;
            assign conf_addr_prev = (i == 0) ? '0 : conf_addr_i[i-1];
            pmp_entry #(
                .PLEN    ( PLEN    ),
                .PMP_LEN ( PMP_LEN )
            ) i_pmp_entry(
                .addr_i           ( addr_i                         ),
                .conf_addr_i      ( conf_addr_i[i]                 ),
                .conf_addr_prev_i ( conf_addr_prev                 ),
                .conf_addr_mode_i ( conf_i[i].addr_mode            ),
                .match_o          ( match[i]                       )
            );
        end
        always_comb begin
            int i;
            allow_o = 1'b0;
            for (i = 0; i < NR_ENTRIES; i++) begin
                
                
                if (priv_lvl_i != riscv::PRIV_LVL_M || conf_i[i].locked) begin
                    if (match[i]) begin
                        if ((access_type_i & conf_i[i].access_type) != access_type_i) allow_o = 1'b0;
                        else allow_o = 1'b1;
                        break;
                    end
                end
            end
            if (i == NR_ENTRIES) begin 
                
                if (priv_lvl_i == riscv::PRIV_LVL_M) allow_o = 1'b1;
                
                else allow_o = 1'b0;
            end
        end
    end else assign allow_o = 1'b1;
    
    
endmodule
module pmp_entry #(
    parameter int unsigned PLEN = 56,
    parameter int unsigned PMP_LEN = 54
) (
    
    input logic [PLEN-1:0] addr_i,
    
    input logic [PMP_LEN-1:0] conf_addr_i,
    input logic [PMP_LEN-1:0] conf_addr_prev_i,
    input riscv::pmp_addr_mode_t conf_addr_mode_i,
    
    output logic match_o
);
    logic [PLEN-1:0] conf_addr_n;
    logic [$clog2(PLEN)-1:0] trail_ones;
    assign conf_addr_n = ~conf_addr_i;
    lzc #(.WIDTH(PLEN), .MODE(1'b0)) i_lzc(
        .in_i    ( conf_addr_n ),
        .cnt_o   ( trail_ones  ),
        .empty_o (             )
    );
    always_comb begin
        case (conf_addr_mode_i)
            riscv::TOR:     begin
                
                
                if (addr_i >= (conf_addr_prev_i << 2) && addr_i < (conf_addr_i << 2)) begin
                    match_o = 1'b1;
                end else match_o = 1'b0;
                
                
            end
            riscv::NA4, riscv::NAPOT:   begin
                logic [PLEN-1:0] base;
                logic [PLEN-1:0] mask;
                int unsigned size;
                if (conf_addr_mode_i == riscv::NA4) size = 2;
                else begin
                    
                    size = trail_ones+3;
                end
                mask = '1 << size;
                base = (conf_addr_i << 2) & mask;
                match_o = (addr_i & mask) == base ? 1'b1 : 1'b0;
                
                
            end
            riscv::OFF: match_o = 1'b0;
            default:    match_o = 0;
        endcase
    end
endmodule
module axi_adapter #(
  parameter int unsigned DATA_WIDTH            = 256,
  parameter logic        CRITICAL_WORD_FIRST   = 0, 
  parameter int unsigned AXI_ID_WIDTH          = 10,
  parameter int unsigned CACHELINE_BYTE_OFFSET = 8
)(
  input  logic                             clk_i,  
  input  logic                             rst_ni, 
  input  logic                             req_i,
  input  ariane_axi::ad_req_t              type_i,
  output logic                             gnt_o,
  output logic [AXI_ID_WIDTH-1:0]          gnt_id_o,
  input  logic [63:0]                      addr_i,
  input  logic                             we_i,
  input  logic [(DATA_WIDTH/64)-1:0][63:0] wdata_i,
  input  logic [(DATA_WIDTH/64)-1:0][7:0]  be_i,
  input  logic [1:0]                       size_i,
  input  logic [AXI_ID_WIDTH-1:0]          id_i,
  
  output logic                             valid_o,
  output logic [(DATA_WIDTH/64)-1:0][63:0] rdata_o,
  output logic [AXI_ID_WIDTH-1:0]          id_o,
  
  output logic [63:0]                      critical_word_o,
  output logic                             critical_word_valid_o,
  
  output ariane_axi::req_t                 axi_req_o,
  input  ariane_axi::resp_t                axi_resp_i
);
  localparam BURST_SIZE = DATA_WIDTH/64-1;
  localparam ADDR_INDEX = ($clog2(DATA_WIDTH/64) > 0) ? $clog2(DATA_WIDTH/64) : 1;
  enum logic [3:0] {
    IDLE, WAIT_B_VALID, WAIT_AW_READY, WAIT_LAST_W_READY, WAIT_LAST_W_READY_AW_READY, WAIT_AW_READY_BURST,
    WAIT_R_VALID, WAIT_R_VALID_MULTIPLE, COMPLETE_READ
  } state_q, state_d;
  
  logic [ADDR_INDEX-1:0] cnt_d, cnt_q;
  logic [(DATA_WIDTH/64)-1:0][63:0] cache_line_d, cache_line_q;
  
  logic [(DATA_WIDTH/64)-1:0] addr_offset_d, addr_offset_q;
  logic [AXI_ID_WIDTH-1:0]    id_d, id_q;
  logic [ADDR_INDEX-1:0]      index;
  always_comb begin : axi_fsm
    
    axi_req_o.aw_valid  = 1'b0;
    axi_req_o.aw.addr   = addr_i;
    axi_req_o.aw.prot   = 3'b0;
    axi_req_o.aw.region = 4'b0;
    axi_req_o.aw.len    = 8'b0;
    axi_req_o.aw.size   = {1'b0, size_i}; 
    axi_req_o.aw.burst  = axi_pkg::BURST_INCR; 
    axi_req_o.aw.lock   = 1'b0;
    axi_req_o.aw.cache  = 4'b0;
    axi_req_o.aw.qos    = 4'b0;
    axi_req_o.aw.id     = id_i;
    axi_req_o.aw.atop   = '0; 
    axi_req_o.aw.user   = '0;
    axi_req_o.ar_valid  = 1'b0;
    
    
    axi_req_o.ar.addr   = (CRITICAL_WORD_FIRST || type_i == ariane_axi::SINGLE_REQ) ? addr_i : { addr_i[63:CACHELINE_BYTE_OFFSET], {{CACHELINE_BYTE_OFFSET}{1'b0}}};
    axi_req_o.ar.prot   = 3'b0;
    axi_req_o.ar.region = 4'b0;
    axi_req_o.ar.len    = 8'b0;
    axi_req_o.ar.size   = {1'b0, size_i}; 
    axi_req_o.ar.burst  = (CRITICAL_WORD_FIRST ? axi_pkg::BURST_WRAP : axi_pkg::BURST_INCR); 
    axi_req_o.ar.lock   = 1'b0;
    axi_req_o.ar.cache  = 4'b0;
    axi_req_o.ar.qos    = 4'b0;
    axi_req_o.ar.id     = id_i;
    axi_req_o.ar.user   = '0;
    axi_req_o.w_valid   = 1'b0;
    axi_req_o.w.data    = wdata_i[0];
    axi_req_o.w.strb    = be_i[0];
    axi_req_o.w.last    = 1'b0;
    axi_req_o.w.user    = '0;
    axi_req_o.b_ready   = 1'b0;
    axi_req_o.r_ready   = 1'b0;
    gnt_o    = 1'b0;
    gnt_id_o = id_i;
    valid_o  = 1'b0;
    id_o     = axi_resp_i.r.id;
    critical_word_o       = axi_resp_i.r.data;
    critical_word_valid_o = 1'b0;
    rdata_o               = cache_line_q;
    state_d       = state_q;
    cnt_d         = cnt_q;
    cache_line_d  = cache_line_q;
    addr_offset_d = addr_offset_q;
    id_d          = id_q;
    index         = '0;
    case (state_q)
      IDLE: begin
        cnt_d = '0;
        
        if (req_i) begin
          
          
          if (we_i) begin
            
            axi_req_o.aw_valid = 1'b1;
            axi_req_o.w_valid  = 1'b1;
            
            if (type_i == ariane_axi::SINGLE_REQ) begin
              
              axi_req_o.w.last   = 1'b1;
              
              gnt_o = axi_resp_i.aw_ready & axi_resp_i.w_ready;
              case ({axi_resp_i.aw_ready, axi_resp_i.w_ready})
                2'b11: state_d = WAIT_B_VALID;
                2'b01: state_d = WAIT_AW_READY;
                2'b10: state_d = WAIT_LAST_W_READY;
                default: state_d = IDLE;
              endcase
            
            end else begin
              axi_req_o.aw.len = BURST_SIZE; 
              axi_req_o.w.data = wdata_i[0];
              axi_req_o.w.strb = be_i[0];
              if (axi_resp_i.w_ready)
                cnt_d = BURST_SIZE - 1;
              else
                cnt_d = BURST_SIZE;
              case ({axi_resp_i.aw_ready, axi_resp_i.w_ready})
                2'b11: state_d = WAIT_LAST_W_READY;
                2'b01: state_d = WAIT_LAST_W_READY_AW_READY;
                2'b10: state_d = WAIT_LAST_W_READY;
                default:;
              endcase
            end
          
          end else begin
            axi_req_o.ar_valid = 1'b1;
            gnt_o = axi_resp_i.ar_ready;
            if (type_i != ariane_axi::SINGLE_REQ) begin
              axi_req_o.ar.len = BURST_SIZE;
              cnt_d = BURST_SIZE;
            end
            if (axi_resp_i.ar_ready) begin
              state_d = (type_i == ariane_axi::SINGLE_REQ) ? WAIT_R_VALID : WAIT_R_VALID_MULTIPLE;
              addr_offset_d = addr_i[ADDR_INDEX-1+3:3];
            end
          end
        end
      end
      
      WAIT_AW_READY: begin
        axi_req_o.aw_valid = 1'b1;
        if (axi_resp_i.aw_ready) begin
          gnt_o   = 1'b1;
          state_d = WAIT_B_VALID;
        end
      end
      
      WAIT_LAST_W_READY_AW_READY: begin
        axi_req_o.w_valid  = 1'b1;
        axi_req_o.w.last   = (cnt_q == '0);
        if (type_i == ariane_axi::SINGLE_REQ) begin
          axi_req_o.w.data = wdata_i[0];
          axi_req_o.w.strb = be_i[0];
        end else begin
          axi_req_o.w.data = wdata_i[BURST_SIZE-cnt_q];
          axi_req_o.w.strb = be_i[BURST_SIZE-cnt_q];
        end
        axi_req_o.aw_valid = 1'b1;
        
        axi_req_o.aw.len   = BURST_SIZE;
        
        case ({axi_resp_i.aw_ready, axi_resp_i.w_ready})
          
          2'b01: begin
            
            if (cnt_q == 0)
              state_d = WAIT_AW_READY_BURST;
            else 
              cnt_d = cnt_q - 1;
          end
          2'b10: state_d = WAIT_LAST_W_READY;
          2'b11: begin
            
            if (cnt_q == 0) begin
              state_d = WAIT_B_VALID;
              gnt_o   = 1'b1;
            
            end else begin
              state_d = WAIT_LAST_W_READY;
              cnt_d   = cnt_q - 1;
            end
          end
          default:;
         endcase
      end
      
      WAIT_AW_READY_BURST: begin
        axi_req_o.aw_valid = 1'b1;
        axi_req_o.aw.len   = BURST_SIZE;
        if (axi_resp_i.aw_ready) begin
          state_d  = WAIT_B_VALID;
          gnt_o    = 1'b1;
        end
      end
      
      WAIT_LAST_W_READY: begin
        axi_req_o.w_valid = 1'b1;
        if (type_i != ariane_axi::SINGLE_REQ) begin
          axi_req_o.w.data = wdata_i[BURST_SIZE-cnt_q];
          axi_req_o.w.strb = be_i[BURST_SIZE-cnt_q];
        end
        
        if (cnt_q == '0) begin
          axi_req_o.w.last = 1'b1;
          if (axi_resp_i.w_ready) begin
            state_d = WAIT_B_VALID;
            gnt_o   = 1'b1;
          end
        end else if (axi_resp_i.w_ready) begin
          cnt_d = cnt_q - 1;
        end
      end
      
      WAIT_B_VALID: begin
        axi_req_o.b_ready = 1'b1;
        id_o = axi_resp_i.b.id;
        
        if (axi_resp_i.b_valid) begin
          state_d = IDLE;
          valid_o = 1'b1;
        end
      end
      
      WAIT_R_VALID_MULTIPLE, WAIT_R_VALID: begin
        if (CRITICAL_WORD_FIRST)
          index = addr_offset_q + (BURST_SIZE-cnt_q);
        else
          index = BURST_SIZE-cnt_q;
        
        axi_req_o.r_ready = 1'b1;
        
        if (axi_resp_i.r_valid) begin
          if (CRITICAL_WORD_FIRST) begin
            
            if (state_q == WAIT_R_VALID_MULTIPLE && cnt_q == BURST_SIZE) begin
              critical_word_valid_o = 1'b1;
              critical_word_o       = axi_resp_i.r.data;
            end
          end else begin
            
            if (index == addr_offset_q) begin
              critical_word_valid_o = 1'b1;
              critical_word_o       = axi_resp_i.r.data;
            end
          end
          
          if (axi_resp_i.r.last) begin
            id_d    = axi_resp_i.r.id;
            state_d = COMPLETE_READ;
          end
          
          if (state_q == WAIT_R_VALID_MULTIPLE) begin
            cache_line_d[index] = axi_resp_i.r.data;
          end else
            cache_line_d[0] = axi_resp_i.r.data;
          
          cnt_d = cnt_q - 1;
        end
      end
      
      COMPLETE_READ: begin
        valid_o = 1'b1;
        state_d = IDLE;
        id_o    = id_q;
      end
    endcase
  end
  
  
  
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (~rst_ni) begin
      
      state_q       <= IDLE;
      cnt_q         <= '0;
      cache_line_q  <= '0;
      addr_offset_q <= '0;
      id_q          <= '0;
    end else begin
      state_q       <= state_d;
      cnt_q         <= cnt_d;
      cache_line_q  <= cache_line_d;
      addr_offset_q <= addr_offset_d;
      id_q          <= id_d;
    end
  end
endmodule
module alu import ariane_pkg::*;(
    input  logic                     clk_i,          
    input  logic                     rst_ni,         
    input  fu_data_t                 fu_data_i,
    output riscv::xlen_t             result_o,
    output logic                     alu_branch_res_o
);
    riscv::xlen_t operand_a_rev;
    logic [31:0] operand_a_rev32;
    logic [riscv::XLEN:0] operand_b_neg;
    logic [riscv::XLEN+1:0] adder_result_ext_o;
    logic        less;  
    
    generate
      genvar k;
      for(k = 0; k < riscv::XLEN; k++)
        assign operand_a_rev[k] = fu_data_i.operand_a[riscv::XLEN-1-k];
      for (k = 0; k < 32; k++)
        assign operand_a_rev32[k] = fu_data_i.operand_a[31-k];
    endgenerate
    
    
    
    logic        adder_op_b_negate;
    logic        adder_z_flag;
    logic [riscv::XLEN:0] adder_in_a, adder_in_b;
    riscv::xlen_t adder_result;
    always_comb begin
      adder_op_b_negate = 1'b0;
      unique case (fu_data_i.operator)
        
        EQ,  NE,
        SUB, SUBW: adder_op_b_negate = 1'b1;
        default: ;
      endcase
    end
    
    assign adder_in_a    = {fu_data_i.operand_a, 1'b1};
    
    assign operand_b_neg = {fu_data_i.operand_b, 1'b0} ^ {riscv::XLEN+1{adder_op_b_negate}};
    assign adder_in_b    =  operand_b_neg ;
    
    assign adder_result_ext_o = $unsigned(adder_in_a) + $unsigned(adder_in_b);
    assign adder_result       = adder_result_ext_o[riscv::XLEN:1];
    assign adder_z_flag       = ~|adder_result;
    
    always_comb begin : branch_resolve
        
        alu_branch_res_o      = 1'b1;
        case (fu_data_i.operator)
            EQ:       alu_branch_res_o = adder_z_flag;
            NE:       alu_branch_res_o = ~adder_z_flag;
            LTS, LTU: alu_branch_res_o = less;
            GES, GEU: alu_branch_res_o = ~less;
            default:  alu_branch_res_o = 1'b1;
        endcase
    end
    
    
    
    
    logic        shift_left;          
    logic        shift_arithmetic;
    riscv::xlen_t shift_amt;           
    riscv::xlen_t shift_op_a;          
    logic [31:0] shift_op_a32;        
    riscv::xlen_t shift_result;
    logic [31:0] shift_result32;
    logic [riscv::XLEN:0] shift_right_result;
    logic [32:0] shift_right_result32;
    riscv::xlen_t shift_left_result;
    logic [31:0] shift_left_result32;
    assign shift_amt = fu_data_i.operand_b;
    assign shift_left = (fu_data_i.operator == SLL) | (fu_data_i.operator == SLLW);
    assign shift_arithmetic = (fu_data_i.operator == SRA) | (fu_data_i.operator == SRAW);
    
    logic [riscv::XLEN:0] shift_op_a_64;
    logic [32:0] shift_op_a_32;
    
    assign shift_op_a    = shift_left ? operand_a_rev   : fu_data_i.operand_a;
    assign shift_op_a32  = shift_left ? operand_a_rev32 : fu_data_i.operand_a[31:0];
    assign shift_op_a_64 = { shift_arithmetic & shift_op_a[riscv::XLEN-1], shift_op_a};
    assign shift_op_a_32 = { shift_arithmetic & shift_op_a[31], shift_op_a32};
    assign shift_right_result     = $unsigned($signed(shift_op_a_64) >>> shift_amt[5:0]);
    assign shift_right_result32   = $unsigned($signed(shift_op_a_32) >>> shift_amt[4:0]);
    
    genvar j;
    generate
      for(j = 0; j < riscv::XLEN; j++)
        assign shift_left_result[j] = shift_right_result[riscv::XLEN-1-j];
      for(j = 0; j < 32; j++)
        assign shift_left_result32[j] = shift_right_result32[31-j];
    endgenerate
    assign shift_result = shift_left ? shift_left_result : shift_right_result[riscv::XLEN-1:0];
    assign shift_result32 = shift_left ? shift_left_result32 : shift_right_result32[31:0];
    
    
    
    always_comb begin
        logic sgn;
        sgn = 1'b0;
        if ((fu_data_i.operator == SLTS) ||
            (fu_data_i.operator == LTS)  ||
            (fu_data_i.operator == GES))
            sgn = 1'b1;
        less = ($signed({sgn & fu_data_i.operand_a[riscv::XLEN-1], fu_data_i.operand_a})  <  $signed({sgn & fu_data_i.operand_b[riscv::XLEN-1], fu_data_i.operand_b}));
    end
    
    
    
    always_comb begin
        result_o   = '0;
        unique case (fu_data_i.operator)
            
            ANDL:  result_o = fu_data_i.operand_a & fu_data_i.operand_b;
            ORL:   result_o = fu_data_i.operand_a | fu_data_i.operand_b;
            XORL:  result_o = fu_data_i.operand_a ^ fu_data_i.operand_b;
            
            ADD, SUB: result_o = adder_result;
            
            ADDW, SUBW: result_o = {{riscv::XLEN-32{adder_result[31]}}, adder_result[31:0]};
            
            SLL,
            SRL, SRA: result_o = (riscv::XLEN == 64) ? shift_result : shift_result32;
            
            SLLW,
            SRLW, SRAW: result_o = {{riscv::XLEN-32{shift_result32[31]}}, shift_result32[31:0]};
            
            SLTS,  SLTU: result_o = {{riscv::XLEN-1{1'b0}}, less};
            default: ; 
        endcase
    end
endmodule
module fpu_wrap import ariane_pkg::*; (
  input  logic                     clk_i,
  input  logic                     rst_ni,
  input  logic                     flush_i,
  input  logic                     fpu_valid_i,
  output logic                     fpu_ready_o,
  input  fu_data_t                 fu_data_i,
  input  logic [1:0]               fpu_fmt_i,
  input  logic [2:0]               fpu_rm_i,
  input  logic [2:0]               fpu_frm_i,
  input  logic [6:0]               fpu_prec_i,
  output logic [TRANS_ID_BITS-1:0] fpu_trans_id_o,
  output logic [FLEN-1:0]          result_o,
  output logic                     fpu_valid_o,
  output exception_t               fpu_exception_o
);
  
  
  enum logic {READY, STALL} state_q, state_d;
  if (FP_PRESENT) begin : fpu_gen
    logic [FLEN-1:0] operand_a_i;
    logic [FLEN-1:0] operand_b_i;
    logic [FLEN-1:0] operand_c_i;
    assign operand_a_i = fu_data_i.operand_a[FLEN-1:0];
    assign operand_b_i = fu_data_i.operand_b[FLEN-1:0];
    assign operand_c_i = fu_data_i.imm[FLEN-1:0];
    
    
    
    localparam OPBITS  =  fpnew_pkg::OP_BITS;
    localparam FMTBITS =  $clog2(fpnew_pkg::NUM_FP_FORMATS);
    localparam IFMTBITS = $clog2(fpnew_pkg::NUM_INT_FORMATS);
    
    localparam fpnew_pkg::fpu_features_t FPU_FEATURES = '{
      Width:         riscv::XLEN, 
      EnableVectors: ariane_pkg::XFVEC,
      EnableNanBox:  1'b1,
      FpFmtMask:     {RVF, RVD, XF16, XF8, XF16ALT},
      IntFmtMask:    {XFVEC && XF8, XFVEC && (XF16 || XF16ALT), 1'b1, 1'b1}
    };
    
    localparam fpnew_pkg::fpu_implementation_t FPU_IMPLEMENTATION = '{
      PipeRegs:  '{
                 '{LAT_COMP_FP32, LAT_COMP_FP64, LAT_COMP_FP16, LAT_COMP_FP8, LAT_COMP_FP16ALT}, 
                 '{default: LAT_DIVSQRT}, 
                 '{default: LAT_NONCOMP}, 
                 '{default: LAT_CONV}},   
      UnitTypes: '{'{default: fpnew_pkg::PARALLEL}, 
                   '{default: fpnew_pkg::MERGED},   
                   '{default: fpnew_pkg::PARALLEL}, 
                   '{default: fpnew_pkg::MERGED}},  
      PipeConfig: fpnew_pkg::DISTRIBUTED
    };
    
    
    
    logic [FLEN-1:0]     operand_a_d,  operand_a_q,  operand_a;
    logic [FLEN-1:0]     operand_b_d,  operand_b_q,  operand_b;
    logic [FLEN-1:0]     operand_c_d,  operand_c_q,  operand_c;
    logic [OPBITS-1:0]   fpu_op_d,     fpu_op_q,     fpu_op;
    logic                fpu_op_mod_d, fpu_op_mod_q, fpu_op_mod;
    logic [FMTBITS-1:0]  fpu_srcfmt_d, fpu_srcfmt_q, fpu_srcfmt;
    logic [FMTBITS-1:0]  fpu_dstfmt_d, fpu_dstfmt_q, fpu_dstfmt;
    logic [IFMTBITS-1:0] fpu_ifmt_d,   fpu_ifmt_q,   fpu_ifmt;
    logic [2:0]          fpu_rm_d,     fpu_rm_q,     fpu_rm;
    logic                fpu_vec_op_d, fpu_vec_op_q, fpu_vec_op;
    logic [TRANS_ID_BITS-1:0] fpu_tag_d, fpu_tag_q, fpu_tag;
    logic fpu_in_ready, fpu_in_valid;
    logic fpu_out_ready, fpu_out_valid;
    logic [4:0] fpu_status;
    
    logic hold_inputs;
    logic use_hold;
    
    
    
    always_comb begin : input_translation
      automatic logic vec_replication; 
      automatic logic replicate_c;     
      automatic logic check_ah;        
      
      operand_a_d         = operand_a_i;
      operand_b_d         = operand_b_i; 
      operand_c_d         = operand_c_i; 
      fpu_op_d            = fpnew_pkg::SGNJ; 
      fpu_op_mod_d        = 1'b0;
      fpu_dstfmt_d        = fpnew_pkg::FP32;
      fpu_ifmt_d          = fpnew_pkg::INT32;
      fpu_rm_d            = fpu_rm_i;
      fpu_vec_op_d        = fu_data_i.fu == FPU_VEC;
      fpu_tag_d           = fu_data_i.trans_id;
      vec_replication     = fpu_rm_i[0]; 
      replicate_c         = 1'b0;
      check_ah            = 1'b0; 
      
      if (!(fpu_rm_i inside {[3'b000:3'b100]}))
        fpu_rm_d = fpu_frm_i;
      
      if (fpu_vec_op_d)
        fpu_rm_d = fpu_frm_i;
      
      unique case (fpu_fmt_i)
        
        2'b00: fpu_dstfmt_d = fpnew_pkg::FP32;
        
        2'b01: fpu_dstfmt_d = fpu_vec_op_d ? fpnew_pkg::FP16ALT : fpnew_pkg::FP64;
        
        2'b10: begin
           if (!fpu_vec_op_d && fpu_rm_i==3'b101)
             fpu_dstfmt_d = fpnew_pkg::FP16ALT;
           else
             fpu_dstfmt_d = fpnew_pkg::FP16;
        end
        
        default: fpu_dstfmt_d = fpnew_pkg::FP8;
      endcase
      
      fpu_srcfmt_d = fpu_dstfmt_d;
      
      unique case (fu_data_i.operator)
        
        FADD: begin
          fpu_op_d    = fpnew_pkg::ADD;
          replicate_c = 1'b1; 
        end
        
        FSUB: begin
          fpu_op_d     = fpnew_pkg::ADD;
          fpu_op_mod_d = 1'b1;
          replicate_c  = 1'b1; 
        end
        
        FMUL: fpu_op_d = fpnew_pkg::MUL;
        
        FDIV: fpu_op_d = fpnew_pkg::DIV;
        
        FMIN_MAX: begin
          fpu_op_d = fpnew_pkg::MINMAX;
          fpu_rm_d = {1'b0, fpu_rm_i[1:0]}; 
          check_ah = 1'b1; 
        end
        
        FSQRT: fpu_op_d = fpnew_pkg::SQRT;
        
        FMADD: fpu_op_d = fpnew_pkg::FMADD;
        
        FMSUB: begin
          fpu_op_d     = fpnew_pkg::FMADD;
          fpu_op_mod_d = 1'b1;
        end
        
        FNMSUB: fpu_op_d = fpnew_pkg::FNMSUB;
        
        FNMADD: begin
          fpu_op_d     = fpnew_pkg::FNMSUB;
          fpu_op_mod_d = 1'b1;
        end
        
        FCVT_F2I: begin
          fpu_op_d     = fpnew_pkg::F2I;
          
          if (fpu_vec_op_d) begin
            fpu_op_mod_d      = fpu_rm_i[0];
            vec_replication = 1'b0; 
            unique case (fpu_fmt_i)
              2'b00: fpu_ifmt_d = fpnew_pkg::INT32;
              2'b01,
              2'b10: fpu_ifmt_d = fpnew_pkg::INT16;
              2'b11: fpu_ifmt_d = fpnew_pkg::INT8;
            endcase
          
          end else begin
            fpu_op_mod_d = operand_c_i[0];
            if (operand_c_i[1])
              fpu_ifmt_d = fpnew_pkg::INT64;
            else
              fpu_ifmt_d = fpnew_pkg::INT32;
          end
        end
        
        FCVT_I2F: begin
          fpu_op_d = fpnew_pkg::I2F;
          
          if (fpu_vec_op_d) begin
            fpu_op_mod_d      = fpu_rm_i[0];
            vec_replication = 1'b0; 
            unique case (fpu_fmt_i)
              2'b00: fpu_ifmt_d = fpnew_pkg::INT32;
              2'b01,
              2'b10: fpu_ifmt_d = fpnew_pkg::INT16;
              2'b11: fpu_ifmt_d = fpnew_pkg::INT8;
            endcase
          
          end else begin
            fpu_op_mod_d = operand_c_i[0];
            if (operand_c_i[1])
              fpu_ifmt_d = fpnew_pkg::INT64;
            else
              fpu_ifmt_d = fpnew_pkg::INT32;
          end
        end
        
        FCVT_F2F: begin
          fpu_op_d = fpnew_pkg::F2F;
          
          if (fpu_vec_op_d) begin
            vec_replication = 1'b0; 
            unique case (operand_c_i[1:0])
              2'b00: fpu_srcfmt_d = fpnew_pkg::FP32;
              2'b01: fpu_srcfmt_d = fpnew_pkg::FP16ALT;
              2'b10: fpu_srcfmt_d = fpnew_pkg::FP16;
              2'b11: fpu_srcfmt_d = fpnew_pkg::FP8;
            endcase
          
          end else begin
            unique case (operand_c_i[2:0])
              3'b000: fpu_srcfmt_d = fpnew_pkg::FP32;
              3'b001: fpu_srcfmt_d = fpnew_pkg::FP64;
              3'b010: fpu_srcfmt_d = fpnew_pkg::FP16;
              3'b110: fpu_srcfmt_d = fpnew_pkg::FP16ALT;
              3'b011: fpu_srcfmt_d = fpnew_pkg::FP8;
            endcase
          end
        end
        
        FSGNJ: begin
          fpu_op_d = fpnew_pkg::SGNJ;
          fpu_rm_d = {1'b0, fpu_rm_i[1:0]}; 
          check_ah = 1'b1; 
        end
        
        FMV_F2X: begin
          fpu_op_d          = fpnew_pkg::SGNJ;
          fpu_rm_d          = 3'b011; 
          fpu_op_mod_d      = 1'b1; 
          check_ah          = 1'b1; 
          vec_replication   = 1'b0; 
        end
        
        FMV_X2F: begin
          fpu_op_d          = fpnew_pkg::SGNJ;
          fpu_rm_d          = 3'b011; 
          check_ah          = 1'b1; 
          vec_replication   = 1'b0; 
        end
        
        FCMP: begin
          fpu_op_d = fpnew_pkg::CMP;
          fpu_rm_d = {1'b0, fpu_rm_i[1:0]}; 
          check_ah = 1'b1; 
        end
        
        FCLASS: begin
          fpu_op_d = fpnew_pkg::CLASSIFY;
          fpu_rm_d = {1'b0, fpu_rm_i[1:0]}; 
          check_ah = 1'b1; 
        end
        
        VFMIN: begin
          fpu_op_d = fpnew_pkg::MINMAX;
          fpu_rm_d = 3'b000; 
        end
        
        VFMAX: begin
          fpu_op_d = fpnew_pkg::MINMAX;
          fpu_rm_d = 3'b001; 
        end
        
        VFSGNJ: begin
          fpu_op_d = fpnew_pkg::SGNJ;
          fpu_rm_d = 3'b000; 
        end
        
        VFSGNJN: begin
          fpu_op_d = fpnew_pkg::SGNJ;
          fpu_rm_d = 3'b001; 
        end
        
        VFSGNJX: begin
          fpu_op_d = fpnew_pkg::SGNJ;
          fpu_rm_d = 3'b010; 
        end
        
        VFEQ: begin
          fpu_op_d = fpnew_pkg::CMP;
          fpu_rm_d = 3'b010; 
        end
        
        VFNE: begin
          fpu_op_d     = fpnew_pkg::CMP;
          fpu_op_mod_d = 1'b1;   
          fpu_rm_d     = 3'b010; 
          end
        
        VFLT: begin
          fpu_op_d = fpnew_pkg::CMP;
          fpu_rm_d = 3'b001; 
        end
        
        VFGE: begin
          fpu_op_d     = fpnew_pkg::CMP;
          fpu_op_mod_d = 1'b1;   
          fpu_rm_d     = 3'b001; 
        end
        
        VFLE: begin
          fpu_op_d = fpnew_pkg::CMP;
          fpu_rm_d = 3'b000; 
        end
        
        VFGT: begin
          fpu_op_d     = fpnew_pkg::CMP;
          fpu_op_mod_d = 1'b1;   
          fpu_rm_d     = 3'b000; 
        end
        
        VFCPKAB_S: begin
          fpu_op_d        = fpnew_pkg::CPKAB;
          fpu_op_mod_d    = fpu_rm_i[0]; 
          vec_replication = 1'b0; 
          fpu_srcfmt_d    = fpnew_pkg::FP32; 
        end
        
        VFCPKCD_S: begin
          fpu_op_d        = fpnew_pkg::CPKCD;
          fpu_op_mod_d    = fpu_rm_i[0]; 
          vec_replication = 1'b0; 
          fpu_srcfmt_d    = fpnew_pkg::FP32; 
        end
        
        VFCPKAB_D: begin
          fpu_op_d        = fpnew_pkg::CPKAB;
          fpu_op_mod_d    = fpu_rm_i[0]; 
          vec_replication = 1'b0; 
          fpu_srcfmt_d    = fpnew_pkg::FP64; 
        end
        
        VFCPKCD_D: begin
          fpu_op_d        = fpnew_pkg::CPKCD;
          fpu_op_mod_d    = fpu_rm_i[0]; 
          vec_replication = 1'b0; 
          fpu_srcfmt_d    = fpnew_pkg::FP64; 
        end
        
        default: ; 
      endcase
      
      if (!fpu_vec_op_d && check_ah)
        if (fpu_rm_i[2])
          fpu_dstfmt_d = fpnew_pkg::FP16ALT;
      
      if (fpu_vec_op_d && vec_replication) begin
        if (replicate_c) begin
          unique case (fpu_dstfmt_d)
            fpnew_pkg::FP32:    operand_c_d = RVD ? {2{operand_c_i[31:0]}} : operand_c_i;
            fpnew_pkg::FP16,
            fpnew_pkg::FP16ALT: operand_c_d = RVD ? {4{operand_c_i[15:0]}} : {2{operand_c_i[15:0]}};
            fpnew_pkg::FP8:     operand_c_d = RVD ? {8{operand_c_i[7:0]}}  : {4{operand_c_i[7:0]}};
          endcase 
        end else begin
          unique case (fpu_dstfmt_d)
            fpnew_pkg::FP32:    operand_b_d = RVD ? {2{operand_b_i[31:0]}} : operand_b_i;
            fpnew_pkg::FP16,
            fpnew_pkg::FP16ALT: operand_b_d = RVD ? {4{operand_b_i[15:0]}} : {2{operand_b_i[15:0]}};
            fpnew_pkg::FP8:     operand_b_d = RVD ? {8{operand_b_i[7:0]}}  : {4{operand_b_i[7:0]}};
          endcase 
        end
      end
    end
    
    
    
    always_comb begin : p_inputFSM
      
      fpu_ready_o  = 1'b0;
      fpu_in_valid = 1'b0;
      hold_inputs = 1'b0;    
      use_hold    = 1'b0;    
      state_d     = state_q; 
      
      unique case (state_q)
        
        READY: begin
          fpu_ready_o  = 1'b1;        
          fpu_in_valid = fpu_valid_i; 
          
          if (fpu_valid_i & ~fpu_in_ready) begin
            fpu_ready_o = 1'b0;  
            hold_inputs = 1'b1;  
            state_d     = STALL; 
          end
        end
        
        STALL: begin
          fpu_in_valid = 1'b1; 
          use_hold     = 1'b1; 
          
          if (fpu_in_ready) begin
            fpu_ready_o = 1'b1;  
            state_d     = READY; 
          end
        end
        
        default: ;
      endcase
      
      if (flush_i) begin
        state_d = READY;
      end
    end
    
    always_ff @(posedge clk_i or negedge rst_ni) begin : fp_hold_reg
      if(~rst_ni) begin
        state_q       <= READY;
        operand_a_q   <= '0;
        operand_b_q   <= '0;
        operand_c_q   <= '0;
        fpu_op_q      <= '0;
        fpu_op_mod_q  <= '0;
        fpu_srcfmt_q  <= '0;
        fpu_dstfmt_q  <= '0;
        fpu_ifmt_q    <= '0;
        fpu_rm_q      <= '0;
        fpu_vec_op_q  <= '0;
        fpu_tag_q     <= '0;
      end else begin
        state_q       <= state_d;
        
        if (hold_inputs) begin
          operand_a_q   <= operand_a_d;
          operand_b_q   <= operand_b_d;
          operand_c_q   <= operand_c_d;
          fpu_op_q      <= fpu_op_d;
          fpu_op_mod_q  <= fpu_op_mod_d;
          fpu_srcfmt_q  <= fpu_srcfmt_d;
          fpu_dstfmt_q  <= fpu_dstfmt_d;
          fpu_ifmt_q    <= fpu_ifmt_d;
          fpu_rm_q      <= fpu_rm_d;
          fpu_vec_op_q  <= fpu_vec_op_d;
          fpu_tag_q     <= fpu_tag_d;
        end
      end
    end
    
    assign operand_a  = use_hold ? operand_a_q  : operand_a_d;
    assign operand_b  = use_hold ? operand_b_q  : operand_b_d;
    assign operand_c  = use_hold ? operand_c_q  : operand_c_d;
    assign fpu_op     = use_hold ? fpu_op_q     : fpu_op_d;
    assign fpu_op_mod = use_hold ? fpu_op_mod_q : fpu_op_mod_d;
    assign fpu_srcfmt = use_hold ? fpu_srcfmt_q : fpu_srcfmt_d;
    assign fpu_dstfmt = use_hold ? fpu_dstfmt_q : fpu_dstfmt_d;
    assign fpu_ifmt   = use_hold ? fpu_ifmt_q   : fpu_ifmt_d;
    assign fpu_rm     = use_hold ? fpu_rm_q     : fpu_rm_d;
    assign fpu_vec_op = use_hold ? fpu_vec_op_q : fpu_vec_op_d;
    assign fpu_tag    = use_hold ? fpu_tag_q    : fpu_tag_d;
    
    logic [2:0][FLEN-1:0] fpu_operands;
    assign fpu_operands[0] = operand_a;
    assign fpu_operands[1] = operand_b;
    assign fpu_operands[2] = operand_c;
    
    
    
    fpnew_top #(
      .Features       ( FPU_FEATURES              ),
      .Implementation ( FPU_IMPLEMENTATION        ),
      .TagType        ( logic [TRANS_ID_BITS-1:0] )
    ) i_fpnew_bulk (
      .clk_i,
      .rst_ni,
      .operands_i     ( fpu_operands                        ),
      .rnd_mode_i     ( fpnew_pkg::roundmode_e'(fpu_rm)     ),
      .op_i           ( fpnew_pkg::operation_e'(fpu_op)     ),
      .op_mod_i       ( fpu_op_mod                          ),
      .src_fmt_i      ( fpnew_pkg::fp_format_e'(fpu_srcfmt) ),
      .dst_fmt_i      ( fpnew_pkg::fp_format_e'(fpu_dstfmt) ),
      .int_fmt_i      ( fpnew_pkg::int_format_e'(fpu_ifmt)  ),
      .vectorial_op_i ( fpu_vec_op                          ),
      .tag_i          ( fpu_tag                             ),
      .in_valid_i     ( fpu_in_valid                        ),
      .in_ready_o     ( fpu_in_ready                        ),
      .flush_i,
      .result_o,
      .status_o       ( fpu_status                          ),
      .tag_o          ( fpu_trans_id_o                      ),
      .out_valid_o    ( fpu_out_valid                       ),
      .out_ready_i    ( fpu_out_ready                       ),
      .busy_o         (                         )
    );
    
    assign fpu_exception_o.cause = {59'h0, fpu_status};
    assign fpu_exception_o.valid = 1'b0;
    
    assign fpu_out_ready = 1'b1;
    
    assign fpu_valid_o = fpu_out_valid;
  end
endmodule
module ariane import ariane_pkg::*; #(
  parameter ariane_pkg::ariane_cfg_t ArianeCfg     = ariane_pkg::ArianeDefaultConfig
) (
  input  logic                         clk_i,
  input  logic                         rst_ni,
  
  input  logic [riscv::VLEN-1:0]       boot_addr_i,  
  input  logic [riscv::XLEN-1:0]       hart_id_i,    
  
  input  logic [1:0]                   irq_i,        
  input  logic                         ipi_i,        
  
  input  logic                         time_irq_i,   
  input  logic                         debug_req_i,  
  
  output wt_cache_pkg::l15_req_t       l15_req_o,
  input  wt_cache_pkg::l15_rtrn_t      l15_rtrn_i
);
  
  
  
  
  riscv::priv_lvl_t           priv_lvl;
  exception_t                 ex_commit; 
  bp_resolve_t                resolved_branch;
  logic [riscv::VLEN-1:0]     pc_commit;
  logic                       eret;
  logic [NR_COMMIT_PORTS-1:0] commit_ack;
  
  
  
  logic [riscv::VLEN-1:0]     trap_vector_base_commit_pcgen;
  logic [riscv::VLEN-1:0]     epc_commit_pcgen;
  
  
  
  fetch_entry_t             fetch_entry_if_id;
  logic                     fetch_valid_if_id;
  logic                     fetch_ready_id_if;
  
  
  
  scoreboard_entry_t        issue_entry_id_issue;
  logic                     issue_entry_valid_id_issue;
  logic                     is_ctrl_fow_id_issue;
  logic                     issue_instr_issue_id;
  
  
  
   logic [riscv::VLEN-1:0] rs1_forwarding_id_ex; 
   logic [riscv::VLEN-1:0] rs2_forwarding_id_ex; 
  fu_data_t                 fu_data_id_ex;
  logic [riscv::VLEN-1:0]   pc_id_ex;
  logic                     is_compressed_instr_id_ex;
  
  logic                     flu_ready_ex_id;
  logic [TRANS_ID_BITS-1:0] flu_trans_id_ex_id;
  logic                     flu_valid_ex_id;
  riscv::xlen_t             flu_result_ex_id;
  exception_t               flu_exception_ex_id;
  
  logic                     alu_valid_id_ex;
  
  logic                     branch_valid_id_ex;
  branchpredict_sbe_t       branch_predict_id_ex;
  logic                     resolve_branch_ex_id;
  
  logic                     lsu_valid_id_ex;
  logic                     lsu_ready_ex_id;
  logic [TRANS_ID_BITS-1:0] load_trans_id_ex_id;
  riscv::xlen_t             load_result_ex_id;
  logic                     load_valid_ex_id;
  exception_t               load_exception_ex_id;
  riscv::xlen_t             store_result_ex_id;
  logic [TRANS_ID_BITS-1:0] store_trans_id_ex_id;
  logic                     store_valid_ex_id;
  exception_t               store_exception_ex_id;
  
  logic                     mult_valid_id_ex;
  
  logic                     fpu_ready_ex_id;
  logic                     fpu_valid_id_ex;
  logic [1:0]               fpu_fmt_id_ex;
  logic [2:0]               fpu_rm_id_ex;
  logic [TRANS_ID_BITS-1:0] fpu_trans_id_ex_id;
  riscv::xlen_t             fpu_result_ex_id;
  logic                     fpu_valid_ex_id;
  exception_t               fpu_exception_ex_id;
  
  logic                     csr_valid_id_ex;
  
  
  
  
  logic                     csr_commit_commit_ex;
  logic                     dirty_fp_state;
  
  logic                     lsu_commit_commit_ex;
  logic                     lsu_commit_ready_ex_commit;
  logic [TRANS_ID_BITS-1:0] lsu_commit_trans_id;
  logic                     no_st_pending_ex;
  logic                     no_st_pending_commit;
  logic                     amo_valid_commit;
  
  
  
  scoreboard_entry_t [NR_COMMIT_PORTS-1:0] commit_instr_id_commit;
  
  
  
  logic [NR_COMMIT_PORTS-1:0][4:0]  waddr_commit_id;
  logic [NR_COMMIT_PORTS-1:0][riscv::XLEN-1:0] wdata_commit_id;
  logic [NR_COMMIT_PORTS-1:0]       we_gpr_commit_id;
  logic [NR_COMMIT_PORTS-1:0]       we_fpr_commit_id;
  
  
  
  logic [4:0]               fflags_csr_commit;
  riscv::xs_t               fs;
  logic [2:0]               frm_csr_id_issue_ex;
  logic [6:0]               fprec_csr_ex;
  logic                     enable_translation_csr_ex;
  logic                     en_ld_st_translation_csr_ex;
  riscv::priv_lvl_t         ld_st_priv_lvl_csr_ex;
  logic                     sum_csr_ex;
  logic                     mxr_csr_ex;
  logic [riscv::PPNW-1:0]   satp_ppn_csr_ex;
  logic [ASID_WIDTH-1:0]    asid_csr_ex;
  logic [11:0]              csr_addr_ex_csr;
  fu_op                     csr_op_commit_csr;
  riscv::xlen_t             csr_wdata_commit_csr;
  riscv::xlen_t             csr_rdata_csr_commit;
  exception_t               csr_exception_csr_commit;
  logic                     tvm_csr_id;
  logic                     tw_csr_id;
  logic                     tsr_csr_id;
  irq_ctrl_t                irq_ctrl_csr_id;
  logic                     dcache_en_csr_nbdcache;
  logic                     csr_write_fflags_commit_cs;
  logic                     icache_en_csr;
  logic                     debug_mode;
  logic                     single_step_csr_commit;
  riscv::pmpcfg_t [15:0]    pmpcfg;
  logic [15:0][riscv::PLEN-3:0] pmpaddr;
  
  
  
  logic [4:0]               addr_csr_perf;
  riscv::xlen_t             data_csr_perf, data_perf_csr;
  logic                     we_csr_perf;
  logic                     icache_flush_ctrl_cache;
  logic                     itlb_miss_ex_perf;
  logic                     dtlb_miss_ex_perf;
  logic                     dcache_miss_cache_perf;
  logic                     icache_miss_cache_perf;
  
  
  
  logic                     set_pc_ctrl_pcgen;
  logic                     flush_csr_ctrl;
  logic                     flush_unissued_instr_ctrl_id;
  logic                     flush_ctrl_if;
  logic                     flush_ctrl_id;
  logic                     flush_ctrl_ex;
  logic                     flush_ctrl_bp;
  logic                     flush_tlb_ctrl_ex;
  logic                     fence_i_commit_controller;
  logic                     fence_commit_controller;
  logic                     sfence_vma_commit_controller;
  logic                     halt_ctrl;
  logic                     halt_csr_ctrl;
  logic                     dcache_flush_ctrl_cache;
  logic                     dcache_flush_ack_cache_ctrl;
  logic                     set_debug_pc;
  logic                     flush_commit;
  icache_areq_i_t           icache_areq_ex_cache;
  icache_areq_o_t           icache_areq_cache_ex;
  icache_dreq_i_t           icache_dreq_if_cache;
  icache_dreq_o_t           icache_dreq_cache_if;
  amo_req_t                 amo_req;
  amo_resp_t                amo_resp;
  logic                     sb_full;
  
  
  
  dcache_req_i_t [2:0]      dcache_req_ports_ex_cache;
  dcache_req_o_t [2:0]      dcache_req_ports_cache_ex;
  logic                     dcache_commit_wbuffer_empty;
  logic                     dcache_commit_wbuffer_not_ni;
  
  
  
  frontend #(
    .ArianeCfg ( ArianeCfg )
  ) i_frontend (
    .flush_i             ( flush_ctrl_if                 ), 
    .flush_bp_i          ( 1'b0                          ),
    .debug_mode_i        ( debug_mode                    ),
    .boot_addr_i         ( boot_addr_i[riscv::VLEN-1:0]  ),
    .icache_dreq_i       ( icache_dreq_cache_if          ),
    .icache_dreq_o       ( icache_dreq_if_cache          ),
    .resolved_branch_i   ( resolved_branch               ),
    .pc_commit_i         ( pc_commit                     ),
    .set_pc_commit_i     ( set_pc_ctrl_pcgen             ),
    .set_debug_pc_i      ( set_debug_pc                  ),
    .epc_i               ( epc_commit_pcgen              ),
    .eret_i              ( eret                          ),
    .trap_vector_base_i  ( trap_vector_base_commit_pcgen ),
    .ex_valid_i          ( ex_commit.valid               ),
    .fetch_entry_o       ( fetch_entry_if_id             ),
    .fetch_entry_valid_o ( fetch_valid_if_id             ),
    .fetch_entry_ready_i ( fetch_ready_id_if             ),
    .*
  );
  
  
  
  id_stage id_stage_i (
    .clk_i,
    .rst_ni,
    .flush_i                    ( flush_ctrl_if              ),
    .debug_req_i,
    .fetch_entry_i              ( fetch_entry_if_id          ),
    .fetch_entry_valid_i        ( fetch_valid_if_id          ),
    .fetch_entry_ready_o        ( fetch_ready_id_if          ),
    .issue_entry_o              ( issue_entry_id_issue       ),
    .issue_entry_valid_o        ( issue_entry_valid_id_issue ),
    .is_ctrl_flow_o             ( is_ctrl_fow_id_issue       ),
    .issue_instr_ack_i          ( issue_instr_issue_id       ),
    .priv_lvl_i                 ( priv_lvl                   ),
    .fs_i                       ( fs                         ),
    .frm_i                      ( frm_csr_id_issue_ex        ),
    .irq_i                      ( irq_i                      ),
    .irq_ctrl_i                 ( irq_ctrl_csr_id            ),
    .debug_mode_i               ( debug_mode                 ),
    .tvm_i                      ( tvm_csr_id                 ),
    .tw_i                       ( tw_csr_id                  ),
    .tsr_i                      ( tsr_csr_id                 )
  );
  
  
  
  issue_stage #(
    .NR_ENTRIES                 ( NR_SB_ENTRIES                ),
    .NR_WB_PORTS                ( NR_WB_PORTS                  ),
    .NR_COMMIT_PORTS            ( NR_COMMIT_PORTS              )
  ) issue_stage_i (
    .clk_i,
    .rst_ni,
    .sb_full_o                  ( sb_full                      ),
    .flush_unissued_instr_i     ( flush_unissued_instr_ctrl_id ),
    .flush_i                    ( flush_ctrl_id                ),
    
    .decoded_instr_i            ( issue_entry_id_issue         ),
    .decoded_instr_valid_i      ( issue_entry_valid_id_issue   ),
    .is_ctrl_flow_i             ( is_ctrl_fow_id_issue         ),
    .decoded_instr_ack_o        ( issue_instr_issue_id         ),
    
    .rs1_forwarding_o           ( rs1_forwarding_id_ex         ),
    .rs2_forwarding_o           ( rs2_forwarding_id_ex         ),
    .fu_data_o                  ( fu_data_id_ex                ),
    .pc_o                       ( pc_id_ex                     ),
    .is_compressed_instr_o      ( is_compressed_instr_id_ex    ),
    
    .flu_ready_i                ( flu_ready_ex_id              ),
    
    .alu_valid_o                ( alu_valid_id_ex              ),
    
    .branch_valid_o             ( branch_valid_id_ex           ), 
    .branch_predict_o           ( branch_predict_id_ex         ), 
    .resolve_branch_i           ( resolve_branch_ex_id         ), 
    
    .lsu_ready_i                ( lsu_ready_ex_id              ),
    .lsu_valid_o                ( lsu_valid_id_ex              ),
    
    .mult_valid_o               ( mult_valid_id_ex             ),
    
    .fpu_ready_i                ( fpu_ready_ex_id              ),
    .fpu_valid_o                ( fpu_valid_id_ex              ),
    .fpu_fmt_o                  ( fpu_fmt_id_ex                ),
    .fpu_rm_o                   ( fpu_rm_id_ex                 ),
    
    .csr_valid_o                ( csr_valid_id_ex              ),
    
    .resolved_branch_i          ( resolved_branch              ),
    .trans_id_i                 ( {flu_trans_id_ex_id,  load_trans_id_ex_id,  store_trans_id_ex_id,   fpu_trans_id_ex_id }),
    .wbdata_i                   ( {flu_result_ex_id,    load_result_ex_id,    store_result_ex_id,       fpu_result_ex_id }),
    .ex_ex_i                    ( {flu_exception_ex_id, load_exception_ex_id, store_exception_ex_id, fpu_exception_ex_id }),
    .wt_valid_i                 ( {flu_valid_ex_id,     load_valid_ex_id,     store_valid_ex_id,         fpu_valid_ex_id }),
    .waddr_i                    ( waddr_commit_id              ),
    .wdata_i                    ( wdata_commit_id              ),
    .we_gpr_i                   ( we_gpr_commit_id             ),
    .we_fpr_i                   ( we_fpr_commit_id             ),
    .commit_instr_o             ( commit_instr_id_commit       ),
    .commit_ack_i               ( commit_ack                   ),
    .*
  );
  
  
  
  ex_stage #(
    .ASID_WIDTH ( ASID_WIDTH ),
    .ArianeCfg  ( ArianeCfg  )
  ) ex_stage_i (
    .clk_i                  ( clk_i                       ),
    .rst_ni                 ( rst_ni                      ),
    .debug_mode_i           ( debug_mode                  ),
    .flush_i                ( flush_ctrl_ex               ),
    .rs1_forwarding_i       ( rs1_forwarding_id_ex        ),
    .rs2_forwarding_i       ( rs2_forwarding_id_ex        ),
    .fu_data_i              ( fu_data_id_ex               ),
    .pc_i                   ( pc_id_ex                    ),
    .is_compressed_instr_i  ( is_compressed_instr_id_ex   ),
    
    .flu_result_o           ( flu_result_ex_id            ),
    .flu_trans_id_o         ( flu_trans_id_ex_id          ),
    .flu_valid_o            ( flu_valid_ex_id             ),
    .flu_exception_o        ( flu_exception_ex_id         ),
    .flu_ready_o            ( flu_ready_ex_id             ),
    
    .alu_valid_i            ( alu_valid_id_ex             ),
    
    .branch_valid_i         ( branch_valid_id_ex          ),
    .branch_predict_i       ( branch_predict_id_ex        ), 
    .resolved_branch_o      ( resolved_branch             ),
    .resolve_branch_o       ( resolve_branch_ex_id        ),
    
    .csr_valid_i            ( csr_valid_id_ex             ),
    .csr_addr_o             ( csr_addr_ex_csr             ),
    .csr_commit_i           ( csr_commit_commit_ex        ), 
    
    .mult_valid_i           ( mult_valid_id_ex            ),
    
    .lsu_ready_o            ( lsu_ready_ex_id             ),
    .lsu_valid_i            ( lsu_valid_id_ex             ),
    .load_result_o          ( load_result_ex_id           ),
    .load_trans_id_o        ( load_trans_id_ex_id         ),
    .load_valid_o           ( load_valid_ex_id            ),
    .load_exception_o       ( load_exception_ex_id        ),
    .store_result_o         ( store_result_ex_id          ),
    .store_trans_id_o       ( store_trans_id_ex_id        ),
    .store_valid_o          ( store_valid_ex_id           ),
    .store_exception_o      ( store_exception_ex_id       ),
    .lsu_commit_i           ( lsu_commit_commit_ex        ), 
    .lsu_commit_ready_o     ( lsu_commit_ready_ex_commit  ), 
    .commit_tran_id_i       ( lsu_commit_trans_id         ), 
    .no_st_pending_o        ( no_st_pending_ex            ),
    
    .fpu_ready_o            ( fpu_ready_ex_id             ),
    .fpu_valid_i            ( fpu_valid_id_ex             ),
    .fpu_fmt_i              ( fpu_fmt_id_ex               ),
    .fpu_rm_i               ( fpu_rm_id_ex                ),
    .fpu_frm_i              ( frm_csr_id_issue_ex         ),
    .fpu_prec_i             ( fprec_csr_ex                ),
    .fpu_trans_id_o         ( fpu_trans_id_ex_id          ),
    .fpu_result_o           ( fpu_result_ex_id            ),
    .fpu_valid_o            ( fpu_valid_ex_id             ),
    .fpu_exception_o        ( fpu_exception_ex_id         ),
    .amo_valid_commit_i     ( amo_valid_commit            ),
    .amo_req_o              ( amo_req                     ),
    .amo_resp_i             ( amo_resp                    ),
    
    .itlb_miss_o            ( itlb_miss_ex_perf           ),
    .dtlb_miss_o            ( dtlb_miss_ex_perf           ),
    
    .enable_translation_i   ( enable_translation_csr_ex   ), 
    .en_ld_st_translation_i ( en_ld_st_translation_csr_ex ),
    .flush_tlb_i            ( flush_tlb_ctrl_ex           ),
    .priv_lvl_i             ( priv_lvl                    ), 
    .ld_st_priv_lvl_i       ( ld_st_priv_lvl_csr_ex       ), 
    .sum_i                  ( sum_csr_ex                  ), 
    .mxr_i                  ( mxr_csr_ex                  ), 
    .satp_ppn_i             ( satp_ppn_csr_ex             ), 
    .asid_i                 ( asid_csr_ex                 ), 
    .icache_areq_i          ( icache_areq_cache_ex        ),
    .icache_areq_o          ( icache_areq_ex_cache        ),
    
    .dcache_req_ports_i     ( dcache_req_ports_cache_ex   ),
    .dcache_req_ports_o     ( dcache_req_ports_ex_cache   ),
    .dcache_wbuffer_empty_i ( dcache_commit_wbuffer_empty ),
    .dcache_wbuffer_not_ni_i ( dcache_commit_wbuffer_not_ni ),
    
    .pmpcfg_i               ( pmpcfg                      ),
    .pmpaddr_i              ( pmpaddr                     )
  );
  
  
  
  
  
  assign no_st_pending_commit = no_st_pending_ex & dcache_commit_wbuffer_empty;
  commit_stage #(
    .NR_COMMIT_PORTS ( NR_COMMIT_PORTS )
  ) commit_stage_i (
    .clk_i,
    .rst_ni,
    .halt_i                 ( halt_ctrl                     ),
    .flush_dcache_i         ( dcache_flush_ctrl_cache       ),
    .exception_o            ( ex_commit                     ),
    .dirty_fp_state_o       ( dirty_fp_state                ),
    .single_step_i          ( single_step_csr_commit        ),
    .commit_instr_i         ( commit_instr_id_commit        ),
    .commit_ack_o           ( commit_ack                    ),
    .no_st_pending_i        ( no_st_pending_commit          ),
    .waddr_o                ( waddr_commit_id               ),
    .wdata_o                ( wdata_commit_id               ),
    .we_gpr_o               ( we_gpr_commit_id              ),
    .we_fpr_o               ( we_fpr_commit_id              ),
    .commit_lsu_o           ( lsu_commit_commit_ex          ),
    .commit_lsu_ready_i     ( lsu_commit_ready_ex_commit    ),
    .commit_tran_id_o       ( lsu_commit_trans_id           ),
    .amo_valid_commit_o     ( amo_valid_commit              ),
    .amo_resp_i             ( amo_resp                      ),
    .commit_csr_o           ( csr_commit_commit_ex          ),
    .pc_o                   ( pc_commit                     ),
    .csr_op_o               ( csr_op_commit_csr             ),
    .csr_wdata_o            ( csr_wdata_commit_csr          ),
    .csr_rdata_i            ( csr_rdata_csr_commit          ),
    .csr_write_fflags_o     ( csr_write_fflags_commit_cs    ),
    .csr_exception_i        ( csr_exception_csr_commit      ),
    .fence_i_o              ( fence_i_commit_controller     ),
    .fence_o                ( fence_commit_controller       ),
    .sfence_vma_o           ( sfence_vma_commit_controller  ),
    .flush_commit_o         ( flush_commit                  ),
    .*
  );
  
  
  
  csr_regfile #(
    .AsidWidth              ( ASID_WIDTH                    ),
    .DmBaseAddress          ( ArianeCfg.DmBaseAddress       ),
    .NrCommitPorts          ( NR_COMMIT_PORTS               ),
    .NrPMPEntries           ( ArianeCfg.NrPMPEntries        )
  ) csr_regfile_i (
    .flush_o                ( flush_csr_ctrl                ),
    .halt_csr_o             ( halt_csr_ctrl                 ),
    .commit_instr_i         ( commit_instr_id_commit        ),
    .commit_ack_i           ( commit_ack                    ),
    .boot_addr_i            ( boot_addr_i[riscv::VLEN-1:0]  ),
    .hart_id_i              ( hart_id_i[riscv::XLEN-1:0]    ),
    .ex_i                   ( ex_commit                     ),
    .csr_op_i               ( csr_op_commit_csr             ),
    .csr_write_fflags_i     ( csr_write_fflags_commit_cs    ),
    .dirty_fp_state_i       ( dirty_fp_state                ),
    .csr_addr_i             ( csr_addr_ex_csr               ),
    .csr_wdata_i            ( csr_wdata_commit_csr          ),
    .csr_rdata_o            ( csr_rdata_csr_commit          ),
    .pc_i                   ( pc_commit                     ),
    .csr_exception_o        ( csr_exception_csr_commit      ),
    .epc_o                  ( epc_commit_pcgen              ),
    .eret_o                 ( eret                          ),
    .set_debug_pc_o         ( set_debug_pc                  ),
    .trap_vector_base_o     ( trap_vector_base_commit_pcgen ),
    .priv_lvl_o             ( priv_lvl                      ),
    .fs_o                   ( fs                            ),
    .fflags_o               ( fflags_csr_commit             ),
    .frm_o                  ( frm_csr_id_issue_ex           ),
    .fprec_o                ( fprec_csr_ex                  ),
    .irq_ctrl_o             ( irq_ctrl_csr_id               ),
    .ld_st_priv_lvl_o       ( ld_st_priv_lvl_csr_ex         ),
    .en_translation_o       ( enable_translation_csr_ex     ),
    .en_ld_st_translation_o ( en_ld_st_translation_csr_ex   ),
    .sum_o                  ( sum_csr_ex                    ),
    .mxr_o                  ( mxr_csr_ex                    ),
    .satp_ppn_o             ( satp_ppn_csr_ex               ),
    .asid_o                 ( asid_csr_ex                   ),
    .tvm_o                  ( tvm_csr_id                    ),
    .tw_o                   ( tw_csr_id                     ),
    .tsr_o                  ( tsr_csr_id                    ),
    .debug_mode_o           ( debug_mode                    ),
    .single_step_o          ( single_step_csr_commit        ),
    .dcache_en_o            ( dcache_en_csr_nbdcache        ),
    .icache_en_o            ( icache_en_csr                 ),
    .perf_addr_o            ( addr_csr_perf                 ),
    .perf_data_o            ( data_csr_perf                 ),
    .perf_data_i            ( data_perf_csr                 ),
    .perf_we_o              ( we_csr_perf                   ),
    .pmpcfg_o               ( pmpcfg                        ),
    .pmpaddr_o              ( pmpaddr                       ),
    .debug_req_i,
    .ipi_i,
    .irq_i,
    .time_irq_i,
    .*
  );
  
  
  
  perf_counters i_perf_counters (
    .clk_i             ( clk_i                  ),
    .rst_ni            ( rst_ni                 ),
    .debug_mode_i      ( debug_mode             ),
    .addr_i            ( addr_csr_perf          ),
    .we_i              ( we_csr_perf            ),
    .data_i            ( data_csr_perf          ),
    .data_o            ( data_perf_csr          ),
    .commit_instr_i    ( commit_instr_id_commit ),
    .commit_ack_i      ( commit_ack             ),
    .l1_icache_miss_i  ( icache_miss_cache_perf ),
    .l1_dcache_miss_i  ( dcache_miss_cache_perf ),
    .itlb_miss_i       ( itlb_miss_ex_perf      ),
    .dtlb_miss_i       ( dtlb_miss_ex_perf      ),
    .sb_full_i         ( sb_full                ),
    .if_empty_i        ( ~fetch_valid_if_id     ),
    .ex_i              ( ex_commit              ),
    .eret_i            ( eret                   ),
    .resolved_branch_i ( resolved_branch        )
  );
  
  
  
  controller controller_i (
    
    .set_pc_commit_o        ( set_pc_ctrl_pcgen             ),
    .flush_unissued_instr_o ( flush_unissued_instr_ctrl_id  ),
    .flush_if_o             ( flush_ctrl_if                 ),
    .flush_id_o             ( flush_ctrl_id                 ),
    .flush_ex_o             ( flush_ctrl_ex                 ),
    .flush_bp_o             ( flush_ctrl_bp                 ),
    .flush_tlb_o            ( flush_tlb_ctrl_ex             ),
    .flush_dcache_o         ( dcache_flush_ctrl_cache       ),
    .flush_dcache_ack_i     ( dcache_flush_ack_cache_ctrl   ),
    .halt_csr_i             ( halt_csr_ctrl                 ),
    .halt_o                 ( halt_ctrl                     ),
    
    .eret_i                 ( eret                          ),
    .ex_valid_i             ( ex_commit.valid               ),
    .set_debug_pc_i         ( set_debug_pc                  ),
    .flush_csr_i            ( flush_csr_ctrl                ),
    .resolved_branch_i      ( resolved_branch               ),
    .fence_i_i              ( fence_i_commit_controller     ),
    .fence_i                ( fence_commit_controller       ),
    .sfence_vma_i           ( sfence_vma_commit_controller  ),
    .flush_commit_i         ( flush_commit                  ),
    .flush_icache_o         ( icache_flush_ctrl_cache       ),
    .*
  );
  
  
  
  std_cache_subsystem #(
    
    
    
    .ArianeCfg             ( ArianeCfg                   )
  ) i_cache_subsystem (
    
    .clk_i                 ( clk_i                       ),
    .rst_ni                ( rst_ni                      ),
    .priv_lvl_i            ( priv_lvl                    ),
    
    .icache_en_i           ( icache_en_csr               ),
    .icache_flush_i        ( icache_flush_ctrl_cache     ),
    .icache_miss_o         ( icache_miss_cache_perf      ),
    .icache_areq_i         ( icache_areq_ex_cache        ),
    .icache_areq_o         ( icache_areq_cache_ex        ),
    .icache_dreq_i         ( icache_dreq_if_cache        ),
    .icache_dreq_o         ( icache_dreq_cache_if        ),
    
    .dcache_enable_i       ( dcache_en_csr_nbdcache      ),
    .dcache_flush_i        ( dcache_flush_ctrl_cache     ),
    .dcache_flush_ack_o    ( dcache_flush_ack_cache_ctrl ),
    
    .amo_req_i             ( amo_req                     ),
    .amo_resp_o            ( amo_resp                    ),
    .dcache_miss_o         ( dcache_miss_cache_perf      ),
    
    .wbuffer_empty_o       ( dcache_commit_wbuffer_empty ),
    
    .dcache_req_ports_i    ( dcache_req_ports_ex_cache   ),
    .dcache_req_ports_o    ( dcache_req_ports_cache_ex   ),
    
    .axi_req_o             ( axi_req_o                   ),
    .axi_resp_i            ( axi_resp_i                  )
  );
  assign dcache_commit_wbuffer_not_ni = 1'b1;
  
  
  
  
  
  
  
  
  
  
  
  
  localparam PC_QUEUE_DEPTH = 16;
  logic        piton_pc_vld;
  logic [riscv::VLEN-1:0] piton_pc;
  logic [NR_COMMIT_PORTS-1:0][riscv::VLEN-1:0] pc_data;
  logic [NR_COMMIT_PORTS-1:0] pc_pop, pc_empty;
  for (genvar i = 0; i < NR_COMMIT_PORTS; i++) begin : gen_pc_fifo
    fifo_v3 #(
      .DATA_WIDTH(64),
      .DEPTH(PC_QUEUE_DEPTH))
    i_pc_fifo (
      .clk_i      ( clk_i                                               ),
      .rst_ni     ( rst_ni                                              ),
      .flush_i    ( '0                                                  ),
      .testmode_i ( '0                                                  ),
      .full_o     (                                                     ),
      .empty_o    ( pc_empty[i]                                         ),
      .usage_o    (                                                     ),
      .data_i     ( commit_instr_id_commit[i].pc                        ),
      .push_i     ( commit_ack[i] & ~commit_instr_id_commit[i].ex.valid ),
      .data_o     ( pc_data[i]                                          ),
      .pop_i      ( pc_pop[i]                                           )
    );
  end
  rr_arb_tree #(
    .NumIn(NR_COMMIT_PORTS),
    .DataWidth(64))
  i_rr_arb_tree (
    .clk_i   ( clk_i        ),
    .rst_ni  ( rst_ni       ),
    .flush_i ( '0           ),
    .rr_i    ( '0           ),
    .req_i   ( ~pc_empty    ),
    .gnt_o   ( pc_pop       ),
    .data_i  ( pc_data      ),
    .gnt_i   ( piton_pc_vld ),
    .req_o   ( piton_pc_vld ),
    .data_o  ( piton_pc     ),
    .idx_o   (              )
  );
 
  int f;
  logic [63:0] cycles;
  initial begin
    f = $fopen("trace_hart_00.dasm", "w");
  end
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (~rst_ni) begin
      cycles <= 0;
    end else begin
      byte mode = "";
      if (debug_mode) mode = "D";
      else begin
        case (priv_lvl)
        riscv::PRIV_LVL_M: mode = "M";
        riscv::PRIV_LVL_S: mode = "S";
        riscv::PRIV_LVL_U: mode = "U";
        endcase
      end
      for (int i = 0; i < NR_COMMIT_PORTS; i++) begin
        if (commit_ack[i] && !commit_instr_id_commit[i].ex.valid) begin
          $fwrite(f, "%d 0x%0h %s (0x%h) DASM(%h)\n", cycles, commit_instr_id_commit[i].pc, mode, commit_instr_id_commit[i].ex.tval[31:0], commit_instr_id_commit[i].ex.tval[31:0]);
        end else if (commit_ack[i] && commit_instr_id_commit[i].ex.valid) begin
          if (commit_instr_id_commit[i].ex.cause == 2) begin
            $fwrite(f, "Exception Cause: Illegal Instructions, DASM(%h) PC=%h\n", commit_instr_id_commit[i].ex.tval[31:0], commit_instr_id_commit[i].pc);
          end else begin
            if (debug_mode) begin
              $fwrite(f, "%d 0x%0h %s (0x%h) DASM(%h)\n", cycles, commit_instr_id_commit[i].pc, mode, commit_instr_id_commit[i].ex.tval[31:0], commit_instr_id_commit[i].ex.tval[31:0]);
            end else begin
              $fwrite(f, "Exception Cause: %5d, DASM(%h) PC=%h\n", commit_instr_id_commit[i].ex.cause, commit_instr_id_commit[i].ex.tval[31:0], commit_instr_id_commit[i].pc);
            end
          end
        end
      end
        cycles <= cycles + 1;
    end
  end
  final begin
    $fclose(f);
  end
 
endmodule 
module branch_unit (
    input  logic                      clk_i,
    input  logic                      rst_ni,
    input  logic                      debug_mode_i,
    input  ariane_pkg::fu_data_t      fu_data_i,
    input  logic [riscv::VLEN-1:0]    pc_i,                   
    input  logic                      is_compressed_instr_i,
    input  logic                      fu_valid_i,             
    input  logic                      branch_valid_i,
    input  logic                      branch_comp_res_i,      
    output logic [riscv::VLEN-1:0]    branch_result_o,
    input  ariane_pkg::branchpredict_sbe_t        branch_predict_i,       
    output ariane_pkg::bp_resolve_t               resolved_branch_o,      
    output logic                      resolve_branch_o,       
                                                              
    output ariane_pkg::exception_t    branch_exception_o      
);
    logic [riscv::VLEN-1:0] target_address;
    logic [riscv::VLEN-1:0] next_pc;
   
    always_comb begin : mispredict_handler
        
        automatic logic [riscv::VLEN-1:0] jump_base;
        
        jump_base = (fu_data_i.operator == ariane_pkg::JALR) ? fu_data_i.operand_a[riscv::VLEN-1:0] : pc_i;
        target_address                   = {riscv::VLEN{1'b0}};
        resolve_branch_o                 = 1'b0;
        resolved_branch_o.target_address = {riscv::VLEN{1'b0}};
        resolved_branch_o.is_taken       = 1'b0;
        resolved_branch_o.valid          = branch_valid_i;
        resolved_branch_o.is_mispredict  = 1'b0;
        resolved_branch_o.cf_type        = branch_predict_i.cf;
        
        
        next_pc                          = pc_i + ((is_compressed_instr_i) ? {{riscv::VLEN-2{1'b0}}, 2'h2} : {{riscv::VLEN-3{1'b0}}, 3'h4});
        
        target_address                   = $unsigned($signed(jump_base) + $signed(fu_data_i.imm[riscv::VLEN-1:0]));
        
        if (fu_data_i.operator == ariane_pkg::JALR) target_address[0] = 1'b0;
        
        branch_result_o = next_pc;
        resolved_branch_o.pc = pc_i;
        
        
        
        if (branch_valid_i) begin
            
            resolved_branch_o.target_address = (branch_comp_res_i) ? target_address : next_pc;
            resolved_branch_o.is_taken = branch_comp_res_i;
            
            if (ariane_pkg::op_is_branch(fu_data_i.operator) && branch_comp_res_i != (branch_predict_i.cf == ariane_pkg::Branch)) begin
                
                
                resolved_branch_o.is_mispredict  = 1'b1;
                resolved_branch_o.cf_type = ariane_pkg::Branch;
            end
            if (fu_data_i.operator == ariane_pkg::JALR
                
                && (branch_predict_i.cf == ariane_pkg::NoCF || target_address != branch_predict_i.predict_address)) begin
                resolved_branch_o.is_mispredict  = 1'b1;
                
                if (branch_predict_i.cf != ariane_pkg::Return) resolved_branch_o.cf_type = ariane_pkg::JumpR;
            end
            
            resolve_branch_o = 1'b1;
        end
    end
    
    
    always_comb begin : exception_handling
        branch_exception_o.cause = riscv::INSTR_ADDR_MISALIGNED;
        branch_exception_o.valid = 1'b0;
        branch_exception_o.tval  = {{riscv::XLEN-riscv::VLEN{pc_i[riscv::VLEN-1]}}, pc_i};
        
        if (branch_valid_i && target_address[0] != 1'b0) branch_exception_o.valid = 1'b1;
    end
endmodule
module compressed_decoder
(
    input  logic [31:0] instr_i,
    output logic [31:0] instr_o,
    output logic        illegal_instr_o,
    output logic        is_compressed_o
);
    
    
    
    always_comb begin
        illegal_instr_o = 1'b0;
        instr_o         = '0;
        is_compressed_o = 1'b1;
        instr_o         = instr_i;
        
        
        unique case (instr_i[1:0])
            
            riscv::OpcodeC0: begin
                unique case (instr_i[15:13])
                    riscv::OpcodeC0Addi4spn: begin
                        
                        instr_o = {2'b0, instr_i[10:7], instr_i[12:11], instr_i[5], instr_i[6], 2'b00, 5'h02, 3'b000, 2'b01, instr_i[4:2], riscv::OpcodeOpImm};
                        if (instr_i[12:5] == 8'b0)  illegal_instr_o = 1'b1;
                    end
                    riscv::OpcodeC0Fld: begin
                        
                        
                        instr_o = {4'b0, instr_i[6:5], instr_i[12:10], 3'b000, 2'b01, instr_i[9:7], 3'b011, 2'b01, instr_i[4:2], riscv::OpcodeLoadFp};
                    end
                    riscv::OpcodeC0Lw: begin
                        
                        instr_o = {5'b0, instr_i[5], instr_i[12:10], instr_i[6], 2'b00, 2'b01, instr_i[9:7], 3'b010, 2'b01, instr_i[4:2], riscv::OpcodeLoad};
                    end
                    riscv::OpcodeC0Ld: begin
                        
                        
                        instr_o = {4'b0, instr_i[6:5], instr_i[12:10], 3'b000, 2'b01, instr_i[9:7], 3'b011, 2'b01, instr_i[4:2], riscv::OpcodeLoad};
                    end
                    riscv::OpcodeC0Fsd: begin
                        
                        instr_o = {4'b0, instr_i[6:5], instr_i[12], 2'b01, instr_i[4:2], 2'b01, instr_i[9:7], 3'b011, instr_i[11:10], 3'b000, riscv::OpcodeStoreFp};
                    end
                    riscv::OpcodeC0Sw: begin
                        
                        instr_o = {5'b0, instr_i[5], instr_i[12], 2'b01, instr_i[4:2], 2'b01, instr_i[9:7], 3'b010, instr_i[11:10], instr_i[6], 2'b00, riscv::OpcodeStore};
                    end
                    riscv::OpcodeC0Sd: begin
                        
                        instr_o = {4'b0, instr_i[6:5], instr_i[12], 2'b01, instr_i[4:2], 2'b01, instr_i[9:7], 3'b011, instr_i[11:10], 3'b000, riscv::OpcodeStore};
                    end
                    default: begin
                        illegal_instr_o = 1'b1;
                    end
              endcase
            end
            
            riscv::OpcodeC1: begin
                unique case (instr_i[15:13])
                    riscv::OpcodeC1Addi: begin
                        
                        
                        instr_o = {{6 {instr_i[12]}}, instr_i[12], instr_i[6:2], instr_i[11:7], 3'b0, instr_i[11:7], riscv::OpcodeOpImm};
                    end
                    
                    riscv::OpcodeC1Addiw: begin 
                        if (riscv::XLEN == 64) begin
                            
                            if (instr_i[11:7] != 5'h0) begin 
                                instr_o = {{6 {instr_i[12]}}, instr_i[12], instr_i[6:2], instr_i[11:7], 3'b0, instr_i[11:7], riscv::OpcodeOpImm32};
                            end else begin
                                illegal_instr_o = 1'b1;
                            end
                        end else begin
                            
                            instr_o = {instr_i[12], instr_i[8], instr_i[10:9], instr_i[6], instr_i[7], instr_i[2], instr_i[11], instr_i[5:3], {9 {instr_i[12]}}, 5'b1, riscv::OpcodeJal};
             
                        end
                    end
                    riscv::OpcodeC1Li: begin
                        
                        instr_o = {{6 {instr_i[12]}}, instr_i[12], instr_i[6:2], 5'b0, 3'b0, instr_i[11:7], riscv::OpcodeOpImm};
                    end
                    riscv::OpcodeC1LuiAddi16sp: begin
                        
                        instr_o = {{15 {instr_i[12]}}, instr_i[6:2], instr_i[11:7], riscv::OpcodeLui};
                        if (instr_i[11:7] == 5'h02) begin
                            
                            instr_o = {{3 {instr_i[12]}}, instr_i[4:3], instr_i[5], instr_i[2], instr_i[6], 4'b0, 5'h02, 3'b000, 5'h02, riscv::OpcodeOpImm};
                        end
                        if ({instr_i[12], instr_i[6:2]} == 6'b0) illegal_instr_o = 1'b1;
                    end
                    riscv::OpcodeC1MiscAlu: begin
                        unique case (instr_i[11:10])
                            2'b00,
                            2'b01: begin
                                
                                
                                instr_o = {1'b0, instr_i[10], 4'b0, instr_i[12], instr_i[6:2], 2'b01, instr_i[9:7], 3'b101, 2'b01, instr_i[9:7], riscv::OpcodeOpImm};
                            end
                            2'b10: begin
                                
                                instr_o = {{6 {instr_i[12]}}, instr_i[12], instr_i[6:2], 2'b01, instr_i[9:7], 3'b111, 2'b01, instr_i[9:7], riscv::OpcodeOpImm};
                            end
                            2'b11: begin
                                unique case ({instr_i[12], instr_i[6:5]})
                                    3'b000: begin
                                        
                                        instr_o = {2'b01, 5'b0, 2'b01, instr_i[4:2], 2'b01, instr_i[9:7], 3'b000, 2'b01, instr_i[9:7], riscv::OpcodeOp};
                                    end
                                    3'b001: begin
                                        
                                        instr_o = {7'b0, 2'b01, instr_i[4:2], 2'b01, instr_i[9:7], 3'b100, 2'b01, instr_i[9:7], riscv::OpcodeOp};
                                    end
                                    3'b010: begin
                                        
                                        instr_o = {7'b0, 2'b01, instr_i[4:2], 2'b01, instr_i[9:7], 3'b110, 2'b01, instr_i[9:7], riscv::OpcodeOp};
                                    end
                                    3'b011: begin
                                        
                                        instr_o = {7'b0, 2'b01, instr_i[4:2], 2'b01, instr_i[9:7], 3'b111, 2'b01, instr_i[9:7], riscv::OpcodeOp};
                                    end
                                    3'b100: begin
                                        
                                        instr_o = {2'b01, 5'b0, 2'b01, instr_i[4:2], 2'b01, instr_i[9:7], 3'b000, 2'b01, instr_i[9:7], riscv::OpcodeOp32};
                                    end
                                    3'b101: begin
                                        
                                        instr_o = {2'b00, 5'b0, 2'b01, instr_i[4:2], 2'b01, instr_i[9:7], 3'b000, 2'b01, instr_i[9:7], riscv::OpcodeOp32};
                                    end
                                    3'b110,
                                    3'b111: begin
                                        
                                        
                                        illegal_instr_o = 1'b1;
                                        instr_o = {16'b0, instr_i};
                                    end
                                endcase
                            end
                        endcase
                    end
                    riscv::OpcodeC1J: begin
                        
                        instr_o = {instr_i[12], instr_i[8], instr_i[10:9], instr_i[6], instr_i[7], instr_i[2], instr_i[11], instr_i[5:3], {9 {instr_i[12]}}, 4'b0, ~instr_i[15], riscv::OpcodeJal};
                    end
                    riscv::OpcodeC1Beqz, riscv::OpcodeC1Bnez: begin
                        
                        
                        instr_o = {{4 {instr_i[12]}}, instr_i[6:5], instr_i[2], 5'b0, 2'b01, instr_i[9:7], 2'b00, instr_i[13], instr_i[11:10], instr_i[4:3], instr_i[12], riscv::OpcodeBranch};
                    end
                endcase
            end
            
            riscv::OpcodeC2: begin
                unique case (instr_i[15:13])
                    riscv::OpcodeC2Slli: begin
                        
                        instr_o = {6'b0, instr_i[12], instr_i[6:2], instr_i[11:7], 3'b001, instr_i[11:7], riscv::OpcodeOpImm};
                    end
                    riscv::OpcodeC2Fldsp: begin
                        
                        instr_o = {3'b0, instr_i[4:2], instr_i[12], instr_i[6:5], 3'b000, 5'h02, 3'b011, instr_i[11:7], riscv::OpcodeLoadFp};
                    end
                    riscv::OpcodeC2Lwsp: begin
                        
                        instr_o = {4'b0, instr_i[3:2], instr_i[12], instr_i[6:4], 2'b00, 5'h02, 3'b010, instr_i[11:7], riscv::OpcodeLoad};
                        if (instr_i[11:7] == 5'b0)  illegal_instr_o = 1'b1;
                    end
                    riscv::OpcodeC2Ldsp: begin
                        
                        instr_o = {3'b0, instr_i[4:2], instr_i[12], instr_i[6:5], 3'b000, 5'h02, 3'b011, instr_i[11:7], riscv::OpcodeLoad};
                        if (instr_i[11:7] == 5'b0)  illegal_instr_o = 1'b1;
                    end
                    riscv::OpcodeC2JalrMvAdd: begin
                        if (instr_i[12] == 1'b0) begin
                            
                            instr_o = {7'b0, instr_i[6:2], 5'b0, 3'b0, instr_i[11:7], riscv::OpcodeOp};
                            if (instr_i[6:2] == 5'b0) begin
                                
                                instr_o = {12'b0, instr_i[11:7], 3'b0, 5'b0, riscv::OpcodeJalr};
                                
                                illegal_instr_o = (instr_i[11:7] != '0) ? 1'b0 : 1'b1;
                            end
                        end else begin
                            
                            instr_o = {7'b0, instr_i[6:2], instr_i[11:7], 3'b0, instr_i[11:7], riscv::OpcodeOp};
                            if (instr_i[11:7] == 5'b0 && instr_i[6:2] == 5'b0) begin
                                
                                instr_o = {32'h00_10_00_73};
                            end else if (instr_i[11:7] != 5'b0 && instr_i[6:2] == 5'b0) begin
                                
                                instr_o = {12'b0, instr_i[11:7], 3'b000, 5'b00001, riscv::OpcodeJalr};
                            end
                        end
                    end
                    riscv::OpcodeC2Fsdsp: begin
                        
                        instr_o = {3'b0, instr_i[9:7], instr_i[12], instr_i[6:2], 5'h02, 3'b011, instr_i[11:10], 3'b000, riscv::OpcodeStoreFp};
                    end
                    riscv::OpcodeC2Swsp: begin
                        
                        instr_o = {4'b0, instr_i[8:7], instr_i[12], instr_i[6:2], 5'h02, 3'b010, instr_i[11:9], 2'b00, riscv::OpcodeStore};
                    end
                    riscv::OpcodeC2Sdsp: begin
                        
                        instr_o = {3'b0, instr_i[9:7], instr_i[12], instr_i[6:2], 5'h02, 3'b011, instr_i[11:10], 3'b000, riscv::OpcodeStore};
                    end
                    default: begin
                        illegal_instr_o = 1'b1;
                    end
                endcase
            end
            
            default: is_compressed_o = 1'b0;
        endcase
        
        if (illegal_instr_o && is_compressed_o) begin
            instr_o = instr_i;
        end
    end
endmodule
module controller import ariane_pkg::*; (
    input  logic            clk_i,
    input  logic            rst_ni,
    output logic            set_pc_commit_o,        
    output logic            flush_if_o,             
    output logic            flush_unissued_instr_o, 
    output logic            flush_id_o,             
    output logic            flush_ex_o,             
    output logic            flush_bp_o,             
    output logic            flush_icache_o,         
    output logic            flush_dcache_o,         
    input  logic            flush_dcache_ack_i,     
    output logic            flush_tlb_o,            
    input  logic            halt_csr_i,             
    output logic            halt_o,                 
    input  logic            eret_i,                 
    input  logic            ex_valid_i,             
    input  logic            set_debug_pc_i,         
    input  bp_resolve_t     resolved_branch_i,      
    input  logic            flush_csr_i,            
    input  logic            fence_i_i,              
    input  logic            fence_i,                
    input  logic            sfence_vma_i,           
    input  logic            flush_commit_i          
);
    
    logic fence_active_d, fence_active_q;
    logic flush_dcache;
    
    
    
    always_comb begin : flush_ctrl
        fence_active_d         = fence_active_q;
        set_pc_commit_o        = 1'b0;
        flush_if_o             = 1'b0;
        flush_unissued_instr_o = 1'b0;
        flush_id_o             = 1'b0;
        flush_ex_o             = 1'b0;
        flush_dcache           = 1'b0;
        flush_icache_o         = 1'b0;
        flush_tlb_o            = 1'b0;
        flush_bp_o             = 1'b0;
        
        
        
        
        if (resolved_branch_i.is_mispredict) begin
            
            flush_unissued_instr_o = 1'b1;
            
            flush_if_o             = 1'b1;
        end
        
        
        
        if (fence_i) begin
            
            set_pc_commit_o        = 1'b1;
            flush_if_o             = 1'b1;
            flush_unissued_instr_o = 1'b1;
            flush_id_o             = 1'b1;
            flush_ex_o             = 1'b1;
            flush_dcache           = 1'b1;
            fence_active_d         = 1'b1;
        end
        
        
        
        if (fence_i_i) begin
            set_pc_commit_o        = 1'b1;
            flush_if_o             = 1'b1;
            flush_unissued_instr_o = 1'b1;
            flush_id_o             = 1'b1;
            flush_ex_o             = 1'b1;
            flush_icache_o         = 1'b1;
            flush_dcache           = 1'b1;
            fence_active_d         = 1'b1;
        end
        
        if (flush_dcache_ack_i && fence_active_q) begin
            fence_active_d = 1'b0;
        
        end else if (fence_active_q) begin
            flush_dcache = 1'b1;
        end
        
        
        
        if (sfence_vma_i) begin
            set_pc_commit_o        = 1'b1;
            flush_if_o             = 1'b1;
            flush_unissued_instr_o = 1'b1;
            flush_id_o             = 1'b1;
            flush_ex_o             = 1'b1;
            flush_tlb_o            = 1'b1;
        end
        
        if (flush_csr_i || flush_commit_i) begin
            set_pc_commit_o        = 1'b1;
            flush_if_o             = 1'b1;
            flush_unissued_instr_o = 1'b1;
            flush_id_o             = 1'b1;
            flush_ex_o             = 1'b1;
        end
        
        
        
        
        if (ex_valid_i || eret_i || set_debug_pc_i) begin
            
            
            set_pc_commit_o        = 1'b0;
            flush_if_o             = 1'b1;
            flush_unissued_instr_o = 1'b1;
            flush_id_o             = 1'b1;
            flush_ex_o             = 1'b1;
            
            
            
            
            flush_bp_o             = 1'b1;
        end
    end
    
    
    
    always_comb begin
        
        halt_o = halt_csr_i || fence_active_q;
    end
    
    
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (~rst_ni) begin
            fence_active_q <= 1'b0;
            flush_dcache_o <= 1'b0;
        end else begin
            fence_active_q <= fence_active_d;
            
            flush_dcache_o <= flush_dcache;
        end
    end
endmodule
module csr_buffer import ariane_pkg::*; (
    input  logic                     clk_i,          
    input  logic                     rst_ni,         
    input  logic                     flush_i,
    input  fu_data_t                 fu_data_i,
    output logic                     csr_ready_o,    
    input  logic                     csr_valid_i,    
    output riscv::xlen_t             csr_result_o,
    input  logic                     csr_commit_i,   
    
    output logic  [11:0]             csr_addr_o      
);
    
    
    struct packed {
        logic [11:0] csr_address;
        logic        valid;
    } csr_reg_n, csr_reg_q;
    
    assign csr_result_o   = fu_data_i.operand_a;
    assign csr_addr_o     = csr_reg_q.csr_address;
    
    always_comb begin : write
        csr_reg_n  = csr_reg_q;
        
        csr_ready_o = 1'b1;
        
        if ((csr_reg_q.valid || csr_valid_i) && ~csr_commit_i)
            csr_ready_o = 1'b0;
        
        
        if (csr_valid_i) begin
            csr_reg_n.csr_address = fu_data_i.operand_b[11:0];
            csr_reg_n.valid       = 1'b1;
        end
        
        if (csr_commit_i && ~csr_valid_i) begin
            csr_reg_n.valid       = 1'b0;
        end
        
        if (flush_i)
            csr_reg_n.valid       = 1'b0;
    end
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if(~rst_ni) begin
            csr_reg_q <= '{default: 0};
        end else begin
            csr_reg_q <= csr_reg_n;
        end
    end
endmodule
module csr_regfile import ariane_pkg::*; #(
    parameter logic [63:0] DmBaseAddress   = 64'h0, 
    parameter int          AsidWidth       = 1,
    parameter int unsigned NrCommitPorts   = 2,
    parameter int unsigned NrPMPEntries    = 8
) (
    input  logic                  clk_i,                      
    input  logic                  rst_ni,                     
    input  logic                  time_irq_i,                 
    
    output logic                  flush_o,
    output logic                  halt_csr_o,                 
    
    input  scoreboard_entry_t [NrCommitPorts-1:0] commit_instr_i, 
    input  logic [NrCommitPorts-1:0]              commit_ack_i,   
    
    input  logic[riscv::VLEN-1:0] boot_addr_i,                
    input  logic[riscv::XLEN-1:0] hart_id_i,                  
    
    input exception_t             ex_i,                       
    input  fu_op                  csr_op_i,                   
    input  logic  [11:0]          csr_addr_i,                 
    input  logic[riscv::XLEN-1:0] csr_wdata_i,                
    output logic[riscv::XLEN-1:0] csr_rdata_o,                
    input  logic                  dirty_fp_state_i,           
    input  logic                  csr_write_fflags_i,         
    input  logic  [riscv::VLEN-1:0]  pc_i,                    
    output exception_t            csr_exception_o,            
                                                              
                                                              
    
    output logic  [riscv::VLEN-1:0] epc_o,                    
    output logic                  eret_o,                     
    output logic  [riscv::VLEN-1:0] trap_vector_base_o,       
    output riscv::priv_lvl_t      priv_lvl_o,                 
    
    output riscv::xs_t            fs_o,                       
    output logic [4:0]            fflags_o,                   
    output logic [2:0]            frm_o,                      
    output logic [6:0]            fprec_o,                    
    
    output irq_ctrl_t             irq_ctrl_o,                 
    
    output logic                  en_translation_o,           
    output logic                  en_ld_st_translation_o,     
    output riscv::priv_lvl_t      ld_st_priv_lvl_o,           
    output logic                  sum_o,
    output logic                  mxr_o,
    output logic[riscv::PPNW-1:0] satp_ppn_o,
    output logic [AsidWidth-1:0] asid_o,
    
    input  logic [1:0]            irq_i,                      
    input  logic                  ipi_i,                      
    input  logic                  debug_req_i,                
    output logic                  set_debug_pc_o,
    
    output logic                  tvm_o,                      
    output logic                  tw_o,                       
    output logic                  tsr_o,                      
    output logic                  debug_mode_o,               
    output logic                  single_step_o,              
    
    output logic                  icache_en_o,                
    output logic                  dcache_en_o,                
    
    output logic  [4:0]           perf_addr_o,                
    output logic[riscv::XLEN-1:0] perf_data_o,                
    input  logic[riscv::XLEN-1:0] perf_data_i,                
    output logic                  perf_we_o,
    
    output riscv::pmpcfg_t [15:0] pmpcfg_o,   
    output logic [15:0][riscv::PLEN-3:0] pmpaddr_o            
);
    
    logic        read_access_exception, update_access_exception, privilege_violation;
    logic        csr_we, csr_read;
    riscv::xlen_t csr_wdata, csr_rdata;
    riscv::priv_lvl_t   trap_to_priv_lvl;
    
    logic        en_ld_st_translation_d, en_ld_st_translation_q;
    logic  mprv;
    logic  mret;  
    logic  sret;  
    logic  dret;  
    
    logic  dirty_fp_state_csr;
    riscv::status_rv_t    mstatus_q,  mstatus_d;
    riscv::xlen_t         mstatus_extended;
    riscv::satp_t         satp_q, satp_d;
    riscv::dcsr_t         dcsr_q,     dcsr_d;
    riscv::csr_t  csr_addr;
    
    riscv::priv_lvl_t   priv_lvl_d, priv_lvl_q;
    
    logic        debug_mode_q, debug_mode_d;
    logic        mtvec_rst_load_q;
    riscv::xlen_t dpc_q,       dpc_d;
    riscv::xlen_t dscratch0_q, dscratch0_d;
    riscv::xlen_t dscratch1_q, dscratch1_d;
    riscv::xlen_t mtvec_q,     mtvec_d;
    riscv::xlen_t medeleg_q,   medeleg_d;
    riscv::xlen_t mideleg_q,   mideleg_d;
    riscv::xlen_t mip_q,       mip_d;
    riscv::xlen_t mie_q,       mie_d;
    riscv::xlen_t mcounteren_q,mcounteren_d;
    riscv::xlen_t mscratch_q,  mscratch_d;
    riscv::xlen_t mepc_q,      mepc_d;
    riscv::xlen_t mcause_q,    mcause_d;
    riscv::xlen_t mtval_q,     mtval_d;
    riscv::xlen_t stvec_q,     stvec_d;
    riscv::xlen_t scounteren_q,scounteren_d;
    riscv::xlen_t sscratch_q,  sscratch_d;
    riscv::xlen_t sepc_q,      sepc_d;
    riscv::xlen_t scause_q,    scause_d;
    riscv::xlen_t stval_q,     stval_d;
    riscv::xlen_t dcache_q,    dcache_d;
    riscv::xlen_t icache_q,    icache_d;
    logic        wfi_d,       wfi_q;
    riscv::xlen_t cycle_q,     cycle_d;
    riscv::xlen_t instret_q,   instret_d;
    riscv::pmpcfg_t [15:0]    pmpcfg_q,  pmpcfg_d;
    logic [15:0][riscv::PLEN-3:0]        pmpaddr_q,  pmpaddr_d;
    assign pmpcfg_o = pmpcfg_q[15:0];
    assign pmpaddr_o = pmpaddr_q;
    riscv::fcsr_t fcsr_q, fcsr_d;
    
    
    
    assign csr_addr = riscv::csr_t'(csr_addr_i);
    assign fs_o = mstatus_q.fs;
    
    
    
    assign mstatus_extended = riscv::IS_XLEN64 ? mstatus_q[riscv::XLEN-1:0] :
                              {mstatus_q.sd, mstatus_q.wpri3[7:0], mstatus_q[22:0]};
    always_comb begin : csr_read_process
        
        read_access_exception = 1'b0;
        csr_rdata = '0;
        perf_addr_o = csr_addr.address[4:0];
        if (csr_read) begin
            unique case (csr_addr.address)
                riscv::CSR_FFLAGS: begin
                    if (mstatus_q.fs == riscv::Off) begin
                        read_access_exception = 1'b1;
                    end else begin
                        csr_rdata = {{riscv::XLEN-5{1'b0}}, fcsr_q.fflags};
                    end
                end
                riscv::CSR_FRM: begin
                    if (mstatus_q.fs == riscv::Off) begin
                        read_access_exception = 1'b1;
                    end else begin
                        csr_rdata = {{riscv::XLEN-3{1'b0}}, fcsr_q.frm};
                    end
                end
                riscv::CSR_FCSR: begin
                    if (mstatus_q.fs == riscv::Off) begin
                        read_access_exception = 1'b1;
                    end else begin
                        csr_rdata = {{riscv::XLEN-8{1'b0}}, fcsr_q.frm, fcsr_q.fflags};
                    end
                end
                
                riscv::CSR_FTRAN: begin
                    if (mstatus_q.fs == riscv::Off) begin
                        read_access_exception = 1'b1;
                    end else begin
                        csr_rdata = {{riscv::XLEN-7{1'b0}}, fcsr_q.fprec};
                    end
                end
                
                riscv::CSR_DCSR:               csr_rdata = {{riscv::XLEN-32{1'b0}}, dcsr_q};
                riscv::CSR_DPC:                csr_rdata = dpc_q;
                riscv::CSR_DSCRATCH0:          csr_rdata = dscratch0_q;
                riscv::CSR_DSCRATCH1:          csr_rdata = dscratch1_q;
                
                riscv::CSR_TSELECT:; 
                riscv::CSR_TDATA1:;  
                riscv::CSR_TDATA2:;  
                riscv::CSR_TDATA3:;  
                
                riscv::CSR_SSTATUS: begin
                    csr_rdata = mstatus_extended & ariane_pkg::SMODE_STATUS_READ_MASK[riscv::XLEN-1:0];
                end
                riscv::CSR_SIE:                csr_rdata = mie_q & mideleg_q;
                riscv::CSR_SIP:                csr_rdata = mip_q & mideleg_q;
                riscv::CSR_STVEC:              csr_rdata = stvec_q;
                riscv::CSR_SCOUNTEREN:         csr_rdata = scounteren_q;
                riscv::CSR_SSCRATCH:           csr_rdata = sscratch_q;
                riscv::CSR_SEPC:               csr_rdata = sepc_q;
                riscv::CSR_SCAUSE:             csr_rdata = scause_q;
                riscv::CSR_STVAL:              csr_rdata = stval_q;
                riscv::CSR_SATP: begin
                    
                    if (priv_lvl_o == riscv::PRIV_LVL_S && mstatus_q.tvm) begin
                        read_access_exception = 1'b1;
                    end else begin
                        csr_rdata = satp_q;
                    end
                end
                
                riscv::CSR_MSTATUS:            csr_rdata = mstatus_extended;
                riscv::CSR_MISA:               csr_rdata = ISA_CODE;
                riscv::CSR_MEDELEG:            csr_rdata = medeleg_q;
                riscv::CSR_MIDELEG:            csr_rdata = mideleg_q;
                riscv::CSR_MIE:                csr_rdata = mie_q;
                riscv::CSR_MTVEC:              csr_rdata = mtvec_q;
                riscv::CSR_MCOUNTEREN:         csr_rdata = mcounteren_q;
                riscv::CSR_MSCRATCH:           csr_rdata = mscratch_q;
                riscv::CSR_MEPC:               csr_rdata = mepc_q;
                riscv::CSR_MCAUSE:             csr_rdata = mcause_q;
                riscv::CSR_MTVAL:              csr_rdata = mtval_q;
                riscv::CSR_MIP:                csr_rdata = mip_q;
                riscv::CSR_MVENDORID:          csr_rdata = '0; 
                riscv::CSR_MARCHID:            csr_rdata = ARIANE_MARCHID;
                riscv::CSR_MIMPID:             csr_rdata = '0; 
                riscv::CSR_MHARTID:            csr_rdata = hart_id_i;
                riscv::CSR_MCYCLE:             csr_rdata = cycle_q;
                riscv::CSR_MINSTRET:           csr_rdata = instret_q;
                
                riscv::CSR_CYCLE:              csr_rdata = cycle_q;
                riscv::CSR_INSTRET:            csr_rdata = instret_q;
                riscv::CSR_ML1_ICACHE_MISS,
                riscv::CSR_ML1_DCACHE_MISS,
                riscv::CSR_MITLB_MISS,
                riscv::CSR_MDTLB_MISS,
                riscv::CSR_MLOAD,
                riscv::CSR_MSTORE,
                riscv::CSR_MEXCEPTION,
                riscv::CSR_MEXCEPTION_RET,
                riscv::CSR_MBRANCH_JUMP,
                riscv::CSR_MCALL,
                riscv::CSR_MRET,
                riscv::CSR_MMIS_PREDICT,
                riscv::CSR_MSB_FULL,
                riscv::CSR_MIF_EMPTY,
                riscv::CSR_MHPM_COUNTER_17,
                riscv::CSR_MHPM_COUNTER_18,
                riscv::CSR_MHPM_COUNTER_19,
                riscv::CSR_MHPM_COUNTER_20,
                riscv::CSR_MHPM_COUNTER_21,
                riscv::CSR_MHPM_COUNTER_22,
                riscv::CSR_MHPM_COUNTER_23,
                riscv::CSR_MHPM_COUNTER_24,
                riscv::CSR_MHPM_COUNTER_25,
                riscv::CSR_MHPM_COUNTER_26,
                riscv::CSR_MHPM_COUNTER_27,
                riscv::CSR_MHPM_COUNTER_28,
                riscv::CSR_MHPM_COUNTER_29,
                riscv::CSR_MHPM_COUNTER_30,
                riscv::CSR_MHPM_COUNTER_31:           csr_rdata   = perf_data_i;
                
                riscv::CSR_DCACHE:           csr_rdata = dcache_q;
                riscv::CSR_ICACHE:           csr_rdata = icache_q;
                
                riscv::CSR_PMPCFG0:          csr_rdata = pmpcfg_q[7:0];
                riscv::CSR_PMPCFG2:          csr_rdata = pmpcfg_q[15:8];
                
                
                
                
                
                riscv::CSR_PMPADDR0:         csr_rdata = {10'b0, pmpaddr_q[ 0][riscv::PLEN-3:1], (pmpcfg_q[ 0].addr_mode[1] == 1'b1 ? pmpaddr_q[ 0][0] : 1'b0)};
                riscv::CSR_PMPADDR1:         csr_rdata = {10'b0, pmpaddr_q[ 1][riscv::PLEN-3:1], (pmpcfg_q[ 1].addr_mode[1] == 1'b1 ? pmpaddr_q[ 1][0] : 1'b0)};
                riscv::CSR_PMPADDR2:         csr_rdata = {10'b0, pmpaddr_q[ 2][riscv::PLEN-3:1], (pmpcfg_q[ 2].addr_mode[1] == 1'b1 ? pmpaddr_q[ 2][0] : 1'b0)};
                riscv::CSR_PMPADDR3:         csr_rdata = {10'b0, pmpaddr_q[ 3][riscv::PLEN-3:1], (pmpcfg_q[ 3].addr_mode[1] == 1'b1 ? pmpaddr_q[ 3][0] : 1'b0)};
                riscv::CSR_PMPADDR4:         csr_rdata = {10'b0, pmpaddr_q[ 4][riscv::PLEN-3:1], (pmpcfg_q[ 4].addr_mode[1] == 1'b1 ? pmpaddr_q[ 4][0] : 1'b0)};
                riscv::CSR_PMPADDR5:         csr_rdata = {10'b0, pmpaddr_q[ 5][riscv::PLEN-3:1], (pmpcfg_q[ 5].addr_mode[1] == 1'b1 ? pmpaddr_q[ 5][0] : 1'b0)};
                riscv::CSR_PMPADDR6:         csr_rdata = {10'b0, pmpaddr_q[ 6][riscv::PLEN-3:1], (pmpcfg_q[ 6].addr_mode[1] == 1'b1 ? pmpaddr_q[ 6][0] : 1'b0)};
                riscv::CSR_PMPADDR7:         csr_rdata = {10'b0, pmpaddr_q[ 7][riscv::PLEN-3:1], (pmpcfg_q[ 7].addr_mode[1] == 1'b1 ? pmpaddr_q[ 7][0] : 1'b0)};
                riscv::CSR_PMPADDR8:         csr_rdata = {10'b0, pmpaddr_q[ 8][riscv::PLEN-3:1], (pmpcfg_q[ 8].addr_mode[1] == 1'b1 ? pmpaddr_q[ 8][0] : 1'b0)};
                riscv::CSR_PMPADDR9:         csr_rdata = {10'b0, pmpaddr_q[ 9][riscv::PLEN-3:1], (pmpcfg_q[ 9].addr_mode[1] == 1'b1 ? pmpaddr_q[ 9][0] : 1'b0)};
                riscv::CSR_PMPADDR10:        csr_rdata = {10'b0, pmpaddr_q[10][riscv::PLEN-3:1], (pmpcfg_q[10].addr_mode[1] == 1'b1 ? pmpaddr_q[10][0] : 1'b0)};
                riscv::CSR_PMPADDR11:        csr_rdata = {10'b0, pmpaddr_q[11][riscv::PLEN-3:1], (pmpcfg_q[11].addr_mode[1] == 1'b1 ? pmpaddr_q[11][0] : 1'b0)};
                riscv::CSR_PMPADDR12:        csr_rdata = {10'b0, pmpaddr_q[12][riscv::PLEN-3:1], (pmpcfg_q[12].addr_mode[1] == 1'b1 ? pmpaddr_q[12][0] : 1'b0)};
                riscv::CSR_PMPADDR13:        csr_rdata = {10'b0, pmpaddr_q[13][riscv::PLEN-3:1], (pmpcfg_q[13].addr_mode[1] == 1'b1 ? pmpaddr_q[13][0] : 1'b0)};
                riscv::CSR_PMPADDR14:        csr_rdata = {10'b0, pmpaddr_q[14][riscv::PLEN-3:1], (pmpcfg_q[14].addr_mode[1] == 1'b1 ? pmpaddr_q[14][0] : 1'b0)};
                riscv::CSR_PMPADDR15:        csr_rdata = {10'b0, pmpaddr_q[15][riscv::PLEN-3:1], (pmpcfg_q[15].addr_mode[1] == 1'b1 ? pmpaddr_q[15][0] : 1'b0)};
                default: read_access_exception = 1'b1;
            endcase
        end
    end
    
    
    
    riscv::xlen_t mask;
    always_comb begin : csr_update
        automatic riscv::satp_t satp;
        automatic riscv::xlen_t instret;
        satp = satp_q;
        instret = instret_q;
        
        
        
        cycle_d = cycle_q;
        instret_d = instret_q;
        if (!debug_mode_q) begin
            
            for (int i = 0; i < NrCommitPorts; i++) begin
                if (commit_ack_i[i] && !ex_i.valid) instret++;
            end
            instret_d = instret;
            
            if (ENABLE_CYCLE_COUNT) cycle_d = cycle_q + 1'b1;
            else cycle_d = instret;
        end
        eret_o                  = 1'b0;
        flush_o                 = 1'b0;
        update_access_exception = 1'b0;
        set_debug_pc_o          = 1'b0;
        perf_we_o               = 1'b0;
        perf_data_o             = 'b0;
        fcsr_d                  = fcsr_q;
        priv_lvl_d              = priv_lvl_q;
        debug_mode_d            = debug_mode_q;
        dcsr_d                  = dcsr_q;
        dpc_d                   = dpc_q;
        dscratch0_d             = dscratch0_q;
        dscratch1_d             = dscratch1_q;
        mstatus_d               = mstatus_q;
        
        
        
        
        
        
        if (mtvec_rst_load_q) begin
            mtvec_d             = {{riscv::XLEN-riscv::VLEN{1'b0}}, boot_addr_i} + 'h40;
        end else begin
            mtvec_d             = mtvec_q;
        end
        medeleg_d               = medeleg_q;
        mideleg_d               = mideleg_q;
        mip_d                   = mip_q;
        mie_d                   = mie_q;
        mepc_d                  = mepc_q;
        mcause_d                = mcause_q;
        mcounteren_d            = mcounteren_q;
        mscratch_d              = mscratch_q;
        mtval_d                 = mtval_q;
        dcache_d                = dcache_q;
        icache_d                = icache_q;
        sepc_d                  = sepc_q;
        scause_d                = scause_q;
        stvec_d                 = stvec_q;
        scounteren_d            = scounteren_q;
        sscratch_d              = sscratch_q;
        stval_d                 = stval_q;
        satp_d                  = satp_q;
        en_ld_st_translation_d  = en_ld_st_translation_q;
        dirty_fp_state_csr      = 1'b0;
        pmpcfg_d                = pmpcfg_q;
        pmpaddr_d               = pmpaddr_q;
        
        if (csr_we) begin
            unique case (csr_addr.address)
                
                riscv::CSR_FFLAGS: begin
                    if (mstatus_q.fs == riscv::Off) begin
                        update_access_exception = 1'b1;
                    end else begin
                        dirty_fp_state_csr = 1'b1;
                        fcsr_d.fflags = csr_wdata[4:0];
                        
                        flush_o = 1'b1;
                    end
                end
                riscv::CSR_FRM: begin
                    if (mstatus_q.fs == riscv::Off) begin
                        update_access_exception = 1'b1;
                    end else begin
                        dirty_fp_state_csr = 1'b1;
                        fcsr_d.frm    = csr_wdata[2:0];
                        
                        flush_o = 1'b1;
                    end
                end
                riscv::CSR_FCSR: begin
                    if (mstatus_q.fs == riscv::Off) begin
                        update_access_exception = 1'b1;
                    end else begin
                        dirty_fp_state_csr = 1'b1;
                        fcsr_d[7:0] = csr_wdata[7:0]; 
                        
                        flush_o = 1'b1;
                    end
                end
                riscv::CSR_FTRAN: begin
                    if (mstatus_q.fs == riscv::Off) begin
                        update_access_exception = 1'b1;
                    end else begin
                        dirty_fp_state_csr = 1'b1;
                        fcsr_d.fprec = csr_wdata[6:0]; 
                        
                        flush_o = 1'b1;
                    end
                end
                
                riscv::CSR_DCSR: begin
                    dcsr_d = csr_wdata[31:0];
                    
                    dcsr_d.xdebugver = 4'h4;
                    
                    dcsr_d.nmip      = 1'b0;
                    dcsr_d.stopcount = 1'b0;
                    dcsr_d.stoptime  = 1'b0;
                end
                riscv::CSR_DPC:                dpc_d = csr_wdata;
                riscv::CSR_DSCRATCH0:          dscratch0_d = csr_wdata;
                riscv::CSR_DSCRATCH1:          dscratch1_d = csr_wdata;
                
                riscv::CSR_TSELECT:; 
                riscv::CSR_TDATA1:;  
                riscv::CSR_TDATA2:;  
                riscv::CSR_TDATA3:;  
                
                riscv::CSR_SSTATUS: begin
                    mask = ariane_pkg::SMODE_STATUS_WRITE_MASK[riscv::XLEN-1:0];
                    mstatus_d = (mstatus_q & ~{{64-riscv::XLEN{1'b0}}, mask}) | {{64-riscv::XLEN{1'b0}}, (csr_wdata & mask)};
                    
                    if (!FP_PRESENT) begin
                        mstatus_d.fs = riscv::Off;
                    end
                    
                    flush_o = 1'b1;
                end
                
                
                riscv::CSR_SIE: begin
                    
                    mie_d = (mie_q & ~mideleg_q) | (csr_wdata & mideleg_q);
                end
                riscv::CSR_SIP: begin
                    
                    mask = riscv::MIP_SSIP & mideleg_q;
                    mip_d = (mip_q & ~mask) | (csr_wdata & mask);
                end
                riscv::CSR_STVEC:              stvec_d     = {csr_wdata[riscv::XLEN-1:2], 1'b0, csr_wdata[0]};
                riscv::CSR_SCOUNTEREN:         scounteren_d = {{riscv::XLEN-32{1'b0}}, csr_wdata[31:0]};
                riscv::CSR_SSCRATCH:           sscratch_d  = csr_wdata;
                riscv::CSR_SEPC:               sepc_d      = {csr_wdata[riscv::XLEN-1:1], 1'b0};
                riscv::CSR_SCAUSE:             scause_d    = csr_wdata;
                riscv::CSR_STVAL:              stval_d     = csr_wdata;
                
                riscv::CSR_SATP: begin
                    
                    if (priv_lvl_o == riscv::PRIV_LVL_S && mstatus_q.tvm)
                        update_access_exception = 1'b1;
                    else begin
                        satp      = riscv::satp_t'(csr_wdata);
                        
                        satp.asid = satp.asid & {{(riscv::ASIDW-AsidWidth){1'b0}}, {AsidWidth{1'b1}}};
                        
                        if (riscv::vm_mode_t'(satp.mode) == riscv::ModeOff ||
                            riscv::vm_mode_t'(satp.mode) == riscv::MODE_SV) satp_d = satp;
                    end
                    
                    
                    flush_o = 1'b1;
                end
                riscv::CSR_MSTATUS: begin
                    mstatus_d      = {{64-riscv::XLEN{1'b0}}, csr_wdata};
                    mstatus_d.xs   = riscv::Off;
                    if (!FP_PRESENT) begin
                        mstatus_d.fs = riscv::Off;
                    end
                    mstatus_d.upie = 1'b0;
                    mstatus_d.uie  = 1'b0;
                    
                    flush_o        = 1'b1;
                end
                
                riscv::CSR_MISA:;
                
                
                riscv::CSR_MEDELEG: begin
                    mask = (1 << riscv::INSTR_ADDR_MISALIGNED) |
                           (1 << riscv::BREAKPOINT) |
                           (1 << riscv::ENV_CALL_UMODE) |
                           (1 << riscv::INSTR_PAGE_FAULT) |
                           (1 << riscv::LOAD_PAGE_FAULT) |
                           (1 << riscv::STORE_PAGE_FAULT);
                    medeleg_d = (medeleg_q & ~mask) | (csr_wdata & mask);
                end
                
                
                riscv::CSR_MIDELEG: begin
                    mask = riscv::MIP_SSIP | riscv::MIP_STIP | riscv::MIP_SEIP;
                    mideleg_d = (mideleg_q & ~mask) | (csr_wdata & mask);
                end
                
                riscv::CSR_MIE: begin
                    mask = riscv::MIP_SSIP | riscv::MIP_STIP | riscv::MIP_SEIP | riscv::MIP_MSIP | riscv::MIP_MTIP | riscv::MIP_MEIP;
                    mie_d = (mie_q & ~mask) | (csr_wdata & mask); 
                end
                riscv::CSR_MTVEC: begin
                    mtvec_d = {csr_wdata[riscv::XLEN-1:2], 1'b0, csr_wdata[0]};
                    
                    
                    if (csr_wdata[0]) mtvec_d = {csr_wdata[riscv::XLEN-1:8], 7'b0, csr_wdata[0]};
                end
                riscv::CSR_MCOUNTEREN:         mcounteren_d = {{riscv::XLEN-32{1'b0}}, csr_wdata[31:0]};
                riscv::CSR_MSCRATCH:           mscratch_d  = csr_wdata;
                riscv::CSR_MEPC:               mepc_d      = {csr_wdata[riscv::XLEN-1:1], 1'b0};
                riscv::CSR_MCAUSE:             mcause_d    = csr_wdata;
                riscv::CSR_MTVAL:              mtval_d     = csr_wdata;
                riscv::CSR_MIP: begin
                    mask = riscv::MIP_SSIP | riscv::MIP_STIP | riscv::MIP_SEIP;
                    mip_d = (mip_q & ~mask) | (csr_wdata & mask);
                end
                
                riscv::CSR_MCYCLE:             cycle_d     = csr_wdata;
                riscv::CSR_MINSTRET:           instret     = csr_wdata;
                riscv::CSR_ML1_ICACHE_MISS,
                riscv::CSR_ML1_DCACHE_MISS,
                riscv::CSR_MITLB_MISS,
                riscv::CSR_MDTLB_MISS,
                riscv::CSR_MLOAD,
                riscv::CSR_MSTORE,
                riscv::CSR_MEXCEPTION,
                riscv::CSR_MEXCEPTION_RET,
                riscv::CSR_MBRANCH_JUMP,
                riscv::CSR_MCALL,
                riscv::CSR_MRET,
                riscv::CSR_MMIS_PREDICT,
                riscv::CSR_MSB_FULL,
                riscv::CSR_MIF_EMPTY,
                riscv::CSR_MHPM_COUNTER_17,
                riscv::CSR_MHPM_COUNTER_18,
                riscv::CSR_MHPM_COUNTER_19,
                riscv::CSR_MHPM_COUNTER_20,
                riscv::CSR_MHPM_COUNTER_21,
                riscv::CSR_MHPM_COUNTER_22,
                riscv::CSR_MHPM_COUNTER_23,
                riscv::CSR_MHPM_COUNTER_24,
                riscv::CSR_MHPM_COUNTER_25,
                riscv::CSR_MHPM_COUNTER_26,
                riscv::CSR_MHPM_COUNTER_27,
                riscv::CSR_MHPM_COUNTER_28,
                riscv::CSR_MHPM_COUNTER_29,
                riscv::CSR_MHPM_COUNTER_30,
                riscv::CSR_MHPM_COUNTER_31: begin
                                        perf_data_o = csr_wdata;
                                        perf_we_o   = 1'b1;
                end
                riscv::CSR_DCACHE:             dcache_d    = {{riscv::XLEN-1{1'b0}}, csr_wdata[0]}; 
                riscv::CSR_ICACHE:             icache_d    = {{riscv::XLEN-1{1'b0}}, csr_wdata[0]}; 
                
                
                
                
                riscv::CSR_PMPCFG0:    for (int i = 0; i < (riscv::XLEN/8); i++) if (!pmpcfg_q[i].locked) pmpcfg_d[i]  = csr_wdata[i*8+:8];
                riscv::CSR_PMPCFG1: begin
                    if (riscv::XLEN == 32) begin
                        for (int i = 0; i < 4; i++) if (!pmpcfg_q[i+4].locked) pmpcfg_d[i+4]  = csr_wdata[i*8+:8];
                    end
                end
                riscv::CSR_PMPCFG2:    for (int i = 0; i < (riscv::XLEN/8); i++) if (!pmpcfg_q[i+8].locked) pmpcfg_d[i+8]  = csr_wdata[i*8+:8];
                riscv::CSR_PMPCFG3: begin
                    if (riscv::XLEN == 32) begin
                        for (int i = 0; i < 4; i++) if (!pmpcfg_q[i+12].locked) pmpcfg_d[i+12]  = csr_wdata[i*8+:8];
                    end
                end
                riscv::CSR_PMPADDR0:   if (!pmpcfg_q[ 0].locked && !(pmpcfg_q[ 1].locked && pmpcfg_q[ 1].addr_mode == riscv::TOR))  pmpaddr_d[0]   = csr_wdata[riscv::PLEN-3:0];
                riscv::CSR_PMPADDR1:   if (!pmpcfg_q[ 1].locked && !(pmpcfg_q[ 2].locked && pmpcfg_q[ 2].addr_mode == riscv::TOR))  pmpaddr_d[1]   = csr_wdata[riscv::PLEN-3:0];
                riscv::CSR_PMPADDR2:   if (!pmpcfg_q[ 2].locked && !(pmpcfg_q[ 3].locked && pmpcfg_q[ 3].addr_mode == riscv::TOR))  pmpaddr_d[2]   = csr_wdata[riscv::PLEN-3:0];
                riscv::CSR_PMPADDR3:   if (!pmpcfg_q[ 3].locked && !(pmpcfg_q[ 4].locked && pmpcfg_q[ 4].addr_mode == riscv::TOR))  pmpaddr_d[3]   = csr_wdata[riscv::PLEN-3:0];
                riscv::CSR_PMPADDR4:   if (!pmpcfg_q[ 4].locked && !(pmpcfg_q[ 5].locked && pmpcfg_q[ 5].addr_mode == riscv::TOR))  pmpaddr_d[4]   = csr_wdata[riscv::PLEN-3:0];
                riscv::CSR_PMPADDR5:   if (!pmpcfg_q[ 5].locked && !(pmpcfg_q[ 6].locked && pmpcfg_q[ 6].addr_mode == riscv::TOR))  pmpaddr_d[5]   = csr_wdata[riscv::PLEN-3:0];
                riscv::CSR_PMPADDR6:   if (!pmpcfg_q[ 6].locked && !(pmpcfg_q[ 7].locked && pmpcfg_q[ 7].addr_mode == riscv::TOR))  pmpaddr_d[6]   = csr_wdata[riscv::PLEN-3:0];
                riscv::CSR_PMPADDR7:   if (!pmpcfg_q[ 7].locked && !(pmpcfg_q[ 8].locked && pmpcfg_q[ 8].addr_mode == riscv::TOR))  pmpaddr_d[7]   = csr_wdata[riscv::PLEN-3:0];
                riscv::CSR_PMPADDR8:   if (!pmpcfg_q[ 8].locked && !(pmpcfg_q[ 9].locked && pmpcfg_q[ 9].addr_mode == riscv::TOR))  pmpaddr_d[8]   = csr_wdata[riscv::PLEN-3:0];
                riscv::CSR_PMPADDR9:   if (!pmpcfg_q[ 9].locked && !(pmpcfg_q[10].locked && pmpcfg_q[10].addr_mode == riscv::TOR))  pmpaddr_d[9]   = csr_wdata[riscv::PLEN-3:0];
                riscv::CSR_PMPADDR10:  if (!pmpcfg_q[10].locked && !(pmpcfg_q[11].locked && pmpcfg_q[11].addr_mode == riscv::TOR))  pmpaddr_d[10]  = csr_wdata[riscv::PLEN-3:0];
                riscv::CSR_PMPADDR11:  if (!pmpcfg_q[11].locked && !(pmpcfg_q[12].locked && pmpcfg_q[12].addr_mode == riscv::TOR))  pmpaddr_d[11]  = csr_wdata[riscv::PLEN-3:0];
                riscv::CSR_PMPADDR12:  if (!pmpcfg_q[12].locked && !(pmpcfg_q[13].locked && pmpcfg_q[13].addr_mode == riscv::TOR))  pmpaddr_d[12]  = csr_wdata[riscv::PLEN-3:0];
                riscv::CSR_PMPADDR13:  if (!pmpcfg_q[13].locked && !(pmpcfg_q[14].locked && pmpcfg_q[14].addr_mode == riscv::TOR))  pmpaddr_d[13]  = csr_wdata[riscv::PLEN-3:0];
                riscv::CSR_PMPADDR14:  if (!pmpcfg_q[14].locked && !(pmpcfg_q[15].locked && pmpcfg_q[15].addr_mode == riscv::TOR))  pmpaddr_d[14]  = csr_wdata[riscv::PLEN-3:0];
                riscv::CSR_PMPADDR15:  if (!pmpcfg_q[15].locked)  pmpaddr_d[15]  = csr_wdata[riscv::PLEN-3:0];
                default: update_access_exception = 1'b1;
            endcase
        end
        mstatus_d.sxl  = riscv::XLEN_64;
        mstatus_d.uxl  = riscv::XLEN_64;
        
        if (FP_PRESENT && (dirty_fp_state_csr || dirty_fp_state_i)) begin
            mstatus_d.fs = riscv::Dirty;
        end
        
        mstatus_d.sd   = (mstatus_q.xs == riscv::Dirty) | (mstatus_q.fs == riscv::Dirty);
        
        if (csr_write_fflags_i) begin
            fcsr_d.fflags = csr_wdata_i[4:0] | fcsr_q.fflags;
        end
        
        
        
        
        mip_d[riscv::IRQ_M_EXT] = irq_i[0];
        
        mip_d[riscv::IRQ_M_SOFT] = ipi_i;
        
        mip_d[riscv::IRQ_M_TIMER] = time_irq_i;
        
        
        
        
        
        trap_to_priv_lvl = riscv::PRIV_LVL_M;
        
        
        if (!debug_mode_q && ex_i.cause != riscv::DEBUG_REQUEST && ex_i.valid) begin
            
            flush_o   = 1'b0;
            
            
            
            
            if ((ex_i.cause[riscv::XLEN-1] && mideleg_q[ex_i.cause[$clog2(riscv::XLEN)-1:0]]) ||
                (~ex_i.cause[riscv::XLEN-1] && medeleg_q[ex_i.cause[$clog2(riscv::XLEN)-1:0]])) begin
                
                
                trap_to_priv_lvl = (priv_lvl_o == riscv::PRIV_LVL_M) ? riscv::PRIV_LVL_M : riscv::PRIV_LVL_S;
            end
            
            if (trap_to_priv_lvl == riscv::PRIV_LVL_S) begin
                
                mstatus_d.sie  = 1'b0;
                mstatus_d.spie = mstatus_q.sie;
                
                mstatus_d.spp  = priv_lvl_q[0];
                
                scause_d       = ex_i.cause;
                
                sepc_d         = {{riscv::XLEN-riscv::VLEN{pc_i[riscv::VLEN-1]}},pc_i};
                
                stval_d        = (ariane_pkg::ZERO_TVAL
                                  && (ex_i.cause inside {
                                    riscv::ILLEGAL_INSTR,
                                    riscv::BREAKPOINT,
                                    riscv::ENV_CALL_UMODE,
                                    riscv::ENV_CALL_SMODE,
                                    riscv::ENV_CALL_MMODE
                                  } || ex_i.cause[riscv::XLEN-1])) ? '0 : ex_i.tval;
            
            end else begin
                
                mstatus_d.mie  = 1'b0;
                mstatus_d.mpie = mstatus_q.mie;
                
                mstatus_d.mpp  = priv_lvl_q;
                mcause_d       = ex_i.cause;
                
                mepc_d         = {{riscv::XLEN-riscv::VLEN{pc_i[riscv::VLEN-1]}},pc_i};
                
                mtval_d        = (ariane_pkg::ZERO_TVAL
                                  && (ex_i.cause inside {
                                    riscv::ILLEGAL_INSTR,
                                    riscv::BREAKPOINT,
                                    riscv::ENV_CALL_UMODE,
                                    riscv::ENV_CALL_SMODE,
                                    riscv::ENV_CALL_MMODE
                                  } || ex_i.cause[riscv::XLEN-1])) ? '0 : ex_i.tval;
            end
            priv_lvl_d = trap_to_priv_lvl;
        end
        
        
        
        
        
        
        
        
        
        
        if (!debug_mode_q) begin
            dcsr_d.prv = priv_lvl_o;
            
            
            if (ex_i.valid && ex_i.cause == riscv::BREAKPOINT) begin
                dcsr_d.prv = priv_lvl_o;
                
                unique case (priv_lvl_o)
                    riscv::PRIV_LVL_M: begin
                        debug_mode_d = dcsr_q.ebreakm;
                        set_debug_pc_o = dcsr_q.ebreakm;
                    end
                    riscv::PRIV_LVL_S: begin
                        debug_mode_d = dcsr_q.ebreaks;
                        set_debug_pc_o = dcsr_q.ebreaks;
                    end
                    riscv::PRIV_LVL_U: begin
                        debug_mode_d = dcsr_q.ebreaku;
                        set_debug_pc_o = dcsr_q.ebreaku;
                    end
                    default:;
                endcase
                
                dpc_d = {{riscv::XLEN-riscv::VLEN{pc_i[riscv::VLEN-1]}},pc_i};
                dcsr_d.cause = dm::CauseBreakpoint;
            end
            
            if (ex_i.valid && ex_i.cause == riscv::DEBUG_REQUEST) begin
                dcsr_d.prv = priv_lvl_o;
                
                dpc_d = {{riscv::XLEN-riscv::VLEN{pc_i[riscv::VLEN-1]}},pc_i};
                
                debug_mode_d = 1'b1;
                
                set_debug_pc_o = 1'b1;
                
                dcsr_d.cause = dm::CauseRequest;
            end
            
            if (dcsr_q.step && commit_ack_i[0]) begin
                dcsr_d.prv = priv_lvl_o;
                
                if (commit_instr_i[0].fu == CTRL_FLOW) begin
                    
                    dpc_d = {{riscv::XLEN-riscv::VLEN{commit_instr_i[0].bp.predict_address[riscv::VLEN-1]}}, commit_instr_i[0].bp.predict_address};
                
                end else if (ex_i.valid) begin
                    dpc_d = {{riscv::XLEN-riscv::VLEN{1'b0}},trap_vector_base_o};
                
                end else if (eret_o) begin
                    dpc_d = {{riscv::XLEN-riscv::VLEN{1'b0}},epc_o};
                
                end else begin
                    dpc_d = {{riscv::XLEN-riscv::VLEN{commit_instr_i[0].pc[riscv::VLEN-1]}}, commit_instr_i[0].pc + (commit_instr_i[0].is_compressed ? 'h2 : 'h4)};
                end
                debug_mode_d = 1'b1;
                set_debug_pc_o = 1'b1;
                dcsr_d.cause = dm::CauseSingleStep;
            end
        end
        
        if (debug_mode_q && ex_i.valid && ex_i.cause == riscv::BREAKPOINT) begin
            set_debug_pc_o = 1'b1;
        end
        
        
        
        
        
        if (mprv && riscv::vm_mode_t'(satp_q.mode) == riscv::MODE_SV && (mstatus_q.mpp != riscv::PRIV_LVL_M))
            en_ld_st_translation_d = 1'b1;
        else 
            en_ld_st_translation_d = en_translation_o;
        ld_st_priv_lvl_o = (mprv) ? mstatus_q.mpp : priv_lvl_o;
        en_ld_st_translation_o = en_ld_st_translation_q;
        
        
        
        
        
        if (mret) begin
            
            eret_o = 1'b1;
            
            
            mstatus_d.mie  = mstatus_q.mpie;
            
            priv_lvl_d     = mstatus_q.mpp;
            
            mstatus_d.mpp  = riscv::PRIV_LVL_U;
            
            mstatus_d.mpie = 1'b1;
        end
        if (sret) begin
            
            eret_o = 1'b1;
            
            mstatus_d.sie  = mstatus_q.spie;
            
            priv_lvl_d     = riscv::priv_lvl_t'({1'b0, mstatus_q.spp});
            
            mstatus_d.spp  = 1'b0;
            
            mstatus_d.spie = 1'b1;
        end
        
        if (dret) begin
            
            eret_o = 1'b1;
            
            priv_lvl_d     = riscv::priv_lvl_t'(dcsr_q.prv);
            
            debug_mode_d = 1'b0;
        end
    end
    
    
    
    always_comb begin : csr_op_logic
        csr_wdata = csr_wdata_i;
        csr_we    = 1'b1;
        csr_read  = 1'b1;
        mret      = 1'b0;
        sret      = 1'b0;
        dret      = 1'b0;
        unique case (csr_op_i)
            CSR_WRITE: csr_wdata = csr_wdata_i;
            CSR_SET:   csr_wdata = csr_wdata_i | csr_rdata;
            CSR_CLEAR: csr_wdata = (~csr_wdata_i) & csr_rdata;
            CSR_READ:  csr_we    = 1'b0;
            SRET: begin
                
                csr_we   = 1'b0;
                csr_read = 1'b0;
                sret     = 1'b1; 
            end
            MRET: begin
                
                csr_we   = 1'b0;
                csr_read = 1'b0;
                mret     = 1'b1; 
            end
            DRET: begin
                
                csr_we   = 1'b0;
                csr_read = 1'b0;
                dret     = 1'b1; 
            end
            default: begin
                csr_we   = 1'b0;
                csr_read = 1'b0;
            end
        endcase
        
        if (privilege_violation) begin
            csr_we = 1'b0;
            csr_read = 1'b0;
        end
    end
    assign irq_ctrl_o.mie = mie_q;
    assign irq_ctrl_o.mip = mip_q;
    assign irq_ctrl_o.sie = mstatus_q.sie;
    assign irq_ctrl_o.mideleg = mideleg_q;
    assign irq_ctrl_o.global_enable = (~debug_mode_q)
                                    
                                    & (~dcsr_q.step | dcsr_q.stepie)
                                    & ((mstatus_q.mie & (priv_lvl_o == riscv::PRIV_LVL_M))
                                    | (priv_lvl_o != riscv::PRIV_LVL_M));
    always_comb begin : privilege_check
        
        
        
        privilege_violation = 1'b0;
        
        
        if (csr_op_i inside {CSR_WRITE, CSR_SET, CSR_CLEAR, CSR_READ}) begin
            if ((riscv::priv_lvl_t'(priv_lvl_o & csr_addr.csr_decode.priv_lvl) != csr_addr.csr_decode.priv_lvl)) begin
                privilege_violation = 1'b1;
            end
            
            if (csr_addr_i[11:4] == 8'h7b && !debug_mode_q) begin
                privilege_violation = 1'b1;
            end
            
            
            if (csr_addr_i inside {[riscv::CSR_CYCLE:riscv::CSR_HPM_COUNTER_31]}) begin
                unique case (priv_lvl_o)
                    riscv::PRIV_LVL_M: privilege_violation = 1'b0;
                    riscv::PRIV_LVL_S: privilege_violation = ~mcounteren_q[csr_addr_i[4:0]];
                    riscv::PRIV_LVL_U: privilege_violation = ~mcounteren_q[csr_addr_i[4:0]] & ~scounteren_q[csr_addr_i[4:0]];
                endcase
            end
        end
    end
    
    
    
    always_comb begin : exception_ctrl
        csr_exception_o = {
            '0, '0, 1'b0
        };
        
        
        
        
        
        if (update_access_exception || read_access_exception) begin
            csr_exception_o.cause = riscv::ILLEGAL_INSTR;
            
            
            csr_exception_o.valid = 1'b1;
        end
        if (privilege_violation) begin
          csr_exception_o.cause = riscv::ILLEGAL_INSTR;
          csr_exception_o.valid = 1'b1;
        end
    end
    
    
    
    always_comb begin : wfi_ctrl
        
        wfi_d = wfi_q;
        
        
        if (|mip_q || debug_req_i || irq_i[1]) begin
            wfi_d = 1'b0;
        
        
        end else if (!debug_mode_q && csr_op_i == WFI && !ex_i.valid) begin
            wfi_d = 1'b1;
        end
    end
    
    always_comb begin : priv_output
        trap_vector_base_o = {mtvec_q[riscv::VLEN-1:2], 2'b0};
        
        if (trap_to_priv_lvl == riscv::PRIV_LVL_S) begin
            trap_vector_base_o = {stvec_q[riscv::VLEN-1:2], 2'b0};
        end
        
        if (debug_mode_q) begin
            trap_vector_base_o = DmBaseAddress[riscv::VLEN-1:0] + dm::ExceptionAddress[riscv::VLEN-1:0];
        end
        
        
        
        if ((mtvec_q[0] || stvec_q[0]) && ex_i.cause[riscv::XLEN-1]) begin
            trap_vector_base_o[7:2] = ex_i.cause[5:0];
        end
        epc_o = mepc_q[riscv::VLEN-1:0];
        
        if (sret) begin
            epc_o = sepc_q[riscv::VLEN-1:0];
        end
        
        if (dret) begin
            epc_o = dpc_q[riscv::VLEN-1:0];
        end
    end
    
    
    
    always_comb begin
        
        
        
        csr_rdata_o = csr_rdata;
        unique case (csr_addr.address)
            riscv::CSR_MIP: csr_rdata_o = csr_rdata | (irq_i[1] << riscv::IRQ_S_EXT);
            
            riscv::CSR_SIP: begin
                csr_rdata_o = csr_rdata
                            | ((irq_i[1] & mideleg_q[riscv::IRQ_S_EXT]) << riscv::IRQ_S_EXT);
            end
            default:;
        endcase
    end
    
    assign priv_lvl_o       = (debug_mode_q) ? riscv::PRIV_LVL_M : priv_lvl_q;
    
    assign fflags_o         = fcsr_q.fflags;
    assign frm_o            = fcsr_q.frm;
    assign fprec_o          = fcsr_q.fprec;
    
    assign satp_ppn_o       = satp_q.ppn;
    assign asid_o           = satp_q.asid[AsidWidth-1:0];
    assign sum_o            = mstatus_q.sum;
    
    assign en_translation_o = (riscv::vm_mode_t'(satp_q.mode) == riscv::MODE_SV &&
                               priv_lvl_o != riscv::PRIV_LVL_M)
                              ? 1'b1
                              : 1'b0;
    assign mxr_o            = mstatus_q.mxr;
    assign tvm_o            = mstatus_q.tvm;
    assign tw_o             = mstatus_q.tw;
    assign tsr_o            = mstatus_q.tsr;
    assign halt_csr_o       = wfi_q;
    assign icache_en_o      = icache_q[0];
    assign dcache_en_o      = dcache_q[0];
    
    assign mprv             = (debug_mode_q && !dcsr_q.mprven) ? 1'b0 : mstatus_q.mprv;
    assign debug_mode_o     = debug_mode_q;
    assign single_step_o    = dcsr_q.step;
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (~rst_ni) begin
            priv_lvl_q             <= riscv::PRIV_LVL_M;
            
            fcsr_q                 <= '0;
            
            debug_mode_q           <= 1'b0;
            dcsr_q                 <= '0;
            dcsr_q.prv             <= riscv::PRIV_LVL_M;
            dcsr_q.xdebugver       <= 4'h4;
            dpc_q                  <= '0;
            dscratch0_q            <= {riscv::XLEN{1'b0}};
            dscratch1_q            <= {riscv::XLEN{1'b0}};
            
            mstatus_q              <= 64'b0;
            
            mtvec_rst_load_q       <= 1'b1;
            mtvec_q                <= '0;
            medeleg_q              <= {riscv::XLEN{1'b0}};
            mideleg_q              <= {riscv::XLEN{1'b0}};
            mip_q                  <= {riscv::XLEN{1'b0}};
            mie_q                  <= {riscv::XLEN{1'b0}};
            mepc_q                 <= {riscv::XLEN{1'b0}};
            mcause_q               <= {riscv::XLEN{1'b0}};
            mcounteren_q           <= {riscv::XLEN{1'b0}};
            mscratch_q             <= {riscv::XLEN{1'b0}};
            mtval_q                <= {riscv::XLEN{1'b0}};
            dcache_q               <= {{riscv::XLEN-1{1'b0}}, 1'b1};
            icache_q               <= {{riscv::XLEN-1{1'b0}}, 1'b1};
            
            sepc_q                 <= {riscv::XLEN{1'b0}};
            scause_q               <= {riscv::XLEN{1'b0}};
            stvec_q                <= {riscv::XLEN{1'b0}};
            scounteren_q           <= {riscv::XLEN{1'b0}};
            sscratch_q             <= {riscv::XLEN{1'b0}};
            stval_q                <= {riscv::XLEN{1'b0}};
            satp_q                 <= {riscv::XLEN{1'b0}};
            
            cycle_q                <= {riscv::XLEN{1'b0}};
            instret_q              <= {riscv::XLEN{1'b0}};
            
            en_ld_st_translation_q <= 1'b0;
            
            wfi_q                  <= 1'b0;
            
            pmpcfg_q               <= '0;
            pmpaddr_q              <= '0;
        end else begin
            priv_lvl_q             <= priv_lvl_d;
            
            fcsr_q                 <= fcsr_d;
            
            debug_mode_q           <= debug_mode_d;
            dcsr_q                 <= dcsr_d;
            dpc_q                  <= dpc_d;
            dscratch0_q            <= dscratch0_d;
            dscratch1_q            <= dscratch1_d;
            
            mstatus_q              <= mstatus_d;
            mtvec_rst_load_q       <= 1'b0;
            mtvec_q                <= mtvec_d;
            medeleg_q              <= medeleg_d;
            mideleg_q              <= mideleg_d;
            mip_q                  <= mip_d;
            mie_q                  <= mie_d;
            mepc_q                 <= mepc_d;
            mcause_q               <= mcause_d;
            mcounteren_q           <= mcounteren_d;
            mscratch_q             <= mscratch_d;
            mtval_q                <= mtval_d;
            dcache_q               <= dcache_d;
            icache_q               <= icache_d;
            
            sepc_q                 <= sepc_d;
            scause_q               <= scause_d;
            stvec_q                <= stvec_d;
            scounteren_q           <= scounteren_d;
            sscratch_q             <= sscratch_d;
            stval_q                <= stval_d;
            satp_q                 <= satp_d;
            
            cycle_q                <= cycle_d;
            instret_q              <= instret_d;
            
            en_ld_st_translation_q <= en_ld_st_translation_d;
            
            wfi_q                  <= wfi_d;
            
            for(int i = 0; i < 16; i++) begin
                if(i < NrPMPEntries) begin
                    
                    if(pmpcfg_q[i].addr_mode != riscv::NA4) 
                        pmpcfg_q[i] <= pmpcfg_d[i];
                    else
                        pmpcfg_q[i] <= pmpcfg_q[i];
                    pmpaddr_q[i] <= pmpaddr_d[i];
                end else begin
                    pmpcfg_q[i] <= '0;
                    pmpaddr_q[i] <= '0;
                end
            end
        end
    end
    
    
    
    
    
    
    
endmodule
module decoder import ariane_pkg::*; (
    input  logic               debug_req_i,             
    input  logic [riscv::VLEN-1:0] pc_i,                
    input  logic               is_compressed_i,         
    input  logic [15:0]        compressed_instr_i,      
    input  logic               is_illegal_i,            
    input  logic [31:0]        instruction_i,           
    input  branchpredict_sbe_t branch_predict_i,
    input  exception_t         ex_i,                    
    input  logic [1:0]         irq_i,                   
    input  irq_ctrl_t          irq_ctrl_i,              
    
    input  riscv::priv_lvl_t   priv_lvl_i,              
    input  logic               debug_mode_i,            
    input  riscv::xs_t         fs_i,                    
    input  logic [2:0]         frm_i,                   
    input  logic               tvm_i,                   
    input  logic               tw_i,                    
    input  logic               tsr_i,                   
    output scoreboard_entry_t  instruction_o,           
    output logic               is_control_flow_instr_o  
);
    logic illegal_instr;
    
    logic ecall;
    
    logic ebreak;
    
    logic check_fprm;
    riscv::instruction_t instr;
    assign instr = riscv::instruction_t'(instruction_i);
    
    
    
    enum logic[3:0] {
        NOIMM, IIMM, SIMM, SBIMM, UIMM, JIMM, RS3
    } imm_select;
    riscv::xlen_t imm_i_type;
    riscv::xlen_t imm_s_type;
    riscv::xlen_t imm_sb_type;
    riscv::xlen_t imm_u_type;
    riscv::xlen_t imm_uj_type;
    riscv::xlen_t imm_bi_type;
    always_comb begin : decoder
        imm_select                  = NOIMM;
        is_control_flow_instr_o     = 1'b0;
        illegal_instr               = 1'b0;
        instruction_o.pc            = pc_i;
        instruction_o.trans_id      = 5'b0;
        instruction_o.fu            = NONE;
        instruction_o.op            = ariane_pkg::ADD;
        instruction_o.rs1           = '0;
        instruction_o.rs2           = '0;
        instruction_o.rd            = '0;
        instruction_o.use_pc        = 1'b0;
        instruction_o.trans_id      = '0;
        instruction_o.is_compressed = is_compressed_i;
        instruction_o.use_zimm      = 1'b0;
        instruction_o.bp            = branch_predict_i;
        ecall                       = 1'b0;
        ebreak                      = 1'b0;
        check_fprm                  = 1'b0;
        if (~ex_i.valid) begin
            case (instr.rtype.opcode)
                riscv::OpcodeSystem: begin
                    instruction_o.fu       = CSR;
                    instruction_o.rs1[4:0] = instr.itype.rs1;
                    instruction_o.rs2[4:0] = instr.rtype.rs2;   
                    instruction_o.rd[4:0]  = instr.itype.rd;
                    unique case (instr.itype.funct3)
                        3'b000: begin
                            
                            if (instr.itype.rs1 != '0 || instr.itype.rd != '0)
                                illegal_instr = 1'b1;
                            
                            case (instr.itype.imm)
                                
                                12'b0: ecall  = 1'b1;
                                
                                12'b1: ebreak = 1'b1;
                                
                                12'b1_0000_0010: begin
                                    instruction_o.op = ariane_pkg::SRET;
                                    
                                    
                                    if (priv_lvl_i == riscv::PRIV_LVL_U) begin
                                        illegal_instr = 1'b1;
                                        
                                        instruction_o.op = ariane_pkg::ADD;
                                    end
                                    
                                    if (priv_lvl_i == riscv::PRIV_LVL_S && tsr_i) begin
                                        illegal_instr = 1'b1;
                                        
                                        instruction_o.op = ariane_pkg::ADD;
                                    end
                                end
                                
                                12'b11_0000_0010: begin
                                    instruction_o.op = ariane_pkg::MRET;
                                    
                                    
                                    if (priv_lvl_i inside {riscv::PRIV_LVL_U, riscv::PRIV_LVL_S})
                                        illegal_instr = 1'b1;
                                end
                                
                                12'b111_1011_0010: begin
                                    instruction_o.op = ariane_pkg::DRET;
                                    
                                    illegal_instr = (!debug_mode_i) ? 1'b1 : 1'b0;
                                end
                                
                                12'b1_0000_0101: begin
                                    if (ENABLE_WFI) instruction_o.op = ariane_pkg::WFI;
                                    
                                    
                                    if (priv_lvl_i == riscv::PRIV_LVL_S && tw_i) begin
                                        illegal_instr = 1'b1;
                                        instruction_o.op = ariane_pkg::ADD;
                                    end
                                    
                                    if (priv_lvl_i == riscv::PRIV_LVL_U) begin
                                        illegal_instr = 1'b1;
                                        instruction_o.op = ariane_pkg::ADD;
                                    end
                                end
                                
                                default: begin
                                    if (instr.instr[31:25] == 7'b1001) begin
                                        
                                        
                                        illegal_instr    = (priv_lvl_i inside {riscv::PRIV_LVL_M, riscv::PRIV_LVL_S}) ? 1'b0 : 1'b1;
                                        instruction_o.op = ariane_pkg::SFENCE_VMA;
                                        
                                        if (priv_lvl_i == riscv::PRIV_LVL_S && tvm_i)
                                            illegal_instr = 1'b1;
                                    end
                                end
                            endcase
                        end
                        
                        3'b001: begin
                            imm_select = IIMM;
                            instruction_o.op = ariane_pkg::CSR_WRITE;
                        end
                        
                        3'b010: begin
                            imm_select = IIMM;
                            
                            if (instr.itype.rs1 == 5'b0)
                                instruction_o.op = ariane_pkg::CSR_READ;
                            else
                                instruction_o.op = ariane_pkg::CSR_SET;
                        end
                        
                        3'b011: begin
                            imm_select = IIMM;
                            
                            if (instr.itype.rs1 == 5'b0)
                                instruction_o.op = ariane_pkg::CSR_READ;
                            else
                                instruction_o.op = ariane_pkg::CSR_CLEAR;
                        end
                        
                        3'b101: begin
                            instruction_o.rs1[4:0] = instr.itype.rs1;
                            imm_select = IIMM;
                            instruction_o.use_zimm = 1'b1;
                            instruction_o.op = ariane_pkg::CSR_WRITE;
                        end
                        3'b110: begin
                            instruction_o.rs1[4:0] = instr.itype.rs1;
                            imm_select = IIMM;
                            instruction_o.use_zimm = 1'b1;
                            
                            if (instr.itype.rs1 == 5'b0)
                                instruction_o.op = ariane_pkg::CSR_READ;
                            else
                                instruction_o.op = ariane_pkg::CSR_SET;
                        end
                        3'b111: begin
                            instruction_o.rs1[4:0] = instr.itype.rs1;
                            imm_select = IIMM;
                            instruction_o.use_zimm = 1'b1;
                            
                            if (instr.itype.rs1 == 5'b0)
                                instruction_o.op = ariane_pkg::CSR_READ;
                            else
                                instruction_o.op = ariane_pkg::CSR_CLEAR;
                        end
                        default: illegal_instr = 1'b1;
                    endcase
                end
                
                riscv::OpcodeMiscMem: begin
                    instruction_o.fu  = CSR;
                    instruction_o.rs1 = '0;
                    instruction_o.rs2 = '0;
                    instruction_o.rd  = '0;
                    case (instr.stype.funct3)
                        
                        
                        3'b000: instruction_o.op  = ariane_pkg::FENCE;
                        
                        3'b001: begin
                            if (instr.instr[31:20] != '0)
                                illegal_instr = 1'b1;
                            instruction_o.op  = ariane_pkg::FENCE_I;
                        end
                        default: illegal_instr = 1'b1;
                    endcase
                    if (instr.stype.rs1 != '0 || instr.stype.imm0 != '0 || instr.instr[31:28] != '0)
                        illegal_instr = 1'b1;
                end
                
                
                
                riscv::OpcodeOp: begin
                    
                    
                    
                    if (instr.rvftype.funct2 == 2'b10) begin 
                        
                        if (FP_PRESENT && XFVEC && fs_i != riscv::Off) begin
                            automatic logic allow_replication; 
                            instruction_o.fu       = FPU_VEC; 
                            instruction_o.rs1[4:0] = instr.rvftype.rs1;
                            instruction_o.rs2[4:0] = instr.rvftype.rs2;
                            instruction_o.rd[4:0]  = instr.rvftype.rd;
                            check_fprm             = 1'b1;
                            allow_replication      = 1'b1;
                            
                            unique case (instr.rvftype.vecfltop)
                                5'b00001 : begin
                                    instruction_o.op  = ariane_pkg::FADD; 
                                    instruction_o.rs1 = '0;                
                                    instruction_o.rs2 = instr.rvftype.rs1; 
                                    imm_select        = IIMM;              
                                end
                                5'b00010 : begin
                                    instruction_o.op  = ariane_pkg::FSUB; 
                                    instruction_o.rs1 = '0;                
                                    instruction_o.rs2 = instr.rvftype.rs1; 
                                    imm_select        = IIMM;              
                                end
                                5'b00011 : instruction_o.op = ariane_pkg::FMUL; 
                                5'b00100 : instruction_o.op = ariane_pkg::FDIV; 
                                5'b00101 : begin
                                    instruction_o.op = ariane_pkg::VFMIN; 
                                    check_fprm       = 1'b0;  
                                end
                                5'b00110 : begin
                                    instruction_o.op = ariane_pkg::VFMAX; 
                                    check_fprm       = 1'b0;  
                                end
                                5'b00111 : begin
                                    instruction_o.op  = ariane_pkg::FSQRT; 
                                    allow_replication = 1'b0;  
                                    if (instr.rvftype.rs2 != 5'b00000) illegal_instr = 1'b1; 
                                end
                                5'b01000 : begin
                                    instruction_o.op = ariane_pkg::FMADD; 
                                    imm_select       = SIMM;  
                                end
                                5'b01001 : begin
                                    instruction_o.op = ariane_pkg::FMSUB; 
                                    imm_select       = SIMM;  
                                end
                                5'b01100 : begin
                                    unique case (instr.rvftype.rs2) inside 
                                        5'b00000 : begin
                                            instruction_o.rs2 = instr.rvftype.rs1; 
                                            if (instr.rvftype.repl)
                                                instruction_o.op = ariane_pkg::FMV_X2F; 
                                            else
                                                instruction_o.op = ariane_pkg::FMV_F2X; 
                                            check_fprm = 1'b0;              
                                        end
                                        5'b00001 : begin
                                            instruction_o.op  = ariane_pkg::FCLASS; 
                                            check_fprm        = 1'b0;   
                                            allow_replication = 1'b0;   
                                        end
                                        5'b00010 : instruction_o.op = ariane_pkg::FCVT_F2I; 
                                        5'b00011 : instruction_o.op = ariane_pkg::FCVT_I2F; 
                                        5'b001?? : begin
                                            instruction_o.op  = ariane_pkg::FCVT_F2F; 
                                            instruction_o.rs2 = instr.rvftype.rd; 
                                            imm_select        = IIMM;     
                                            
                                            
                                            unique case (instr.rvftype.rs2[21:20])
                                                
                                                2'b00: if (~RVFVEC)     illegal_instr = 1'b1;
                                                2'b01: if (~XF16ALTVEC) illegal_instr = 1'b1;
                                                2'b10: if (~XF16VEC)    illegal_instr = 1'b1;
                                                2'b11: if (~XF8VEC)     illegal_instr = 1'b1;
                                                default : illegal_instr = 1'b1;
                                            endcase
                                        end
                                        default : illegal_instr = 1'b1;
                                    endcase
                                end
                                5'b01101 : begin
                                    check_fprm = 1'b0;         
                                    instruction_o.op = ariane_pkg::VFSGNJ; 
                                end
                                5'b01110 : begin
                                    check_fprm = 1'b0;          
                                    instruction_o.op = ariane_pkg::VFSGNJN; 
                                end
                                5'b01111 : begin
                                    check_fprm = 1'b0;          
                                    instruction_o.op = ariane_pkg::VFSGNJX; 
                                end
                                5'b10000 : begin
                                    check_fprm = 1'b0;          
                                    instruction_o.op = ariane_pkg::VFEQ;    
                                end
                                5'b10001 : begin
                                    check_fprm = 1'b0;          
                                    instruction_o.op = ariane_pkg::VFNE;    
                                end
                                5'b10010 : begin
                                    check_fprm = 1'b0;          
                                    instruction_o.op = ariane_pkg::VFLT;    
                                end
                                5'b10011 : begin
                                    check_fprm = 1'b0;          
                                    instruction_o.op = ariane_pkg::VFGE;    
                                end
                                5'b10100 : begin
                                    check_fprm = 1'b0;          
                                    instruction_o.op = ariane_pkg::VFLE;    
                                end
                                5'b10101 : begin
                                    check_fprm = 1'b0;          
                                    instruction_o.op = ariane_pkg::VFGT;    
                                end
                                5'b11000 : begin
                                    instruction_o.op  = ariane_pkg::VFCPKAB_S; 
                                    imm_select        = SIMM;      
                                    if (~RVF) illegal_instr = 1'b1; 
                                    
                                    unique case (instr.rvftype.vfmt)
                                        
                                        2'b00: begin
                                            if (~RVFVEC)            illegal_instr = 1'b1; 
                                            if (instr.rvftype.repl) illegal_instr = 1'b1; 
                                        end
                                        2'b01: begin
                                            if (~XF16ALTVEC) illegal_instr = 1'b1; 
                                        end
                                        2'b10: begin
                                            if (~XF16VEC) illegal_instr = 1'b1; 
                                        end
                                        2'b11: begin
                                            if (~XF8VEC) illegal_instr = 1'b1; 
                                        end
                                        default : illegal_instr = 1'b1;
                                    endcase
                                end
                                5'b11001 : begin
                                    instruction_o.op  = ariane_pkg::VFCPKCD_S; 
                                    imm_select        = SIMM;      
                                    if (~RVF) illegal_instr = 1'b1; 
                                    
                                    unique case (instr.rvftype.vfmt)
                                        
                                        2'b00: illegal_instr = 1'b1; 
                                        2'b01: illegal_instr = 1'b1; 
                                        2'b10: illegal_instr = 1'b1; 
                                        2'b11: begin
                                            if (~XF8VEC) illegal_instr = 1'b1; 
                                        end
                                        default : illegal_instr = 1'b1;
                                    endcase
                                end
                                5'b11010 : begin
                                    instruction_o.op  = ariane_pkg::VFCPKAB_D; 
                                    imm_select        = SIMM;      
                                    if (~RVD) illegal_instr = 1'b1; 
                                    
                                    unique case (instr.rvftype.vfmt)
                                        
                                        2'b00: begin
                                            if (~RVFVEC)            illegal_instr = 1'b1; 
                                            if (instr.rvftype.repl) illegal_instr = 1'b1; 
                                        end
                                        2'b01: begin
                                            if (~XF16ALTVEC) illegal_instr = 1'b1; 
                                        end
                                        2'b10: begin
                                            if (~XF16VEC) illegal_instr = 1'b1; 
                                        end
                                        2'b11: begin
                                            if (~XF8VEC) illegal_instr = 1'b1; 
                                        end
                                        default : illegal_instr = 1'b1;
                                    endcase
                                end
                                5'b11011 : begin
                                    instruction_o.op  = ariane_pkg::VFCPKCD_D; 
                                    imm_select        = SIMM;      
                                    if (~RVD) illegal_instr = 1'b1; 
                                    
                                    unique case (instr.rvftype.vfmt)
                                        
                                        2'b00: illegal_instr = 1'b1; 
                                        2'b01: illegal_instr = 1'b1; 
                                        2'b10: illegal_instr = 1'b1; 
                                        2'b11: begin
                                            if (~XF8VEC) illegal_instr = 1'b1; 
                                        end
                                        default : illegal_instr = 1'b1;
                                    endcase
                                end
                                default : illegal_instr = 1'b1;
                            endcase
                            
                            unique case (instr.rvftype.vfmt)
                                
                                2'b00: if (~RVFVEC)     illegal_instr = 1'b1;
                                2'b01: if (~XF16ALTVEC) illegal_instr = 1'b1;
                                2'b10: if (~XF16VEC)    illegal_instr = 1'b1;
                                2'b11: if (~XF8VEC)     illegal_instr = 1'b1;
                                default: illegal_instr = 1'b1;
                            endcase
                            
                            if (~allow_replication & instr.rvftype.repl) illegal_instr = 1'b1;
                            
                            if (check_fprm) begin
                                unique case (frm_i) inside 
                                    [3'b000:3'b100]: ; 
                                    default : illegal_instr = 1'b1;
                                endcase
                            end
                        end else begin 
                            illegal_instr = 1'b1;
                        end
                    
                    
                    
                    end else begin
                        instruction_o.fu  = (instr.rtype.funct7 == 7'b000_0001) ? MULT : ALU;
                        instruction_o.rs1 = instr.rtype.rs1;
                        instruction_o.rs2 = instr.rtype.rs2;
                        instruction_o.rd  = instr.rtype.rd;
                        unique case ({instr.rtype.funct7, instr.rtype.funct3})
                            {7'b000_0000, 3'b000}: instruction_o.op = ariane_pkg::ADD;   
                            {7'b010_0000, 3'b000}: instruction_o.op = ariane_pkg::SUB;   
                            {7'b000_0000, 3'b010}: instruction_o.op = ariane_pkg::SLTS;  
                            {7'b000_0000, 3'b011}: instruction_o.op = ariane_pkg::SLTU;  
                            {7'b000_0000, 3'b100}: instruction_o.op = ariane_pkg::XORL;  
                            {7'b000_0000, 3'b110}: instruction_o.op = ariane_pkg::ORL;   
                            {7'b000_0000, 3'b111}: instruction_o.op = ariane_pkg::ANDL;  
                            {7'b000_0000, 3'b001}: instruction_o.op = ariane_pkg::SLL;   
                            {7'b000_0000, 3'b101}: instruction_o.op = ariane_pkg::SRL;   
                            {7'b010_0000, 3'b101}: instruction_o.op = ariane_pkg::SRA;   
                            
                            {7'b000_0001, 3'b000}: instruction_o.op = ariane_pkg::MUL;
                            {7'b000_0001, 3'b001}: instruction_o.op = ariane_pkg::MULH;
                            {7'b000_0001, 3'b010}: instruction_o.op = ariane_pkg::MULHSU;
                            {7'b000_0001, 3'b011}: instruction_o.op = ariane_pkg::MULHU;
                            {7'b000_0001, 3'b100}: instruction_o.op = ariane_pkg::DIV;
                            {7'b000_0001, 3'b101}: instruction_o.op = ariane_pkg::DIVU;
                            {7'b000_0001, 3'b110}: instruction_o.op = ariane_pkg::REM;
                            {7'b000_0001, 3'b111}: instruction_o.op = ariane_pkg::REMU;
                            default: begin
                                illegal_instr = 1'b1;
                            end
                        endcase
                    end
                end
                
                
                
                riscv::OpcodeOp32: begin
                    instruction_o.fu  = (instr.rtype.funct7 == 7'b000_0001) ? MULT : ALU;
                    instruction_o.rs1[4:0] = instr.rtype.rs1;
                    instruction_o.rs2[4:0] = instr.rtype.rs2;
                    instruction_o.rd[4:0]  = instr.rtype.rd;
                      if (riscv::IS_XLEN64) begin
                        unique case ({instr.rtype.funct7, instr.rtype.funct3})
                            {7'b000_0000, 3'b000}: instruction_o.op = ariane_pkg::ADDW; 
                            {7'b010_0000, 3'b000}: instruction_o.op = ariane_pkg::SUBW; 
                            {7'b000_0000, 3'b001}: instruction_o.op = ariane_pkg::SLLW; 
                            {7'b000_0000, 3'b101}: instruction_o.op = ariane_pkg::SRLW; 
                            {7'b010_0000, 3'b101}: instruction_o.op = ariane_pkg::SRAW; 
                            
                            {7'b000_0001, 3'b000}: instruction_o.op = ariane_pkg::MULW;
                            {7'b000_0001, 3'b100}: instruction_o.op = ariane_pkg::DIVW;
                            {7'b000_0001, 3'b101}: instruction_o.op = ariane_pkg::DIVUW;
                            {7'b000_0001, 3'b110}: instruction_o.op = ariane_pkg::REMW;
                            {7'b000_0001, 3'b111}: instruction_o.op = ariane_pkg::REMUW;
                            default: illegal_instr = 1'b1;
                        endcase
                      end else illegal_instr = 1'b1;
                end
                
                
                
                riscv::OpcodeOpImm: begin
                    instruction_o.fu  = ALU;
                    imm_select = IIMM;
                    instruction_o.rs1[4:0] = instr.itype.rs1;
                    instruction_o.rd[4:0]  = instr.itype.rd;
                    unique case (instr.itype.funct3)
                        3'b000: instruction_o.op = ariane_pkg::ADD;   
                        3'b010: instruction_o.op = ariane_pkg::SLTS;  
                        3'b011: instruction_o.op = ariane_pkg::SLTU;  
                        3'b100: instruction_o.op = ariane_pkg::XORL;  
                        3'b110: instruction_o.op = ariane_pkg::ORL;   
                        3'b111: instruction_o.op = ariane_pkg::ANDL;  
                        3'b001: begin
                          instruction_o.op = ariane_pkg::SLL;  
                          if (instr.instr[31:26] != 6'b0)
                            illegal_instr = 1'b1;
                          if (instr.instr[25] != 1'b0 && riscv::XLEN==32) illegal_instr = 1'b1;
                        end
                        3'b101: begin
                            if (instr.instr[31:26] == 6'b0)
                                instruction_o.op = ariane_pkg::SRL;  
                            else if (instr.instr[31:26] == 6'b010_000)
                                instruction_o.op = ariane_pkg::SRA;  
                            else
                                illegal_instr = 1'b1;
                            if (instr.instr[25] != 1'b0 && riscv::XLEN==32) illegal_instr = 1'b1;
                        end
                    endcase
                end
                
                
                
                riscv::OpcodeOpImm32: begin
                    instruction_o.fu  = ALU;
                    imm_select = IIMM;
                    instruction_o.rs1[4:0] = instr.itype.rs1;
                    instruction_o.rd[4:0]  = instr.itype.rd;
                    if (riscv::IS_XLEN64)
                    unique case (instr.itype.funct3)
                        3'b000: instruction_o.op = ariane_pkg::ADDW;  
                        3'b001: begin
                          instruction_o.op = ariane_pkg::SLLW;  
                          if (instr.instr[31:25] != 7'b0)
                              illegal_instr = 1'b1;
                        end
                        3'b101: begin
                            if (instr.instr[31:25] == 7'b0)
                                instruction_o.op = ariane_pkg::SRLW;  
                            else if (instr.instr[31:25] == 7'b010_0000)
                                instruction_o.op = ariane_pkg::SRAW;  
                            else
                                illegal_instr = 1'b1;
                        end
                        default: illegal_instr = 1'b1;
                    endcase
                    else illegal_instr = 1'b1;
                end
                
                
                
                riscv::OpcodeStore: begin
                    instruction_o.fu  = STORE;
                    imm_select = SIMM;
                    instruction_o.rs1[4:0]  = instr.stype.rs1;
                    instruction_o.rs2[4:0]  = instr.stype.rs2;
                    
                    unique case (instr.stype.funct3)
                        3'b000: instruction_o.op  = ariane_pkg::SB;
                        3'b001: instruction_o.op  = ariane_pkg::SH;
                        3'b010: instruction_o.op  = ariane_pkg::SW;
                        3'b011: if (riscv::XLEN==64) instruction_o.op  = ariane_pkg::SD; 
                                else illegal_instr = 1'b1;
                        default: illegal_instr = 1'b1;
                    endcase
                end
                riscv::OpcodeLoad: begin
                    instruction_o.fu  = LOAD;
                    imm_select = IIMM;
                    instruction_o.rs1[4:0] = instr.itype.rs1;
                    instruction_o.rd[4:0]  = instr.itype.rd;
                    
                    unique case (instr.itype.funct3)
                        3'b000: instruction_o.op  = ariane_pkg::LB;
                        3'b001: instruction_o.op  = ariane_pkg::LH;
                        3'b010: instruction_o.op  = ariane_pkg::LW;
                        3'b100: instruction_o.op  = ariane_pkg::LBU;
                        3'b101: instruction_o.op  = ariane_pkg::LHU;
                        3'b110: instruction_o.op  = ariane_pkg::LWU;
                        3'b011: if (riscv::XLEN==64) instruction_o.op  = ariane_pkg::LD; 
                                else illegal_instr = 1'b1;
                        default: illegal_instr = 1'b1;
                    endcase
                end
                
                
                
                riscv::OpcodeStoreFp: begin
                    if (FP_PRESENT && fs_i != riscv::Off) begin 
                        instruction_o.fu  = STORE;
                        imm_select = SIMM;
                        instruction_o.rs1        = instr.stype.rs1;
                        instruction_o.rs2        = instr.stype.rs2;
                        
                        unique case (instr.stype.funct3)
                            
                            3'b000: if (XF8) instruction_o.op = ariane_pkg::FSB;
                                    else illegal_instr = 1'b1;
                            3'b001: if (XF16 | XF16ALT) instruction_o.op = ariane_pkg::FSH;
                                    else illegal_instr = 1'b1;
                            3'b010: if (RVF) instruction_o.op = ariane_pkg::FSW;
                                    else illegal_instr = 1'b1;
                            3'b011: if (RVD) instruction_o.op = ariane_pkg::FSD;
                                    else illegal_instr = 1'b1;
                            default: illegal_instr = 1'b1;
                        endcase
                    end else
                        illegal_instr = 1'b1;
                end
                riscv::OpcodeLoadFp: begin
                    if (FP_PRESENT && fs_i != riscv::Off) begin 
                        instruction_o.fu  = LOAD;
                        imm_select = IIMM;
                        instruction_o.rs1       = instr.itype.rs1;
                        instruction_o.rd        = instr.itype.rd;
                        
                        unique case (instr.itype.funct3)
                            
                            3'b000: if (XF8) instruction_o.op = ariane_pkg::FLB;
                                    else illegal_instr = 1'b1;
                            3'b001: if (XF16 | XF16ALT) instruction_o.op = ariane_pkg::FLH;
                                    else illegal_instr = 1'b1;
                            3'b010: if (RVF) instruction_o.op  = ariane_pkg::FLW;
                                    else illegal_instr = 1'b1;
                            3'b011: if (RVD) instruction_o.op  = ariane_pkg::FLD;
                                    else illegal_instr = 1'b1;
                            default: illegal_instr = 1'b1;
                        endcase
                    end else
                        illegal_instr = 1'b1;
                end
                
                
                
                riscv::OpcodeMadd,
                riscv::OpcodeMsub,
                riscv::OpcodeNmsub,
                riscv::OpcodeNmadd: begin
                    if (FP_PRESENT && fs_i != riscv::Off) begin 
                        instruction_o.fu  = FPU;
                        instruction_o.rs1 = instr.r4type.rs1;
                        instruction_o.rs2 = instr.r4type.rs2;
                        instruction_o.rd  = instr.r4type.rd;
                        imm_select        = RS3; 
                        check_fprm        = 1'b1;
                        
                        unique case (instr.r4type.opcode)
                            default:      instruction_o.op = ariane_pkg::FMADD;  
                            riscv::OpcodeMsub:  instruction_o.op = ariane_pkg::FMSUB;  
                            riscv::OpcodeNmsub: instruction_o.op = ariane_pkg::FNMSUB; 
                            riscv::OpcodeNmadd: instruction_o.op = ariane_pkg::FNMADD; 
                        endcase
                        
                        unique case (instr.r4type.funct2)
                            
                            2'b00: if (~RVF)             illegal_instr = 1'b1;
                            2'b01: if (~RVD)             illegal_instr = 1'b1;
                            2'b10: if (~XF16 & ~XF16ALT) illegal_instr = 1'b1;
                            2'b11: if (~XF8)             illegal_instr = 1'b1;
                            default: illegal_instr = 1'b1;
                        endcase
                        
                        if (check_fprm) begin
                            unique case (instr.rftype.rm) inside
                                [3'b000:3'b100]: ; 
                                3'b101: begin      
                                    if (~XF16ALT || instr.rftype.fmt != 2'b10)
                                        illegal_instr = 1'b1;
                                    unique case (frm_i) inside 
                                        [3'b000:3'b100]: ; 
                                        default : illegal_instr = 1'b1;
                                    endcase
                                end
                                3'b111: begin
                                    
                                    unique case (frm_i) inside
                                        [3'b000:3'b100]: ; 
                                        default : illegal_instr = 1'b1;
                                    endcase
                                end
                                default : illegal_instr = 1'b1;
                            endcase
                        end
                    end else begin
                        illegal_instr = 1'b1;
                    end
                end
                riscv::OpcodeOpFp: begin
                    if (FP_PRESENT && fs_i != riscv::Off) begin 
                        instruction_o.fu  = FPU;
                        instruction_o.rs1 = instr.rftype.rs1;
                        instruction_o.rs2 = instr.rftype.rs2;
                        instruction_o.rd  = instr.rftype.rd;
                        check_fprm        = 1'b1;
                        
                        unique case (instr.rftype.funct5)
                            5'b00000: begin
                                instruction_o.op  = ariane_pkg::FADD;             
                                instruction_o.rs1 = '0;               
                                instruction_o.rs2 = instr.rftype.rs1; 
                                imm_select        = IIMM;             
                            end
                            5'b00001: begin
                                instruction_o.op  = ariane_pkg::FSUB;  
                                instruction_o.rs1 = '0;               
                                instruction_o.rs2 = instr.rftype.rs1; 
                                imm_select        = IIMM;             
                            end
                            5'b00010: instruction_o.op = ariane_pkg::FMUL;  
                            5'b00011: instruction_o.op = ariane_pkg::FDIV;  
                            5'b01011: begin
                                instruction_o.op = ariane_pkg::FSQRT; 
                                
                                if (instr.rftype.rs2 != 5'b00000) illegal_instr = 1'b1;
                            end
                            5'b00100: begin
                                instruction_o.op = ariane_pkg::FSGNJ; 
                                check_fprm       = 1'b0;  
                                if (XF16ALT) begin        
                                    if (!(instr.rftype.rm inside {[3'b000:3'b010], [3'b100:3'b110]}))
                                        illegal_instr = 1'b1;
                                end else begin
                                    if (!(instr.rftype.rm inside {[3'b000:3'b010]}))
                                        illegal_instr = 1'b1;
                                end
                            end
                            5'b00101: begin
                                instruction_o.op = ariane_pkg::FMIN_MAX; 
                                check_fprm       = 1'b0;     
                                if (XF16ALT) begin           
                                    if (!(instr.rftype.rm inside {[3'b000:3'b001], [3'b100:3'b101]}))
                                        illegal_instr = 1'b1;
                                end else begin
                                    if (!(instr.rftype.rm inside {[3'b000:3'b001]}))
                                        illegal_instr = 1'b1;
                                end
                            end
                            5'b01000: begin
                                instruction_o.op  = ariane_pkg::FCVT_F2F; 
                                instruction_o.rs2 = instr.rvftype.rs1; 
                                imm_select        = IIMM;     
                                if (instr.rftype.rs2[24:23]) illegal_instr = 1'b1; 
                                
                                unique case (instr.rftype.rs2[22:20])
                                    
                                    3'b000: if (~RVF)     illegal_instr = 1'b1;
                                    3'b001: if (~RVD)     illegal_instr = 1'b1;
                                    3'b010: if (~XF16)    illegal_instr = 1'b1;
                                    3'b110: if (~XF16ALT) illegal_instr = 1'b1;
                                    3'b011: if (~XF8)     illegal_instr = 1'b1;
                                    default: illegal_instr = 1'b1;
                                endcase
                            end
                            5'b10100: begin
                                instruction_o.op = ariane_pkg::FCMP; 
                                check_fprm       = 1'b0; 
                                if (XF16ALT) begin       
                                    if (!(instr.rftype.rm inside {[3'b000:3'b010], [3'b100:3'b110]}))
                                        illegal_instr = 1'b1;
                                end else begin
                                    if (!(instr.rftype.rm inside {[3'b000:3'b010]}))
                                        illegal_instr = 1'b1;
                                end
                            end
                            5'b11000: begin
                                instruction_o.op = ariane_pkg::FCVT_F2I; 
                                imm_select       = IIMM;     
                                if (instr.rftype.rs2[24:22]) illegal_instr = 1'b1; 
                            end
                            5'b11010: begin
                                instruction_o.op = ariane_pkg::FCVT_I2F;  
                                imm_select       = IIMM;     
                                if (instr.rftype.rs2[24:22]) illegal_instr = 1'b1; 
                            end
                            5'b11100: begin
                                instruction_o.rs2 = instr.rftype.rs1; 
                                check_fprm        = 1'b0; 
                                if (instr.rftype.rm == 3'b000 || (XF16ALT && instr.rftype.rm == 3'b100)) 
                                    instruction_o.op = ariane_pkg::FMV_F2X;       
                                else if (instr.rftype.rm == 3'b001 || (XF16ALT && instr.rftype.rm == 3'b101)) 
                                    instruction_o.op = ariane_pkg::FCLASS; 
                                else illegal_instr = 1'b1;
                                
                                if (instr.rftype.rs2 != 5'b00000) illegal_instr = 1'b1;
                            end
                            5'b11110: begin
                                instruction_o.op = ariane_pkg::FMV_X2F;   
                                instruction_o.rs2 = instr.rftype.rs1; 
                                check_fprm       = 1'b0; 
                                if (!(instr.rftype.rm == 3'b000 || (XF16ALT && instr.rftype.rm == 3'b100)))
                                    illegal_instr = 1'b1;
                                
                                if (instr.rftype.rs2 != 5'b00000) illegal_instr = 1'b1;
                            end
                            default : illegal_instr = 1'b1;
                        endcase
                        
                        unique case (instr.rftype.fmt)
                            
                            2'b00: if (~RVF)             illegal_instr = 1'b1;
                            2'b01: if (~RVD)             illegal_instr = 1'b1;
                            2'b10: if (~XF16 & ~XF16ALT) illegal_instr = 1'b1;
                            2'b11: if (~XF8)             illegal_instr = 1'b1;
                            default: illegal_instr = 1'b1;
                        endcase
                        
                        if (check_fprm) begin
                            unique case (instr.rftype.rm) inside
                                [3'b000:3'b100]: ; 
                                3'b101: begin      
                                    if (~XF16ALT || instr.rftype.fmt != 2'b10)
                                        illegal_instr = 1'b1;
                                    unique case (frm_i) inside 
                                        [3'b000:3'b100]: ; 
                                        default : illegal_instr = 1'b1;
                                    endcase
                                end
                                3'b111: begin
                                    
                                    unique case (frm_i) inside
                                        [3'b000:3'b100]: ; 
                                        default : illegal_instr = 1'b1;
                                    endcase
                                end
                                default : illegal_instr = 1'b1;
                            endcase
                        end
                    end else begin
                        illegal_instr = 1'b1;
                    end
                end
                
                
                
                riscv::OpcodeAmo: begin
                    
                    instruction_o.fu  = STORE;
                    instruction_o.rs1[4:0] = instr.atype.rs1;
                    instruction_o.rs2[4:0] = instr.atype.rs2;
                    instruction_o.rd[4:0]  = instr.atype.rd;
                    
                    
                    if (RVA && instr.stype.funct3 == 3'h2) begin
                        unique case (instr.instr[31:27])
                            5'h0:  instruction_o.op = ariane_pkg::AMO_ADDW;
                            5'h1:  instruction_o.op = ariane_pkg::AMO_SWAPW;
                            5'h2: begin
                                instruction_o.op = ariane_pkg::AMO_LRW;
                                if (instr.atype.rs2 != 0) illegal_instr = 1'b1;
                            end
                            5'h3:  instruction_o.op = ariane_pkg::AMO_SCW;
                            5'h4:  instruction_o.op = ariane_pkg::AMO_XORW;
                            5'h8:  instruction_o.op = ariane_pkg::AMO_ORW;
                            5'hC:  instruction_o.op = ariane_pkg::AMO_ANDW;
                            5'h10: instruction_o.op = ariane_pkg::AMO_MINW;
                            5'h14: instruction_o.op = ariane_pkg::AMO_MAXW;
                            5'h18: instruction_o.op = ariane_pkg::AMO_MINWU;
                            5'h1C: instruction_o.op = ariane_pkg::AMO_MAXWU;
                            default: illegal_instr = 1'b1;
                        endcase
                    
                    end else if (RVA && instr.stype.funct3 == 3'h3) begin
                        unique case (instr.instr[31:27])
                            5'h0:  instruction_o.op = ariane_pkg::AMO_ADDD;
                            5'h1:  instruction_o.op = ariane_pkg::AMO_SWAPD;
                            5'h2: begin
                                instruction_o.op = ariane_pkg::AMO_LRD;
                                if (instr.atype.rs2 != 0) illegal_instr = 1'b1;
                            end
                            5'h3:  instruction_o.op = ariane_pkg::AMO_SCD;
                            5'h4:  instruction_o.op = ariane_pkg::AMO_XORD;
                            5'h8:  instruction_o.op = ariane_pkg::AMO_ORD;
                            5'hC:  instruction_o.op = ariane_pkg::AMO_ANDD;
                            5'h10: instruction_o.op = ariane_pkg::AMO_MIND;
                            5'h14: instruction_o.op = ariane_pkg::AMO_MAXD;
                            5'h18: instruction_o.op = ariane_pkg::AMO_MINDU;
                            5'h1C: instruction_o.op = ariane_pkg::AMO_MAXDU;
                            default: illegal_instr = 1'b1;
                        endcase
                    end else begin
                        illegal_instr = 1'b1;
                    end
                end
                
                
                
                riscv::OpcodeBranch: begin
                    imm_select              = SBIMM;
                    instruction_o.fu        = CTRL_FLOW;
                    instruction_o.rs1[4:0]  = instr.stype.rs1;
                    instruction_o.rs2[4:0]  = instr.stype.rs2;
                    is_control_flow_instr_o = 1'b1;
                    case (instr.stype.funct3)
                        3'b000: instruction_o.op = ariane_pkg::EQ;
                        3'b001: instruction_o.op = ariane_pkg::NE;
                        3'b100: instruction_o.op = ariane_pkg::LTS;
                        3'b101: instruction_o.op = ariane_pkg::GES;
                        3'b110: instruction_o.op = ariane_pkg::LTU;
                        3'b111: instruction_o.op = ariane_pkg::GEU;
                        default: begin
                            is_control_flow_instr_o = 1'b0;
                            illegal_instr           = 1'b1;
                        end
                    endcase
                end
                
                riscv::OpcodeJalr: begin
                    instruction_o.fu        = CTRL_FLOW;
                    instruction_o.op        = ariane_pkg::JALR;
                    instruction_o.rs1[4:0]  = instr.itype.rs1;
                    imm_select              = IIMM;
                    instruction_o.rd[4:0]   = instr.itype.rd;
                    is_control_flow_instr_o = 1'b1;
                    
                    if (instr.itype.funct3 != 3'b0) illegal_instr = 1'b1;
                end
                
                riscv::OpcodeJal: begin
                    instruction_o.fu        = CTRL_FLOW;
                    imm_select              = JIMM;
                    instruction_o.rd[4:0]   = instr.utype.rd;
                    is_control_flow_instr_o = 1'b1;
                end
                riscv::OpcodeAuipc: begin
                    instruction_o.fu      = ALU;
                    imm_select            = UIMM;
                    instruction_o.use_pc  = 1'b1;
                    instruction_o.rd[4:0] = instr.utype.rd;
                end
                riscv::OpcodeLui: begin
                    imm_select            = UIMM;
                    instruction_o.fu      = ALU;
                    instruction_o.rd[4:0] = instr.utype.rd;
                end
                default: illegal_instr = 1'b1;
            endcase
        end
    end
    
    
    
    always_comb begin : sign_extend
        imm_i_type  = { {riscv::XLEN-12{instruction_i[31]}}, instruction_i[31:20] };
        imm_s_type  = { {riscv::XLEN-12{instruction_i[31]}}, instruction_i[31:25], instruction_i[11:7] };
        imm_sb_type = { {riscv::XLEN-13{instruction_i[31]}}, instruction_i[31], instruction_i[7], instruction_i[30:25], instruction_i[11:8], 1'b0 };
        imm_u_type  = { {riscv::XLEN-32{instruction_i[31]}}, instruction_i[31:12], 12'b0 }; 
        imm_uj_type = { {riscv::XLEN-20{instruction_i[31]}}, instruction_i[19:12], instruction_i[20], instruction_i[30:21], 1'b0 };
        imm_bi_type = { {riscv::XLEN-5{instruction_i[24]}}, instruction_i[24:20] };
        
        
        case (imm_select)
            IIMM: begin
                instruction_o.result = imm_i_type;
                instruction_o.use_imm = 1'b1;
            end
            SIMM: begin
                instruction_o.result = imm_s_type;
                instruction_o.use_imm = 1'b1;
            end
            SBIMM: begin
                instruction_o.result = imm_sb_type;
                instruction_o.use_imm = 1'b1;
            end
            UIMM: begin
                instruction_o.result = imm_u_type;
                instruction_o.use_imm = 1'b1;
            end
            JIMM: begin
                instruction_o.result = imm_uj_type;
                instruction_o.use_imm = 1'b1;
            end
            RS3: begin
                
                instruction_o.result = {{riscv::XLEN-5{1'b0}}, instr.r4type.rs3};
                instruction_o.use_imm = 1'b0;
            end
            default: begin
                instruction_o.result = {riscv::XLEN{1'b0}};
                instruction_o.use_imm = 1'b0;
            end
        endcase
    end
    
    
    
    riscv::xlen_t interrupt_cause;
    
    assign instruction_o.valid   = instruction_o.ex.valid;
    always_comb begin : exception_handling
        interrupt_cause       = '0;
        instruction_o.ex      = ex_i;
        
        
        if (~ex_i.valid) begin
            
            
            instruction_o.ex.tval  = (is_compressed_i) ? {{riscv::XLEN-16{1'b0}}, compressed_instr_i} : {{riscv::XLEN-32{1'b0}}, instruction_i};
            
            
            
            
            if (illegal_instr || is_illegal_i) begin
                instruction_o.ex.valid = 1'b1;
                
                instruction_o.ex.cause = riscv::ILLEGAL_INSTR;
            
            end else if (ecall) begin
                
                instruction_o.ex.valid = 1'b1;
                
                case (priv_lvl_i)
                    riscv::PRIV_LVL_M: instruction_o.ex.cause = riscv::ENV_CALL_MMODE;
                    riscv::PRIV_LVL_S: instruction_o.ex.cause = riscv::ENV_CALL_SMODE;
                    riscv::PRIV_LVL_U: instruction_o.ex.cause = riscv::ENV_CALL_UMODE;
                    default:; 
                endcase
            end else if (ebreak) begin
                
                instruction_o.ex.valid = 1'b1;
                
                instruction_o.ex.cause = riscv::BREAKPOINT;
            end
            
            
            
            
            
            
            
            
            if (irq_ctrl_i.mie[riscv::S_TIMER_INTERRUPT[$clog2(riscv::XLEN)-1:0]] && irq_ctrl_i.mip[riscv::S_TIMER_INTERRUPT[$clog2(riscv::XLEN)-1:0]]) begin
                interrupt_cause = riscv::S_TIMER_INTERRUPT;
            end
            
            if (irq_ctrl_i.mie[riscv::S_SW_INTERRUPT[$clog2(riscv::XLEN)-1:0]] && irq_ctrl_i.mip[riscv::S_SW_INTERRUPT[$clog2(riscv::XLEN)-1:0]]) begin
                interrupt_cause = riscv::S_SW_INTERRUPT;
            end
            
            
            
            if (irq_ctrl_i.mie[riscv::S_EXT_INTERRUPT[$clog2(riscv::XLEN)-1:0]] && (irq_ctrl_i.mip[riscv::S_EXT_INTERRUPT[$clog2(riscv::XLEN)-1:0]] | irq_i[ariane_pkg::SupervisorIrq])) begin
                interrupt_cause = riscv::S_EXT_INTERRUPT;
            end
            
            if (irq_ctrl_i.mip[riscv::M_TIMER_INTERRUPT[$clog2(riscv::XLEN)-1:0]] && irq_ctrl_i.mie[riscv::M_TIMER_INTERRUPT[$clog2(riscv::XLEN)-1:0]]) begin
                interrupt_cause = riscv::M_TIMER_INTERRUPT;
            end
            
            if (irq_ctrl_i.mip[riscv::M_SW_INTERRUPT[$clog2(riscv::XLEN)-1:0]] && irq_ctrl_i.mie[riscv::M_SW_INTERRUPT[$clog2(riscv::XLEN)-1:0]]) begin
                interrupt_cause = riscv::M_SW_INTERRUPT;
            end
            
            if (irq_ctrl_i.mip[riscv::M_EXT_INTERRUPT[$clog2(riscv::XLEN)-1:0]] && irq_ctrl_i.mie[riscv::M_EXT_INTERRUPT[$clog2(riscv::XLEN)-1:0]]) begin
                interrupt_cause = riscv::M_EXT_INTERRUPT;
            end
            if (interrupt_cause[riscv::XLEN-1] && irq_ctrl_i.global_enable) begin
                
                
                
                if (irq_ctrl_i.mideleg[interrupt_cause[$clog2(riscv::XLEN)-1:0]]) begin
                    if ((irq_ctrl_i.sie && priv_lvl_i == riscv::PRIV_LVL_S) || priv_lvl_i == riscv::PRIV_LVL_U) begin
                        instruction_o.ex.valid = 1'b1;
                        instruction_o.ex.cause = interrupt_cause;
                    end
                end else begin
                    instruction_o.ex.valid = 1'b1;
                    instruction_o.ex.cause = interrupt_cause;
                end
            end
        end
        
        if (debug_req_i && !debug_mode_i) begin
          instruction_o.ex.valid = 1'b1;
          instruction_o.ex.cause = riscv::DEBUG_REQUEST;
        end
    end
endmodule
module ex_stage import ariane_pkg::*; #(
    parameter int unsigned ASID_WIDTH = 1,
    parameter ariane_pkg::ariane_cfg_t ArianeCfg = ariane_pkg::ArianeDefaultConfig
) (
    input  logic                                   clk_i,    
    input  logic                                   rst_ni,   
    input  logic                                   flush_i,
    input  logic                                   debug_mode_i,
    input  logic [riscv::VLEN-1:0]                 rs1_forwarding_i,
    input  logic [riscv::VLEN-1:0]                 rs2_forwarding_i,
    input  fu_data_t                               fu_data_i,
    input  logic [riscv::VLEN-1:0]                 pc_i,                  
    input  logic                                   is_compressed_instr_i, 
                                                                          
    
    output riscv::xlen_t                           flu_result_o,
    output logic [TRANS_ID_BITS-1:0]               flu_trans_id_o,        
    output exception_t                             flu_exception_o,
    output logic                                   flu_ready_o,           
    output logic                                   flu_valid_o,           
    
    
    input  logic                                   alu_valid_i,           
    
    input  logic                                   branch_valid_i,        
    input  branchpredict_sbe_t                     branch_predict_i,
    output bp_resolve_t                            resolved_branch_o,     
    output logic                                   resolve_branch_o,      
    
    input  logic                                   csr_valid_i,
    output logic [11:0]                            csr_addr_o,
    input  logic                                   csr_commit_i,
    
    input  logic                                   mult_valid_i,      
    
    output logic                                   lsu_ready_o,        
    input  logic                                   lsu_valid_i,        
    output logic                                   load_valid_o,
    output riscv::xlen_t                           load_result_o,
    output logic [TRANS_ID_BITS-1:0]               load_trans_id_o,
    output exception_t                             load_exception_o,
    output logic                                   store_valid_o,
    output riscv::xlen_t                           store_result_o,
    output logic [TRANS_ID_BITS-1:0]               store_trans_id_o,
    output exception_t                             store_exception_o,
    input  logic                                   lsu_commit_i,
    output logic                                   lsu_commit_ready_o, 
    input  logic [TRANS_ID_BITS-1:0]               commit_tran_id_i,
    output logic                                   no_st_pending_o,
    input  logic                                   amo_valid_commit_i,
    
    output logic                                   fpu_ready_o,      
    input  logic                                   fpu_valid_i,      
    input  logic [1:0]                             fpu_fmt_i,        
    input  logic [2:0]                             fpu_rm_i,         
    input  logic [2:0]                             fpu_frm_i,        
    input  logic [6:0]                             fpu_prec_i,       
    output logic [TRANS_ID_BITS-1:0]               fpu_trans_id_o,
    output riscv::xlen_t                           fpu_result_o,
    output logic                                   fpu_valid_o,
    output exception_t                             fpu_exception_o,
    
    input  logic                                   enable_translation_i,
    input  logic                                   en_ld_st_translation_i,
    input  logic                                   flush_tlb_i,
    input  riscv::priv_lvl_t                       priv_lvl_i,
    input  riscv::priv_lvl_t                       ld_st_priv_lvl_i,
    input  logic                                   sum_i,
    input  logic                                   mxr_i,
    input  logic [riscv::PPNW-1:0]                 satp_ppn_i,
    input  logic [ASID_WIDTH-1:0]                  asid_i,
    
    input  icache_areq_o_t                         icache_areq_i,
    output icache_areq_i_t                         icache_areq_o,
    
    input  dcache_req_o_t [2:0]                    dcache_req_ports_i,
    output dcache_req_i_t [2:0]                    dcache_req_ports_o,
    input  logic                                   dcache_wbuffer_empty_i,
    input  logic                                   dcache_wbuffer_not_ni_i,
    output amo_req_t                               amo_req_o,          
    input  amo_resp_t                              amo_resp_i,         
    
    output logic                                   itlb_miss_o,
    output logic                                   dtlb_miss_o,
    
    input  riscv::pmpcfg_t [15:0]                  pmpcfg_i,
    input  logic[15:0][riscv::PLEN-3:0]            pmpaddr_i
);
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    logic current_instruction_is_sfence_vma;
    
    
    logic [ASID_WIDTH-1:0] asid_to_be_flushed;
    logic [riscv::VLEN-1:0] vaddr_to_be_flushed;
    
    logic alu_branch_res; 
    riscv::xlen_t alu_result, csr_result, mult_result;
    logic [riscv::VLEN-1:0] branch_result;
    logic csr_ready, mult_ready;
    logic [TRANS_ID_BITS-1:0] mult_trans_id;
    logic mult_valid;
    
    
    fu_data_t alu_data;
    assign alu_data = (alu_valid_i | branch_valid_i) ? fu_data_i  : '0;
    alu alu_i (
        .clk_i,
        .rst_ni,
        .fu_data_i        ( alu_data       ),
        .result_o         ( alu_result     ),
        .alu_branch_res_o ( alu_branch_res )
    );
    
    
    
    branch_unit branch_unit_i (
        .clk_i,
        .rst_ni,
        .debug_mode_i,
        .fu_data_i,
        .pc_i,
        .is_compressed_instr_i,
        
        .fu_valid_i ( alu_valid_i || lsu_valid_i || csr_valid_i || mult_valid_i || fpu_valid_i ) ,
        .branch_valid_i,
        .branch_comp_res_i ( alu_branch_res ),
        .branch_result_o   ( branch_result ),
        .branch_predict_i,
        .resolved_branch_o,
        .resolve_branch_o,
        .branch_exception_o ( flu_exception_o )
    );
    
    csr_buffer csr_buffer_i (
        .clk_i,
        .rst_ni,
        .flush_i,
        .fu_data_i,
        .csr_valid_i,
        .csr_ready_o    ( csr_ready    ),
        .csr_result_o   ( csr_result   ),
        .csr_commit_i,
        .csr_addr_o
    );
    assign flu_valid_o = alu_valid_i | branch_valid_i | csr_valid_i | mult_valid;
    
    always_comb begin
        
        flu_result_o = {{riscv::XLEN-riscv::VLEN{1'b0}}, branch_result};
        flu_trans_id_o = fu_data_i.trans_id;
        
        if (alu_valid_i) begin
            flu_result_o = alu_result;
        
        end else if (csr_valid_i) begin
            flu_result_o = csr_result;
        end else if (mult_valid) begin
            flu_result_o = mult_result;
            flu_trans_id_o = mult_trans_id;
        end
    end
    
    always_comb begin
        flu_ready_o = csr_ready & mult_ready;
    end
    
    fu_data_t mult_data;
    
    assign mult_data  = mult_valid_i ? fu_data_i  : '0;
    mult i_mult (
        .clk_i,
        .rst_ni,
        .flush_i,
        .mult_valid_i,
        .fu_data_i       ( mult_data     ),
        .result_o        ( mult_result   ),
        .mult_valid_o    ( mult_valid    ),
        .mult_ready_o    ( mult_ready    ),
        .mult_trans_id_o ( mult_trans_id )
    );
    
    
    
    generate
        if (FP_PRESENT) begin : fpu_gen
            fu_data_t fpu_data;
            assign fpu_data  = fpu_valid_i ? fu_data_i  : '0;
            fpu_wrap fpu_i (
                .clk_i,
                .rst_ni,
                .flush_i,
                .fpu_valid_i,
                .fpu_ready_o,
                .fu_data_i ( fpu_data ),
                .fpu_fmt_i,
                .fpu_rm_i,
                .fpu_frm_i,
                .fpu_prec_i,
                .fpu_trans_id_o,
                .result_o ( fpu_result_o ),
                .fpu_valid_o,
                .fpu_exception_o
            );
        end else begin : no_fpu_gen
            assign fpu_ready_o     = '0;
            assign fpu_trans_id_o  = '0;
            assign fpu_result_o    = '0;
            assign fpu_valid_o     = '0;
            assign fpu_exception_o = '0;
        end
    endgenerate
    
    
    
    fu_data_t lsu_data;
    assign lsu_data  = lsu_valid_i ? fu_data_i  : '0;
    load_store_unit #(
        .ASID_WIDTH ( ASID_WIDTH ),
        .ArianeCfg ( ArianeCfg )
    ) lsu_i (
        .clk_i,
        .rst_ni,
        .flush_i,
        .no_st_pending_o,
        .fu_data_i             ( lsu_data ),
        .lsu_ready_o,
        .lsu_valid_i,
        .load_trans_id_o,
        .load_result_o,
        .load_valid_o,
        .load_exception_o,
        .store_trans_id_o,
        .store_result_o,
        .store_valid_o,
        .store_exception_o,
        .commit_i              ( lsu_commit_i       ),
        .commit_ready_o        ( lsu_commit_ready_o ),
        .commit_tran_id_i,
        .enable_translation_i,
        .en_ld_st_translation_i,
        .icache_areq_i,
        .icache_areq_o,
        .priv_lvl_i,
        .ld_st_priv_lvl_i,
        .sum_i,
        .mxr_i,
        .satp_ppn_i,
        .asid_i,
        .asid_to_be_flushed_i (asid_to_be_flushed),
        .vaddr_to_be_flushed_i (vaddr_to_be_flushed),
        .flush_tlb_i,
        .itlb_miss_o,
        .dtlb_miss_o,
        .dcache_req_ports_i,
        .dcache_req_ports_o,
        .dcache_wbuffer_empty_i,
        .dcache_wbuffer_not_ni_i,
        .amo_valid_commit_i,
        .amo_req_o,
        .amo_resp_i,
        .pmpcfg_i,
        .pmpaddr_i
    );
	always_ff @(posedge clk_i or negedge rst_ni) begin
	    if (~rst_ni) begin
          current_instruction_is_sfence_vma <= 1'b0;
		  end else begin
          if (flush_i) begin
              current_instruction_is_sfence_vma <= 1'b0;
          end else if ((fu_data_i.operator == SFENCE_VMA) && csr_valid_i) begin
              current_instruction_is_sfence_vma <= 1'b1;
          end
      end
  end
  
	always_ff @(posedge clk_i or negedge rst_ni) begin
		if (~rst_ni) begin
		    asid_to_be_flushed  <= '0;
			  vaddr_to_be_flushed <=  '0;
    
		end else if ((~current_instruction_is_sfence_vma) && (~((fu_data_i.operator == SFENCE_VMA) && csr_valid_i))) begin
			  vaddr_to_be_flushed <=  rs1_forwarding_i;
			  asid_to_be_flushed  <= rs2_forwarding_i[ASID_WIDTH-1:0];
		end
	end
endmodule
module instr_realign import ariane_pkg::*; (
    input  logic                              clk_i,
    input  logic                              rst_ni,
    input  logic                              flush_i,
    input  logic                              valid_i,
    output logic                              serving_unaligned_o, 
    input  logic [riscv::VLEN-1:0]            address_i,
    input  logic [FETCH_WIDTH-1:0]            data_i,
    output logic [INSTR_PER_FETCH-1:0]        valid_o,
    output logic [INSTR_PER_FETCH-1:0][riscv::VLEN-1:0]  addr_o,
    output logic [INSTR_PER_FETCH-1:0][31:0]  instr_o
);
    
    logic [3:0] instr_is_compressed;
    for (genvar i = 0; i < INSTR_PER_FETCH; i ++) begin
        
        assign instr_is_compressed[i] = ~&data_i[i * 16 +: 2];
    end
    
    logic [15:0] unaligned_instr_d,   unaligned_instr_q;
    
    logic        unaligned_d,         unaligned_q;
    
    logic [riscv::VLEN-1:0] unaligned_address_d, unaligned_address_q;
    
    assign serving_unaligned_o = unaligned_q;
    
    if (FETCH_WIDTH == 32) begin : realign_bp_32
        always_comb begin : re_align
            unaligned_d = unaligned_q;
            unaligned_address_d = {address_i[riscv::VLEN-1:2], 2'b10};
            unaligned_instr_d = data_i[31:16];
            valid_o[0] = valid_i;
            instr_o[0] = (unaligned_q) ? {data_i[15:0], unaligned_instr_q} : data_i[31:0];
            addr_o[0]  = (unaligned_q) ? unaligned_address_q : address_i;
            valid_o[1] = 1'b0;
            instr_o[1] = '0;
            addr_o[1]  = {address_i[riscv::VLEN-1:2], 2'b10};
            
            if (instr_is_compressed[0] || unaligned_q) begin
                
                
                
                
                
                
                if (instr_is_compressed[1]) begin
                    unaligned_d = 1'b0;
                    valid_o[1] = valid_i;
                    instr_o[1] = {16'b0, data_i[31:16]};
                end else begin
                    
                    unaligned_d = 1'b1;
                    unaligned_instr_d = data_i[31:16];
                    unaligned_address_d = {address_i[riscv::VLEN-1:2], 2'b10};
                end
            end 
            
            
            if (valid_i && address_i[1]) begin
                
                if (!instr_is_compressed[0]) begin
                    valid_o = '0;
                    unaligned_d = 1'b1;
                    unaligned_address_d = {address_i[riscv::VLEN-1:2], 2'b10};
                    unaligned_instr_d = data_i[15:0];
                
                end else begin
                    valid_o = 1'b1;
                end
            end
        end
    
    end else if (FETCH_WIDTH == 64) begin : realign_bp_64
        initial begin
          $error("Not propperly implemented");
        end
        always_comb begin : re_align
            unaligned_d = unaligned_q;
            unaligned_address_d = unaligned_address_q;
            unaligned_instr_d = unaligned_instr_q;
            valid_o    = '0;
            valid_o[0] = valid_i;
            instr_o[0] = data_i[31:0];
            addr_o[0]  = address_i;
            instr_o[1] = '0;
            addr_o[1]  = {address_i[riscv::VLEN-1:3], 3'b010};
            instr_o[2] = {16'b0, data_i[47:32]};
            addr_o[2]  = {address_i[riscv::VLEN-1:3], 3'b100};
            instr_o[3] = {16'b0, data_i[63:48]};
            addr_o[3]  = {address_i[riscv::VLEN-1:3], 3'b110};
            
            if (unaligned_q) begin
                instr_o[0] = {data_i[15:0], unaligned_instr_q};
                addr_o[0] = unaligned_address_q;
                
                
                
                
                
                
                
                
                
                
                if (instr_is_compressed[1]) begin
                    instr_o[1] = {16'b0, data_i[31:16]};
                    valid_o[1] = valid_i;
                    if (instr_is_compressed[2]) begin
                        if (instr_is_compressed[3]) begin
                            unaligned_d = 1'b0;
                            valid_o[3] = valid_i;
                        end else begin
                            
                        end
                    end else begin
                        unaligned_d = 1'b0;
                        instr_o[2] = data_i[63:32];
                        valid_o[2] = valid_i;
                    end
                
                end else begin
                    instr_o[1] = data_i[47:16];
                    valid_o[1] = valid_i;
                    addr_o[2] = {address_i[riscv::VLEN-1:3], 3'b110};
                    if (instr_is_compressed[2]) begin
                        unaligned_d = 1'b0;
                        instr_o[2] = {16'b0, data_i[63:48]};
                        valid_o[2] = valid_i;
                    end else begin
                        
                    end
                end
            end else if (instr_is_compressed[0]) begin 
                
                
                
                
                
                
                
                if (instr_is_compressed[1]) begin
                    instr_o[1] = {16'b0, data_i[31:16]};
                    valid_o[1] = valid_i;
                    if (instr_is_compressed[2]) begin
                        valid_o[2] = valid_i;
                        if (instr_is_compressed[3]) begin
                            valid_o[3] = valid_i;
                        end else begin
                            
                            unaligned_d = 1'b1;
                            unaligned_instr_d = data_i[63:48];
                            unaligned_address_d = addr_o[3];
                        end
                    end else begin
                        instr_o[2] = data_i[63:32];
                        valid_o[2] = valid_i;
                    end
                
                end else begin
                    instr_o[1] = data_i[47:16];
                    valid_o[1] = valid_i;
                    addr_o[2] = {address_i[riscv::VLEN-1:3], 3'b110};
                    if (instr_is_compressed[3]) begin
                        instr_o[2] = data_i[63:48];
                        valid_o[2] = valid_i;
                    end else begin
                        unaligned_d = 1'b1;
                        unaligned_instr_d = data_i[63:48];
                        unaligned_address_d = addr_o[2];
                    end
                end
            
            
            
            
            
            
            end else begin
                addr_o[1] = {address_i[riscv::VLEN-1:3], 3'b100};
                if (instr_is_compressed[2]) begin
                    instr_o[1] = {16'b0, data_i[47:32]};
                    valid_o[1] = valid_i;
                    addr_o[2] = {address_i[riscv::VLEN-1:3], 3'b110};
                    if (instr_is_compressed[3]) begin
                        
                        valid_o[2] = valid_i;
                        addr_o[2] = {16'b0, data_i[63:48]};
                    end else begin
                        
                        unaligned_d = 1'b1;
                        unaligned_instr_d = data_i[63:48];
                        unaligned_address_d = addr_o[2];
                    end
                end else begin
                    
                    instr_o[1] = data_i[63:32];
                    valid_o[1] = valid_i;
                end
            end
            
            
            
            
            case (address_i[2:1])
                
                
                2'b01: begin
                    
                    
                    
                    
                    
                    
                    
                    addr_o[0] = {address_i[riscv::VLEN-1:3], 3'b010};
                    if (instr_is_compressed[1]) begin
                        instr_o[0] = {16'b0, data_i[31:16]};
                        valid_o[0] = valid_i;
                        if (instr_is_compressed[2]) begin
                            valid_o[1] = valid_i;
                            instr_o[1] = {16'b0, data_i[47:32]};
                            addr_o[1] = {address_i[riscv::VLEN-1:3], 3'b100};
                            if (instr_is_compressed[3]) begin
                                instr_o[2] = {16'b0, data_i[63:48]};
                                addr_o[2] = {address_i[riscv::VLEN-1:3], 3'b110};
                                valid_o[2] = valid_i;
                            end else begin
                                
                                unaligned_d = 1'b1;
                                unaligned_instr_d = data_i[63:48];
                                unaligned_address_d = addr_o[3];
                            end
                        end else begin
                            instr_o[1] = data_i[63:32];
                            addr_o[1] = {address_i[riscv::VLEN-1:3], 3'b100};
                            valid_o[1] = valid_i;
                        end
                    
                    end else begin
                        instr_o[0] = data_i[47:16];
                        valid_o[0] = valid_i;
                        addr_o[1] = {address_i[riscv::VLEN-1:3], 3'b110};
                        if (instr_is_compressed[3]) begin
                            instr_o[1] = data_i[63:48];
                            valid_o[1] = valid_i;
                        end else begin
                            unaligned_d = 1'b1;
                            unaligned_instr_d = data_i[63:48];
                            unaligned_address_d = addr_o[1];
                        end
                    end
                end
                2'b10: begin
                    valid_o = '0;
                    
                    
                    
                    
                    
                    if (instr_is_compressed[2]) begin
                        valid_o[0] = valid_i;
                        instr_o[0] = data_i[47:32];
                        
                        if (instr_is_compressed[3]) begin
                            valid_o[1] = valid_i;
                            instr_o[1] = data_i[63:48];
                        
                        end else begin
                            unaligned_d = 1'b1;
                            unaligned_address_d = {address_i[riscv::VLEN-1:3], 3'b110};
                            unaligned_instr_d = data_i[63:48];
                        end
                    
                    end else begin
                        valid_o[0] = valid_i;
                        instr_o[0] = data_i[63:32];
                        addr_o[0] = address_i;
                    end
                end
                
                
                2'b11: begin
                    valid_o = '0;
                    if (!instr_is_compressed[3]) begin
                        unaligned_d = 1'b1;
                        unaligned_address_d = {address_i[riscv::VLEN-1:3], 3'b110};
                        unaligned_instr_d = data_i[63:48];
                    end else begin
                        valid_o[3] = valid_i;
                    end
                end
            endcase
        end
    end
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (~rst_ni) begin
            unaligned_q         <= 1'b0;
            unaligned_address_q <= '0;
            unaligned_instr_q   <= '0;
        end else begin
            if (valid_i) begin
                unaligned_address_q <= unaligned_address_d;
                unaligned_instr_q   <= unaligned_instr_d;
            end
            if (flush_i) begin
                unaligned_q <= 1'b0;
            end else if (valid_i) begin
                unaligned_q <= unaligned_d;
            end
        end
    end
endmodule
module btb #(
    parameter int NR_ENTRIES = 8
)(
    input  logic                        clk_i,           
    input  logic                        rst_ni,          
    input  logic                        flush_i,         
    input  logic                        debug_mode_i,
    input  logic [riscv::VLEN-1:0]      vpc_i,           
    input  ariane_pkg::btb_update_t     btb_update_i,    
    output ariane_pkg::btb_prediction_t [ariane_pkg::INSTR_PER_FETCH-1:0] btb_prediction_o 
);
    
    localparam OFFSET = 1;
    
    localparam NR_ROWS = NR_ENTRIES / ariane_pkg::INSTR_PER_FETCH;
    
    localparam ROW_ADDR_BITS = $clog2(ariane_pkg::INSTR_PER_FETCH);
    
    localparam PREDICTION_BITS = $clog2(NR_ROWS) + OFFSET + ROW_ADDR_BITS;
    
    localparam ANTIALIAS_BITS = 8;
    
    unread i_unread (.d_i(|vpc_i));
    
    
    ariane_pkg::btb_prediction_t btb_d [NR_ROWS-1:0][ariane_pkg::INSTR_PER_FETCH-1:0],
                                 btb_q [NR_ROWS-1:0][ariane_pkg::INSTR_PER_FETCH-1:0];
    logic [$clog2(NR_ROWS)-1:0]  index, update_pc;
    logic [ROW_ADDR_BITS-1:0]    update_row_index;
    assign index     = vpc_i[PREDICTION_BITS - 1:ROW_ADDR_BITS + OFFSET];
    assign update_pc = btb_update_i.pc[PREDICTION_BITS - 1:ROW_ADDR_BITS + OFFSET];
    assign update_row_index = btb_update_i.pc[ROW_ADDR_BITS + OFFSET - 1:OFFSET];
    
    for (genvar i = 0; i < ariane_pkg::INSTR_PER_FETCH; i++) begin : gen_btb_output
        assign btb_prediction_o[i] = btb_q[index][i]; 
    end
    
    
    
    
    always_comb begin : update_branch_predict
        btb_d = btb_q;
        if (btb_update_i.valid && !debug_mode_i) begin
            btb_d[update_pc][update_row_index].valid = 1'b1;
            
            btb_d[update_pc][update_row_index].target_address = btb_update_i.target_address;
        end
    end
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (!rst_ni) begin
            
            for (int i = 0; i < NR_ROWS; i++)
                btb_q[i] <= '{default: 0};
        end else begin
            
            if (flush_i) begin
                for (int i = 0; i < NR_ROWS; i++) begin
                    for (int j = 0; j < ariane_pkg::INSTR_PER_FETCH; j++) begin
                        btb_q[i][j].valid <=  1'b0;
                    end
                end
            end else begin
                btb_q <=  btb_d;
            end
        end
    end
endmodule
module bht #(
    parameter int unsigned NR_ENTRIES = 1024
)(
    input  logic                        clk_i,
    input  logic                        rst_ni,
    input  logic                        flush_i,
    input  logic                        debug_mode_i,
    input  logic [riscv::VLEN-1:0]      vpc_i,
    input  ariane_pkg::bht_update_t     bht_update_i,
    
    output ariane_pkg::bht_prediction_t [ariane_pkg::INSTR_PER_FETCH-1:0] bht_prediction_o
);
    
    localparam OFFSET = 1;
    
    localparam NR_ROWS = NR_ENTRIES / ariane_pkg::INSTR_PER_FETCH;
    
    localparam ROW_ADDR_BITS = $clog2(ariane_pkg::INSTR_PER_FETCH);
    
    localparam PREDICTION_BITS = $clog2(NR_ROWS) + OFFSET + ROW_ADDR_BITS;
    
    unread i_unread (.d_i(|vpc_i));
    struct packed {
        logic       valid;
        logic [1:0] saturation_counter;
    } bht_d[NR_ROWS-1:0][ariane_pkg::INSTR_PER_FETCH-1:0], bht_q[NR_ROWS-1:0][ariane_pkg::INSTR_PER_FETCH-1:0];
    logic [$clog2(NR_ROWS)-1:0]  index, update_pc;
    logic [ROW_ADDR_BITS-1:0]    update_row_index;
    logic [1:0]                  saturation_counter;
    assign index     = vpc_i[PREDICTION_BITS - 1:ROW_ADDR_BITS + OFFSET];
    assign update_pc = bht_update_i.pc[PREDICTION_BITS - 1:ROW_ADDR_BITS + OFFSET];
    assign update_row_index = bht_update_i.pc[ROW_ADDR_BITS + OFFSET - 1:OFFSET];
    
    for (genvar i = 0; i < ariane_pkg::INSTR_PER_FETCH; i++) begin : gen_bht_output
        assign bht_prediction_o[i].valid = bht_q[index][i].valid;
        assign bht_prediction_o[i].taken = bht_q[index][i].saturation_counter[1] == 1'b1;
    end
    always_comb begin : update_bht
        bht_d = bht_q;
        saturation_counter = bht_q[update_pc][update_row_index].saturation_counter;
        if (bht_update_i.valid && !debug_mode_i) begin
            bht_d[update_pc][update_row_index].valid = 1'b1;
            if (saturation_counter == 2'b11) begin
                
                if (!bht_update_i.taken)
                    bht_d[update_pc][update_row_index].saturation_counter = saturation_counter - 1;
            
            end else if (saturation_counter == 2'b00) begin
                
                if (bht_update_i.taken)
                    bht_d[update_pc][update_row_index].saturation_counter = saturation_counter + 1;
            end else begin 
                if (bht_update_i.taken)
                    bht_d[update_pc][update_row_index].saturation_counter = saturation_counter + 1;
                else
                    bht_d[update_pc][update_row_index].saturation_counter = saturation_counter - 1;
            end
        end
    end
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (!rst_ni) begin
            for (int unsigned i = 0; i < NR_ROWS; i++) begin
                for (int j = 0; j < ariane_pkg::INSTR_PER_FETCH; j++) begin
                    bht_q[i][j] <= '0;
                end
            end
        end else begin
            
            if (flush_i) begin
                for (int i = 0; i < NR_ROWS; i++) begin
                    for (int j = 0; j < ariane_pkg::INSTR_PER_FETCH; j++) begin
                        bht_q[i][j].valid <=  1'b0;
                        bht_q[i][j].saturation_counter <= 2'b10;
                    end
                end
            end else begin
                bht_q <= bht_d;
            end
        end
    end
endmodule
module ras #(
    parameter int unsigned DEPTH = 2
)(
    input  logic             clk_i,
    input  logic             rst_ni,
    input  logic             flush_i,
    input  logic             push_i,
    input  logic             pop_i,
    input  logic [riscv::VLEN-1:0]      data_i,
    output ariane_pkg::ras_t data_o
);
    ariane_pkg::ras_t [DEPTH-1:0] stack_d, stack_q;
    assign data_o = stack_q[0];
    always_comb begin
        stack_d = stack_q;
        
        if (push_i) begin
            stack_d[0].ra = data_i;
            
            stack_d[0].valid = 1'b1;
            stack_d[DEPTH-1:1] = stack_q[DEPTH-2:0];
        end
        if (pop_i) begin
            stack_d[DEPTH-2:0] = stack_q[DEPTH-1:1];
            
            stack_d[DEPTH-1].valid = 1'b0;
            stack_d[DEPTH-1].ra = 'b0;
        end
        
        
        if (pop_i && push_i) begin
           stack_d = stack_q;
           stack_d[0].ra = data_i;
           stack_d[0].valid = 1'b1;
        end
        if (flush_i) begin
          stack_d = '0;
        end
    end
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (~rst_ni) begin
            stack_q <= '0;
        end else begin
            stack_q <= stack_d;
        end
    end
endmodule
module instr_scan (
    input  logic [31:0] instr_i,        
    output logic        rvi_return_o,
    output logic        rvi_call_o,
    output logic        rvi_branch_o,
    output logic        rvi_jalr_o,
    output logic        rvi_jump_o,
    output logic [riscv::VLEN-1:0] rvi_imm_o,
    output logic        rvc_branch_o,
    output logic        rvc_jump_o,
    output logic        rvc_jr_o,
    output logic        rvc_return_o,
    output logic        rvc_jalr_o,
    output logic        rvc_call_o,
    output logic [riscv::VLEN-1:0] rvc_imm_o
);
    logic is_rvc;
    assign is_rvc     = (instr_i[1:0] != 2'b11);
    logic rv32_rvc_jal;
    assign rv32_rvc_jal = (riscv::XLEN == 32) & ((instr_i[15:13] == riscv::OpcodeC1Jal) & is_rvc & (instr_i[1:0] == riscv::OpcodeC1));
    
    assign rvi_return_o = rvi_jalr_o & ((instr_i[19:15] == 5'd1) | instr_i[19:15] == 5'd5)
                                     & (instr_i[19:15] != instr_i[11:7]);
    
    assign rvi_call_o   = (rvi_jalr_o | rvi_jump_o) & ((instr_i[11:7] == 5'd1) | instr_i[11:7] == 5'd5);
    
    assign rvi_imm_o    = (instr_i[3]) ? ariane_pkg::uj_imm(instr_i) : ariane_pkg::sb_imm(instr_i);
    assign rvi_branch_o = (instr_i[6:0] == riscv::OpcodeBranch);
    assign rvi_jalr_o   = (instr_i[6:0] == riscv::OpcodeJalr);
    assign rvi_jump_o   = (instr_i[6:0] == riscv::OpcodeJal);
    
    assign rvc_jump_o   = ((instr_i[15:13] == riscv::OpcodeC1J) & is_rvc & (instr_i[1:0] == riscv::OpcodeC1)) | rv32_rvc_jal;
    
    logic is_jal_r;
    assign is_jal_r     = (instr_i[15:13] == riscv::OpcodeC2JalrMvAdd)
                        & (instr_i[6:2] == 5'b00000)
                        & (instr_i[1:0] == riscv::OpcodeC2)
                        & is_rvc;
    assign rvc_jr_o     = is_jal_r & ~instr_i[12];
    
    assign rvc_jalr_o   = is_jal_r & instr_i[12];
    assign rvc_call_o   = rvc_jalr_o | rv32_rvc_jal;
    assign rvc_branch_o = ((instr_i[15:13] == riscv::OpcodeC1Beqz) | (instr_i[15:13] == riscv::OpcodeC1Bnez))
                        & (instr_i[1:0] == riscv::OpcodeC1)
                        & is_rvc;
    
    assign rvc_return_o = ((instr_i[11:7] == 5'd1) | (instr_i[11:7] == 5'd5))  & rvc_jr_o ;
    
    assign rvc_imm_o    = (instr_i[14]) ? {{56+riscv::VLEN-64{instr_i[12]}}, instr_i[6:5], instr_i[2], instr_i[11:10], instr_i[4:3], 1'b0}
                                       : {{53+riscv::VLEN-64{instr_i[12]}}, instr_i[8], instr_i[10:9], instr_i[6], instr_i[7], instr_i[2], instr_i[11], instr_i[5:3], 1'b0};
endmodule
module instr_queue (
  input  logic                                               clk_i,
  input  logic                                               rst_ni,
  input  logic                                               flush_i,
  input  logic [ariane_pkg::INSTR_PER_FETCH-1:0][31:0]       instr_i,
  input  logic [ariane_pkg::INSTR_PER_FETCH-1:0][riscv::VLEN-1:0] addr_i,
  input  logic [ariane_pkg::INSTR_PER_FETCH-1:0]             valid_i,
  output logic                                               ready_o,
  output logic [ariane_pkg::INSTR_PER_FETCH-1:0]             consumed_o,
  
  input  ariane_pkg::frontend_exception_t                    exception_i,
  input  logic [riscv::VLEN-1:0]                             exception_addr_i,
  
  input  logic [riscv::VLEN-1:0]                             predict_address_i,
  input  ariane_pkg::cf_t  [ariane_pkg::INSTR_PER_FETCH-1:0] cf_type_i,
  
  output logic                                               replay_o,
  output logic [riscv::VLEN-1:0]                             replay_addr_o, 
  
  output ariane_pkg::fetch_entry_t                           fetch_entry_o,
  output logic                                               fetch_entry_valid_o,
  input  logic                                               fetch_entry_ready_i
);
  typedef struct packed {
    logic [31:0]     instr; 
    ariane_pkg::cf_t cf;    
    ariane_pkg::frontend_exception_t ex;    
    logic [riscv::VLEN-1:0] ex_vaddr;       
  } instr_data_t;
  logic [$clog2(ariane_pkg::INSTR_PER_FETCH)-1:0] branch_index;
  
  logic [ariane_pkg::INSTR_PER_FETCH-1:0]
        [$clog2(ariane_pkg::FETCH_FIFO_DEPTH)-1:0] instr_queue_usage;
  instr_data_t [ariane_pkg::INSTR_PER_FETCH-1:0]   instr_data_in, instr_data_out;
  logic [ariane_pkg::INSTR_PER_FETCH-1:0]          push_instr, push_instr_fifo;
  logic [ariane_pkg::INSTR_PER_FETCH-1:0]          pop_instr;
  logic [ariane_pkg::INSTR_PER_FETCH-1:0]          instr_queue_full;
  logic [ariane_pkg::INSTR_PER_FETCH-1:0]          instr_queue_empty;
  logic instr_overflow;
  
  logic [$clog2(ariane_pkg::FETCH_FIFO_DEPTH)-1:0] address_queue_usage;
  logic [riscv::VLEN-1:0] address_out;
  logic pop_address;
  logic push_address;
  logic full_address;
  logic empty_address;
  logic address_overflow;
  
  logic [$clog2(ariane_pkg::INSTR_PER_FETCH)-1:0] idx_is_d, idx_is_q;
  
  
  logic [ariane_pkg::INSTR_PER_FETCH-1:0] idx_ds_d, idx_ds_q;
  logic [riscv::VLEN-1:0] pc_d, pc_q; 
  logic reset_address_d, reset_address_q; 
  logic [ariane_pkg::INSTR_PER_FETCH*2-2:0] branch_mask_extended;
  logic [ariane_pkg::INSTR_PER_FETCH-1:0] branch_mask;
  logic branch_empty;
  logic [ariane_pkg::INSTR_PER_FETCH-1:0] taken;
  
  logic [$clog2(ariane_pkg::INSTR_PER_FETCH):0] popcount;
  logic [$clog2(ariane_pkg::INSTR_PER_FETCH)-1:0] shamt;
  logic [ariane_pkg::INSTR_PER_FETCH-1:0] valid;
  logic [ariane_pkg::INSTR_PER_FETCH*2-1:0] consumed_extended;
  
  logic [ariane_pkg::INSTR_PER_FETCH*2-1:0] fifo_pos_extended;
  logic [ariane_pkg::INSTR_PER_FETCH-1:0] fifo_pos;
  logic [ariane_pkg::INSTR_PER_FETCH*2-1:0][31:0] instr;
  ariane_pkg::cf_t [ariane_pkg::INSTR_PER_FETCH*2-1:0] cf;
  
  logic [ariane_pkg::INSTR_PER_FETCH-1:0] instr_overflow_fifo;
  assign ready_o = ~(|instr_queue_full) & ~full_address;
  for (genvar i = 0; i < ariane_pkg::INSTR_PER_FETCH; i++) begin : gen_unpack_taken
    assign taken[i] = cf_type_i[i] != ariane_pkg::NoCF;
  end
  
  lzc #(
    .WIDTH   ( ariane_pkg::INSTR_PER_FETCH ),
    .MODE    ( 0                           ) 
  ) i_lzc_branch_index (
    .in_i    ( taken          ), 
    .cnt_o   ( branch_index   ), 
    .empty_o ( branch_empty   )
  );
  
  
  
  
  
  
  assign branch_mask_extended = {{{ariane_pkg::INSTR_PER_FETCH-1}{1'b0}}, {{ariane_pkg::INSTR_PER_FETCH}{1'b1}}} << branch_index;
  assign branch_mask = branch_mask_extended[ariane_pkg::INSTR_PER_FETCH * 2 - 2:ariane_pkg::INSTR_PER_FETCH - 1];
  
  assign valid = valid_i & branch_mask;
  
  assign consumed_extended = {push_instr_fifo, push_instr_fifo} >> idx_is_q;
  assign consumed_o = consumed_extended[ariane_pkg::INSTR_PER_FETCH-1:0];
  
  popcount #(
    .INPUT_WIDTH   ( ariane_pkg::INSTR_PER_FETCH )
  ) i_popcount (
    .data_i     ( push_instr_fifo ),
    .popcount_o ( popcount        )
  );
  assign shamt = popcount[$bits(shamt)-1:0];
  
  assign idx_is_d = idx_is_q + shamt;
  
  
  
  
  assign fifo_pos_extended = { valid, valid } << idx_is_q;
  
  assign fifo_pos = fifo_pos_extended[ariane_pkg::INSTR_PER_FETCH*2-1:ariane_pkg::INSTR_PER_FETCH];
  
  
  assign push_instr = fifo_pos & ~instr_queue_full;
  
  for (genvar i = 0; i < ariane_pkg::INSTR_PER_FETCH; i++) begin : gen_duplicate_instr_input
    assign instr[i] = instr_i[i];
    assign instr[i + ariane_pkg::INSTR_PER_FETCH] = instr_i[i];
    assign cf[i] = cf_type_i[i];
    assign cf[i + ariane_pkg::INSTR_PER_FETCH] = cf_type_i[i];
  end
  
  for (genvar i = 0; i < ariane_pkg::INSTR_PER_FETCH; i++) begin : gen_fifo_input_select
    
    assign instr_data_in[i].instr = instr[i + idx_is_q];
    assign instr_data_in[i].cf = cf[i + idx_is_q];
    assign instr_data_in[i].ex = exception_i; 
    assign instr_data_in[i].ex_vaddr = exception_addr_i;
    
  end
  
  
  
  
  
  
  
  
  assign instr_overflow_fifo = instr_queue_full & fifo_pos;
  assign instr_overflow = |instr_overflow_fifo; 
  assign address_overflow = full_address & push_address;
  assign replay_o = instr_overflow | address_overflow;
  
  
  
  
  assign replay_addr_o = (address_overflow) ? addr_i[0] : addr_i[shamt];
  
  
  
  
  assign fetch_entry_valid_o = ~(&instr_queue_empty);
  always_comb begin
    idx_ds_d = idx_ds_q;
    pop_instr = '0;
    
    fetch_entry_o.instruction = '0;
    fetch_entry_o.address = pc_q;
    fetch_entry_o.ex.valid = 1'b0;
    fetch_entry_o.ex.cause = '0;
    fetch_entry_o.ex.tval = '0;
    fetch_entry_o.branch_predict.predict_address = address_out;
    fetch_entry_o.branch_predict.cf = ariane_pkg::NoCF;
    
    for (int unsigned i = 0; i < ariane_pkg::INSTR_PER_FETCH; i++) begin
      if (idx_ds_q[i]) begin
        if (instr_data_out[i].ex == ariane_pkg::FE_INSTR_ACCESS_FAULT) begin
            fetch_entry_o.ex.cause = riscv::INSTR_ACCESS_FAULT;
        end else begin
            fetch_entry_o.ex.cause = riscv::INSTR_PAGE_FAULT;
        end
        fetch_entry_o.instruction = instr_data_out[i].instr;
        fetch_entry_o.ex.valid = instr_data_out[i].ex != ariane_pkg::FE_NONE;
        fetch_entry_o.ex.tval  = {{64-riscv::VLEN{1'b0}}, instr_data_out[i].ex_vaddr};
        fetch_entry_o.branch_predict.cf = instr_data_out[i].cf;
        pop_instr[i] = fetch_entry_valid_o & fetch_entry_ready_i;
      end
    end
    
    if (fetch_entry_ready_i) begin
      idx_ds_d = {idx_ds_q[ariane_pkg::INSTR_PER_FETCH-2:0], idx_ds_q[ariane_pkg::INSTR_PER_FETCH-1]};
    end
  end
  
  
  assign pop_address = ((fetch_entry_o.branch_predict.cf != ariane_pkg::NoCF) & |pop_instr);
  
  
  
  always_comb begin
    pc_d = pc_q;
    reset_address_d = flush_i ? 1'b1 : reset_address_q;
    if (fetch_entry_ready_i) begin
      
      
      pc_d =  pc_q + ((fetch_entry_o.instruction[1:0] != 2'b11) ? 'd2 : 'd4);
    end
    if (pop_address) pc_d = address_out;
      
    if (valid_i[0] && reset_address_q) begin
      
      pc_d = addr_i[0];
      reset_address_d = 1'b0;
    end
  end
  
  for (genvar i = 0; i < ariane_pkg::INSTR_PER_FETCH; i++) begin : gen_instr_fifo
    
    assign push_instr_fifo[i] = push_instr[i] & ~address_overflow;
    fifo_v3 #(
      .DEPTH      ( ariane_pkg::FETCH_FIFO_DEPTH ),
      .dtype      ( instr_data_t                 )
    ) i_fifo_instr_data (
      .clk_i      ( clk_i                ),
      .rst_ni     ( rst_ni               ),
      .flush_i    ( flush_i              ),
      .testmode_i ( 1'b0                 ),
      .full_o     ( instr_queue_full[i]  ),
      .empty_o    ( instr_queue_empty[i] ),
      .usage_o    ( instr_queue_usage[i] ),
      .data_i     ( instr_data_in[i]     ),
      .push_i     ( push_instr_fifo[i]   ),
      .data_o     ( instr_data_out[i]    ),
      .pop_i      ( pop_instr[i]         )
    );
  end
  
  
  always_comb begin
    push_address = 1'b0;
    
    for (int i = 0; i < ariane_pkg::INSTR_PER_FETCH; i++) begin
      push_address |= push_instr[i] & (instr_data_in[i].cf != ariane_pkg::NoCF);
    end
  end
  fifo_v3 #(
    .DEPTH      ( ariane_pkg::FETCH_FIFO_DEPTH ), 
    .DATA_WIDTH ( riscv::VLEN                  )
  ) i_fifo_address (
    .clk_i      ( clk_i                        ),
    .rst_ni     ( rst_ni                       ),
    .flush_i    ( flush_i                      ),
    .testmode_i ( 1'b0                         ),
    .full_o     ( full_address                 ),
    .empty_o    ( empty_address                ),
    .usage_o    ( address_queue_usage          ),
    .data_i     ( predict_address_i            ),
    .push_i     ( push_address & ~full_address ),
    .data_o     ( address_out                  ),
    .pop_i      ( pop_address                  )
  );
  unread i_unread_address_fifo (.d_i(|{empty_address, address_queue_usage}));
  unread i_unread_branch_mask (.d_i(|branch_mask_extended));
  unread i_unread_lzc (.d_i(|{branch_empty}));
  unread i_unread_fifo_pos (.d_i(|fifo_pos_extended)); 
  unread i_unread_instr_fifo (.d_i(|instr_queue_usage));
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      idx_ds_q        <= 'b1;
      idx_is_q        <= '0;
      pc_q            <= '0;
      reset_address_q <= 1'b1;
    end else begin
      pc_q            <= pc_d;
      reset_address_q <= reset_address_d;
      if (flush_i) begin
          
          idx_ds_q        <= 'b1;
          
          idx_is_q        <= '0;
          reset_address_q <= 1'b1;
      end else begin
          idx_ds_q        <= idx_ds_d;
          idx_is_q        <= idx_is_d;
      end
    end
  end
  
  
  
  
endmodule
module frontend import ariane_pkg::*; #(
  parameter ariane_pkg::ariane_cfg_t ArianeCfg = ariane_pkg::ArianeDefaultConfig
) (
  input  logic               clk_i,              
  input  logic               rst_ni,             
  input  logic               flush_i,            
  input  logic               flush_bp_i,         
  input  logic               debug_mode_i,
  
  input  logic [riscv::VLEN-1:0]        boot_addr_i,
  
  
  input  bp_resolve_t        resolved_branch_i,  
  
  input  logic               set_pc_commit_i,    
  input  logic [riscv::VLEN-1:0] pc_commit_i,        
  
  input  logic [riscv::VLEN-1:0] epc_i,              
  input  logic               eret_i,             
  input  logic [riscv::VLEN-1:0] trap_vector_base_i, 
  input  logic               ex_valid_i,         
  input  logic               set_debug_pc_i,     
  
  output icache_dreq_i_t     icache_dreq_o,
  input  icache_dreq_o_t     icache_dreq_i,
  
  output fetch_entry_t       fetch_entry_o,       
  output logic               fetch_entry_valid_o, 
  input  logic               fetch_entry_ready_i  
);
    
    logic [FETCH_WIDTH-1:0] icache_data_q;
    logic                   icache_valid_q;
    ariane_pkg::frontend_exception_t icache_ex_valid_q;
    logic [riscv::VLEN-1:0] icache_vaddr_q;
    logic                   instr_queue_ready;
    logic [ariane_pkg::INSTR_PER_FETCH-1:0] instr_queue_consumed;
    
    btb_prediction_t        btb_q;
    bht_prediction_t        bht_q;
    
    logic                   if_ready;
    logic [riscv::VLEN-1:0] npc_d, npc_q; 
    
    logic                   npc_rst_load_q;
    logic                   replay;
    logic [riscv::VLEN-1:0] replay_addr;
    
    logic [$clog2(ariane_pkg::INSTR_PER_FETCH)-1:0] shamt;
    
    assign shamt = icache_dreq_i.vaddr[$clog2(ariane_pkg::INSTR_PER_FETCH):1];
    
    
    
    
    logic [INSTR_PER_FETCH-1:0]       rvi_return, rvi_call, rvi_branch,
                                      rvi_jalr, rvi_jump;
    logic [INSTR_PER_FETCH-1:0][riscv::VLEN-1:0] rvi_imm;
    
    logic [INSTR_PER_FETCH-1:0]       rvc_branch, rvc_jump, rvc_jr, rvc_return,
                                      rvc_jalr, rvc_call;
    logic [INSTR_PER_FETCH-1:0][riscv::VLEN-1:0] rvc_imm;
    
    logic [INSTR_PER_FETCH-1:0][31:0] instr;
    logic [INSTR_PER_FETCH-1:0][riscv::VLEN-1:0] addr;
    logic [INSTR_PER_FETCH-1:0]       instruction_valid;
    
    bht_prediction_t [INSTR_PER_FETCH-1:0] bht_prediction;
    btb_prediction_t [INSTR_PER_FETCH-1:0] btb_prediction;
    bht_prediction_t [INSTR_PER_FETCH-1:0] bht_prediction_shifted;
    btb_prediction_t [INSTR_PER_FETCH-1:0] btb_prediction_shifted;
    ras_t            ras_predict;
    
    logic            is_mispredict;
    logic            ras_push, ras_pop;
    logic [riscv::VLEN-1:0]     ras_update;
    
    logic [riscv::VLEN-1:0]                 predict_address;
    cf_t  [ariane_pkg::INSTR_PER_FETCH-1:0] cf_type;
    logic [ariane_pkg::INSTR_PER_FETCH-1:0] taken_rvi_cf;
    logic [ariane_pkg::INSTR_PER_FETCH-1:0] taken_rvc_cf;
    logic serving_unaligned;
    
    instr_realign i_instr_realign (
      .clk_i               ( clk_i                 ),
      .rst_ni              ( rst_ni                ),
      .flush_i             ( icache_dreq_o.kill_s2 ),
      .valid_i             ( icache_valid_q        ),
      .serving_unaligned_o ( serving_unaligned     ),
      .address_i           ( icache_vaddr_q        ),
      .data_i              ( icache_data_q         ),
      .valid_o             ( instruction_valid     ),
      .addr_o              ( addr                  ),
      .instr_o             ( instr                 )
    );
    
    
    
    
    
    
    assign bht_prediction_shifted[0] = (serving_unaligned) ? bht_q : bht_prediction[0];
    assign btb_prediction_shifted[0] = (serving_unaligned) ? btb_q : btb_prediction[0];
    
    
    for (genvar i = 1; i < INSTR_PER_FETCH; i++) begin : gen_prediction_address
      assign bht_prediction_shifted[i] = bht_prediction[addr[i][$clog2(INSTR_PER_FETCH):1]];
      assign btb_prediction_shifted[i] = btb_prediction[addr[i][$clog2(INSTR_PER_FETCH):1]];
    end
    
    
    logic bp_valid;
    logic [INSTR_PER_FETCH-1:0] is_branch;
    logic [INSTR_PER_FETCH-1:0] is_call;
    logic [INSTR_PER_FETCH-1:0] is_jump;
    logic [INSTR_PER_FETCH-1:0] is_return;
    logic [INSTR_PER_FETCH-1:0] is_jalr;
    for (genvar i = 0; i < INSTR_PER_FETCH; i++) begin
      
      assign is_branch[i] =  instruction_valid[i] & (rvi_branch[i] | rvc_branch[i]);
      
      assign is_call[i] = instruction_valid[i] & (rvi_call[i] | rvc_call[i]);
      
      assign is_return[i] = instruction_valid[i] & (rvi_return[i] | rvc_return[i]);
      
      assign is_jump[i] = instruction_valid[i] & (rvi_jump[i] | rvc_jump[i]);
      
      assign is_jalr[i] = instruction_valid[i] & ~is_return[i] & ~is_call[i] & (rvi_jalr[i] | rvc_jalr[i] | rvc_jr[i]);
    end
    
    always_comb begin
      taken_rvi_cf = '0;
      taken_rvc_cf = '0;
      predict_address = '0;
      for (int i = 0; i < INSTR_PER_FETCH; i++)  cf_type[i] = ariane_pkg::NoCF;
      ras_push = 1'b0;
      ras_pop = 1'b0;
      ras_update = '0;
      
      for (int i = INSTR_PER_FETCH - 1; i >= 0 ; i--) begin
        unique case ({is_branch[i], is_return[i], is_jump[i], is_jalr[i]})
          4'b0000:; 
          
          4'b0001: begin
            ras_pop = 1'b0;
            ras_push = 1'b0;
            if (btb_prediction_shifted[i].valid) begin
              predict_address = btb_prediction_shifted[i].target_address;
              cf_type[i] = ariane_pkg::JumpR;
            end
          end
          
          4'b0010: begin
            ras_pop = 1'b0;
            ras_push = 1'b0;
            taken_rvi_cf[i] = rvi_jump[i];
            taken_rvc_cf[i] = rvc_jump[i];
            cf_type[i] = ariane_pkg::Jump;
          end
          
          4'b0100: begin
            
            ras_pop = ras_predict.valid & instr_queue_consumed[i];
            ras_push = 1'b0;
            predict_address = ras_predict.ra;
            cf_type[i] = ariane_pkg::Return;
          end
          
          4'b1000: begin
            ras_pop = 1'b0;
            ras_push = 1'b0;
            
            if (bht_prediction_shifted[i].valid) begin
              taken_rvi_cf[i] = rvi_branch[i] & bht_prediction_shifted[i].taken;
              taken_rvc_cf[i] = rvc_branch[i] & bht_prediction_shifted[i].taken;
            
            end else begin
              
              taken_rvi_cf[i] = rvi_branch[i] & rvi_imm[i][riscv::VLEN-1];
              taken_rvc_cf[i] = rvc_branch[i] & rvc_imm[i][riscv::VLEN-1];
            end
            if (taken_rvi_cf[i] || taken_rvc_cf[i]) cf_type[i] = ariane_pkg::Branch;
          end
          default:;
            
        endcase
          
          
          if (is_call[i]) begin
            ras_push = instr_queue_consumed[i];
            ras_update = addr[i] + (rvc_call[i] ? 2 : 4);
          end
          
          if (taken_rvc_cf[i] || taken_rvi_cf[i]) begin
            predict_address = addr[i] + (taken_rvc_cf[i] ? rvc_imm[i] : rvi_imm[i]);
          end
      end
    end
    
    always_comb begin
      bp_valid = 1'b0;
      
      
      
      for (int i = 0; i < INSTR_PER_FETCH; i++) bp_valid |= ((cf_type[i] != NoCF & cf_type[i] != Return) | ((cf_type[i] == Return) & ras_predict.valid));
    end
    assign is_mispredict = resolved_branch_i.valid & resolved_branch_i.is_mispredict;
    
    assign icache_dreq_o.req = instr_queue_ready;
    assign if_ready = icache_dreq_i.ready & instr_queue_ready;
    
    
    
    
    assign icache_dreq_o.kill_s1 = is_mispredict | flush_i | replay;
    
    
    assign icache_dreq_o.kill_s2 = icache_dreq_o.kill_s1 | bp_valid;
    
    bht_update_t bht_update;
    btb_update_t btb_update;
    
    logic speculative_q,speculative_d;
    assign speculative_d = (speculative_q && !resolved_branch_i.valid || |is_branch || |is_return || |is_jalr) && !flush_i;
    assign icache_dreq_o.spec = speculative_d;
    assign bht_update.valid = resolved_branch_i.valid
                                & (resolved_branch_i.cf_type == ariane_pkg::Branch);
    assign bht_update.pc    = resolved_branch_i.pc;
    assign bht_update.taken = resolved_branch_i.is_taken;
    
    assign btb_update.valid = resolved_branch_i.valid
                                & resolved_branch_i.is_mispredict
                                & (resolved_branch_i.cf_type == ariane_pkg::JumpR);
    assign btb_update.pc    = resolved_branch_i.pc;
    assign btb_update.target_address = resolved_branch_i.target_address;
    
    
    
    
    
    
    
    
    
    
    
    
    always_comb begin : npc_select
      automatic logic [riscv::VLEN-1:0] fetch_address;
      
      
      
      
      
      
      if (npc_rst_load_q) begin
        npc_d         = boot_addr_i;
        fetch_address = boot_addr_i;
      end else begin
        fetch_address    = npc_q;
        
        npc_d            = npc_q;
      end
      
      if (bp_valid) begin
        fetch_address = predict_address;
        npc_d = predict_address;
      end
      
      if (if_ready) npc_d = {fetch_address[riscv::VLEN-1:2], 2'b0}  + 'h4;
      
      if (replay) npc_d = replay_addr;
      
      if (is_mispredict) npc_d = resolved_branch_i.target_address;
      
      if (eret_i) npc_d = epc_i;
      
      if (ex_valid_i) npc_d = trap_vector_base_i;
      
      
      
      
      
      
      
      if (set_pc_commit_i) npc_d = pc_commit_i + {{riscv::VLEN-3{1'b0}}, 3'b100};
      
      
      if (set_debug_pc_i) npc_d = ArianeCfg.DmBaseAddress[riscv::VLEN-1:0] + dm::HaltAddress[riscv::VLEN-1:0];
      icache_dreq_o.vaddr = fetch_address;
    end
    logic [FETCH_WIDTH-1:0] icache_data;
    
    assign icache_data = icache_dreq_i.data >> {shamt, 4'b0};
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        npc_rst_load_q    <= 1'b1;
        npc_q             <= '0;
        speculative_q     <= '0;
        icache_data_q     <= '0;
        icache_valid_q    <= 1'b0;
        icache_vaddr_q    <= 'b0;
        icache_ex_valid_q <= ariane_pkg::FE_NONE;
        btb_q             <= '0;
        bht_q             <= '0;
      end else begin
        npc_rst_load_q    <= 1'b0;
        npc_q             <= npc_d;
        speculative_q    <= speculative_d;
        icache_valid_q    <= icache_dreq_i.valid;
        if (icache_dreq_i.valid) begin
          icache_data_q        <= icache_data;
          icache_vaddr_q       <= icache_dreq_i.vaddr;
          
          if (icache_dreq_i.ex.cause == riscv::INSTR_PAGE_FAULT) begin
            icache_ex_valid_q <= ariane_pkg::FE_INSTR_PAGE_FAULT;
          end else if (icache_dreq_i.ex.cause == riscv::INSTR_ACCESS_FAULT) begin
            icache_ex_valid_q <= ariane_pkg::FE_INSTR_ACCESS_FAULT;
          end else icache_ex_valid_q <= ariane_pkg::FE_NONE;
          
          btb_q                <= btb_prediction[INSTR_PER_FETCH-1];
          bht_q                <= bht_prediction[INSTR_PER_FETCH-1];
        end
      end
    end
    ras #(
      .DEPTH  ( ArianeCfg.RASDepth  )
    ) i_ras (
      .clk_i,
      .rst_ni,
      .flush_i( flush_bp_i  ),
      .push_i ( ras_push    ),
      .pop_i  ( ras_pop     ),
      .data_i ( ras_update  ),
      .data_o ( ras_predict )
    );
    btb #(
      .NR_ENTRIES       ( ArianeCfg.BTBEntries   )
    ) i_btb (
      .clk_i,
      .rst_ni,
      .flush_i          ( flush_bp_i       ),
      .debug_mode_i,
      .vpc_i            ( icache_vaddr_q   ),
      .btb_update_i     ( btb_update       ),
      .btb_prediction_o ( btb_prediction   )
    );
    bht #(
      .NR_ENTRIES       ( ArianeCfg.BHTEntries   )
    ) i_bht (
      .clk_i,
      .rst_ni,
      .flush_i          ( flush_bp_i       ),
      .debug_mode_i,
      .vpc_i            ( icache_vaddr_q   ),
      .bht_update_i     ( bht_update       ),
      .bht_prediction_o ( bht_prediction   )
    );
    
    
    for (genvar i = 0; i < INSTR_PER_FETCH; i++) begin : gen_instr_scan
      instr_scan i_instr_scan (
        .instr_i      ( instr[i]      ),
        .rvi_return_o ( rvi_return[i] ),
        .rvi_call_o   ( rvi_call[i]   ),
        .rvi_branch_o ( rvi_branch[i] ),
        .rvi_jalr_o   ( rvi_jalr[i]   ),
        .rvi_jump_o   ( rvi_jump[i]   ),
        .rvi_imm_o    ( rvi_imm[i]    ),
        .rvc_branch_o ( rvc_branch[i] ),
        .rvc_jump_o   ( rvc_jump[i]   ),
        .rvc_jr_o     ( rvc_jr[i]     ),
        .rvc_return_o ( rvc_return[i] ),
        .rvc_jalr_o   ( rvc_jalr[i]   ),
        .rvc_call_o   ( rvc_call[i]   ),
        .rvc_imm_o    ( rvc_imm[i]    )
      );
    end
    instr_queue i_instr_queue (
      .clk_i               ( clk_i                ),
      .rst_ni              ( rst_ni               ),
      .flush_i             ( flush_i              ),
      .instr_i             ( instr                ), 
      .addr_i              ( addr                 ), 
      .exception_i         ( icache_ex_valid_q    ), 
      .exception_addr_i    ( icache_vaddr_q       ),
      .predict_address_i   ( predict_address      ),
      .cf_type_i           ( cf_type              ),
      .valid_i             ( instruction_valid    ), 
      .consumed_o          ( instr_queue_consumed ),
      .ready_o             ( instr_queue_ready    ),
      .replay_o            ( replay               ),
      .replay_addr_o       ( replay_addr          ),
      .fetch_entry_o       ( fetch_entry_o        ), 
      .fetch_entry_valid_o ( fetch_entry_valid_o  ), 
      .fetch_entry_ready_i ( fetch_entry_ready_i  )  
    );
    
    
    
    
endmodule
module id_stage (
    input  logic                          clk_i,
    input  logic                          rst_ni,
    input  logic                          flush_i,
    input  logic                          debug_req_i,
    
    input  ariane_pkg::fetch_entry_t      fetch_entry_i,
    input  logic                          fetch_entry_valid_i,
    output logic                          fetch_entry_ready_o, 
    
    output ariane_pkg::scoreboard_entry_t issue_entry_o,       
    output logic                          issue_entry_valid_o, 
    output logic                          is_ctrl_flow_o,      
    input  logic                          issue_instr_ack_i,   
    
    input  riscv::priv_lvl_t              priv_lvl_i,          
    input  riscv::xs_t                    fs_i,                
    input  logic [2:0]                    frm_i,               
    input  logic [1:0]                    irq_i,
    input  ariane_pkg::irq_ctrl_t         irq_ctrl_i,
    input  logic                          debug_mode_i,        
    input  logic                          tvm_i,
    input  logic                          tw_i,
    input  logic                          tsr_i
);
    
    struct packed {
        logic                          valid;
        ariane_pkg::scoreboard_entry_t sbe;
        logic                          is_ctrl_flow;
    } issue_n, issue_q;
    logic                            is_control_flow_instr;
    ariane_pkg::scoreboard_entry_t   decoded_instruction;
    logic                is_illegal;
    logic                [31:0] instruction;
    logic                is_compressed;
    
    
    
    compressed_decoder compressed_decoder_i (
        .instr_i                 ( fetch_entry_i.instruction   ),
        .instr_o                 ( instruction                 ),
        .illegal_instr_o         ( is_illegal                  ),
        .is_compressed_o         ( is_compressed               )
    );
    
    
    
    decoder decoder_i (
        .debug_req_i,
        .irq_ctrl_i,
        .irq_i,
        .pc_i                    ( fetch_entry_i.address           ),
        .is_compressed_i         ( is_compressed                   ),
        .is_illegal_i            ( is_illegal                      ),
        .instruction_i           ( instruction                     ),
        .compressed_instr_i      ( fetch_entry_i.instruction[15:0] ),
        .branch_predict_i        ( fetch_entry_i.branch_predict    ),
        .ex_i                    ( fetch_entry_i.ex                ),
        .priv_lvl_i              ( priv_lvl_i                      ),
        .debug_mode_i            ( debug_mode_i                    ),
        .fs_i,
        .frm_i,
        .tvm_i,
        .tw_i,
        .tsr_i,
        .instruction_o           ( decoded_instruction          ),
        .is_control_flow_instr_o ( is_control_flow_instr        )
    );
    
    
    
    assign issue_entry_o = issue_q.sbe;
    assign issue_entry_valid_o = issue_q.valid;
    assign is_ctrl_flow_o = issue_q.is_ctrl_flow;
    always_comb begin
        issue_n     = issue_q;
        fetch_entry_ready_o = 1'b0;
        
        if (issue_instr_ack_i)
            issue_n.valid = 1'b0;
        
        
        
        if ((!issue_q.valid || issue_instr_ack_i) && fetch_entry_valid_i) begin
            fetch_entry_ready_o = 1'b1;
            issue_n = '{1'b1, decoded_instruction, is_control_flow_instr};
        end
        
        if (flush_i)
            issue_n.valid = 1'b0;
    end
    
    
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if(~rst_ni) begin
            issue_q <= '0;
        end else begin
            issue_q <= issue_n;
        end
    end
endmodule
module issue_read_operands import ariane_pkg::*; #(
    parameter int unsigned NR_COMMIT_PORTS = 2
)(
    input  logic                                   clk_i,    
    input  logic                                   rst_ni,   
    
    input  logic                                   flush_i,
    
    input  scoreboard_entry_t                      issue_instr_i,
    input  logic                                   issue_instr_valid_i,
    output logic                                   issue_ack_o,
    
    output logic [REG_ADDR_SIZE-1:0]               rs1_o,
    input  riscv::xlen_t                           rs1_i,
    input  logic                                   rs1_valid_i,
    output logic [REG_ADDR_SIZE-1:0]               rs2_o,
    input  riscv::xlen_t                           rs2_i,
    input  logic                                   rs2_valid_i,
    output logic [REG_ADDR_SIZE-1:0]               rs3_o,
    input  logic [FLEN-1:0]                        rs3_i,
    input  logic                                   rs3_valid_i,
    
    input  fu_t [2**REG_ADDR_SIZE-1:0]             rd_clobber_gpr_i,
    input  fu_t [2**REG_ADDR_SIZE-1:0]             rd_clobber_fpr_i,
    
    output fu_data_t                               fu_data_o,
    output logic [riscv::VLEN-1:0]                 rs1_forwarding_o,  
    output logic [riscv::VLEN-1:0]                 rs2_forwarding_o,  
    output logic [riscv::VLEN-1:0]                 pc_o,
    output logic                                   is_compressed_instr_o,
    
    input  logic                                   flu_ready_i,      
    output logic                                   alu_valid_o,      
    
    output logic                                   branch_valid_o,   
    output branchpredict_sbe_t                     branch_predict_o,
    
    input  logic                                   lsu_ready_i,      
    output logic                                   lsu_valid_o,      
    
    output logic                                   mult_valid_o,     
    
    input  logic                                   fpu_ready_i,      
    output logic                                   fpu_valid_o,      
    output logic [1:0]                             fpu_fmt_o,        
    output logic [2:0]                             fpu_rm_o,         
    
    output logic                                   csr_valid_o,      
    
    input  logic [NR_COMMIT_PORTS-1:0][4:0]        waddr_i,
    input  logic [NR_COMMIT_PORTS-1:0][riscv::XLEN-1:0] wdata_i,
    input  logic [NR_COMMIT_PORTS-1:0]             we_gpr_i,
    input  logic [NR_COMMIT_PORTS-1:0]             we_fpr_i
    
    
    
    
);
    logic stall;   
    logic fu_busy; 
    riscv::xlen_t    operand_a_regfile, operand_b_regfile;  
    logic [FLEN-1:0] operand_c_regfile; 
    
    riscv::xlen_t operand_a_n, operand_a_q,
                 operand_b_n, operand_b_q,
                 imm_n, imm_q;
    logic          alu_valid_q;
    logic         mult_valid_q;
    logic          fpu_valid_q;
    logic [1:0]      fpu_fmt_q;
    logic [2:0]       fpu_rm_q;
    logic          lsu_valid_q;
    logic          csr_valid_q;
    logic       branch_valid_q;
    logic [TRANS_ID_BITS-1:0] trans_id_n, trans_id_q;
    fu_op operator_n, operator_q; 
    fu_t  fu_n,       fu_q; 
    
    logic forward_rs1, forward_rs2, forward_rs3;
    
    riscv::instruction_t orig_instr;
    assign orig_instr = riscv::instruction_t'(issue_instr_i.ex.tval[31:0]);
    
    assign rs1_forwarding_o = operand_a_n[riscv::VLEN-1:0];  
    assign rs2_forwarding_o = operand_b_n[riscv::VLEN-1:0];  
    assign fu_data_o.operand_a = operand_a_q;
    assign fu_data_o.operand_b = operand_b_q;
    assign fu_data_o.fu        = fu_q;
    assign fu_data_o.operator  = operator_q;
    assign fu_data_o.trans_id  = trans_id_q;
    assign fu_data_o.imm       = imm_q;
    assign alu_valid_o         = alu_valid_q;
    assign branch_valid_o      = branch_valid_q;
    assign lsu_valid_o         = lsu_valid_q;
    assign csr_valid_o         = csr_valid_q;
    assign mult_valid_o        = mult_valid_q;
    assign fpu_valid_o         = fpu_valid_q;
    assign fpu_fmt_o           = fpu_fmt_q;
    assign fpu_rm_o            = fpu_rm_q;
    
    
    
    
    
    always_comb begin : unit_busy
        unique case (issue_instr_i.fu)
            NONE:
                fu_busy = 1'b0;
            ALU, CTRL_FLOW, CSR, MULT:
                fu_busy = ~flu_ready_i;
            FPU, FPU_VEC:
                fu_busy = ~fpu_ready_i;
            LOAD, STORE:
                fu_busy = ~lsu_ready_i;
            default:
                fu_busy = 1'b0;
        endcase
    end
    
    
    
    
    
    always_comb begin : operands_available
        stall = 1'b0;
        
        forward_rs1 = 1'b0;
        forward_rs2 = 1'b0;
        forward_rs3 = 1'b0; 
        
        rs1_o = issue_instr_i.rs1;
        rs2_o = issue_instr_i.rs2;
        rs3_o = issue_instr_i.result[REG_ADDR_SIZE-1:0]; 
        
        
        
        
        if (!issue_instr_i.use_zimm && (is_rs1_fpr(issue_instr_i.op) ? rd_clobber_fpr_i[issue_instr_i.rs1] != NONE
                                                                     : rd_clobber_gpr_i[issue_instr_i.rs1] != NONE)) begin
            
            
            
            if (rs1_valid_i && (is_rs1_fpr(issue_instr_i.op) ? 1'b1 : ((rd_clobber_gpr_i[issue_instr_i.rs1] != CSR) || (issue_instr_i.op == SFENCE_VMA)))) begin
                forward_rs1 = 1'b1;
            end else begin 
                stall = 1'b1;
            end
        end
        if (is_rs2_fpr(issue_instr_i.op) ? rd_clobber_fpr_i[issue_instr_i.rs2] != NONE
                                         : rd_clobber_gpr_i[issue_instr_i.rs2] != NONE) begin
            
            if (rs2_valid_i && (is_rs2_fpr(issue_instr_i.op) ? 1'b1 : ( (rd_clobber_gpr_i[issue_instr_i.rs2] != CSR) || (issue_instr_i.op == SFENCE_VMA))))  begin
                forward_rs2 = 1'b1;
            end else begin 
                stall = 1'b1;
            end
        end
        if (is_imm_fpr(issue_instr_i.op) && rd_clobber_fpr_i[issue_instr_i.result[REG_ADDR_SIZE-1:0]] != NONE) begin
            
            if (rs3_valid_i) begin
                forward_rs3 = 1'b1;
            end else begin 
                stall = 1'b1;
            end
        end
    end
    
    always_comb begin : forwarding_operand_select
        
        operand_a_n = operand_a_regfile;
        operand_b_n = operand_b_regfile;
        
        
        imm_n      = is_imm_fpr(issue_instr_i.op) ? {{riscv::XLEN-FLEN{1'b0}}, operand_c_regfile} : issue_instr_i.result;
        trans_id_n = issue_instr_i.trans_id;
        fu_n       = issue_instr_i.fu;
        operator_n = issue_instr_i.op;
        
        if (forward_rs1) begin
            operand_a_n  = rs1_i;
        end
        if (forward_rs2) begin
            operand_b_n  = rs2_i;
        end
        if (forward_rs3) begin
            imm_n  = {{riscv::XLEN-FLEN{1'b0}}, rs3_i};
        end
        
        if (issue_instr_i.use_pc) begin
            operand_a_n = {{riscv::XLEN-riscv::VLEN{issue_instr_i.pc[riscv::VLEN-1]}}, issue_instr_i.pc};
        end
        
        if (issue_instr_i.use_zimm) begin
            
            operand_a_n = {{riscv::XLEN-5{1'b0}}, issue_instr_i.rs1[4:0]};
        end
        
        
        if (issue_instr_i.use_imm && (issue_instr_i.fu != STORE) && (issue_instr_i.fu != CTRL_FLOW) && !is_rs2_fpr(issue_instr_i.op)) begin
            operand_b_n = issue_instr_i.result;
        end
    end
    
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        alu_valid_q    <= 1'b0;
        lsu_valid_q    <= 1'b0;
        mult_valid_q   <= 1'b0;
        fpu_valid_q    <= 1'b0;
        fpu_fmt_q      <= 2'b0;
        fpu_rm_q       <= 3'b0;
        csr_valid_q    <= 1'b0;
        branch_valid_q <= 1'b0;
      end else begin
        alu_valid_q    <= 1'b0;
        lsu_valid_q    <= 1'b0;
        mult_valid_q   <= 1'b0;
        fpu_valid_q    <= 1'b0;
        fpu_fmt_q      <= 2'b0;
        fpu_rm_q       <= 3'b0;
        csr_valid_q    <= 1'b0;
        branch_valid_q <= 1'b0;
        
        
        
        if (!issue_instr_i.ex.valid && issue_instr_valid_i && issue_ack_o) begin
            case (issue_instr_i.fu)
                ALU:
                    alu_valid_q    <= 1'b1;
                CTRL_FLOW:
                    branch_valid_q <= 1'b1;
                MULT:
                    mult_valid_q   <= 1'b1;
                FPU : begin
                    fpu_valid_q    <= 1'b1;
                    fpu_fmt_q      <= orig_instr.rftype.fmt; 
                    fpu_rm_q       <= orig_instr.rftype.rm;  
                end
                FPU_VEC : begin
                    fpu_valid_q    <= 1'b1;
                    fpu_fmt_q      <= orig_instr.rvftype.vfmt;         
                    fpu_rm_q       <= {2'b0, orig_instr.rvftype.repl}; 
                end
                LOAD, STORE:
                    lsu_valid_q    <= 1'b1;
                CSR:
                    csr_valid_q    <= 1'b1;
                default:;
            endcase
        end
        
        
        if (flush_i) begin
            alu_valid_q    <= 1'b0;
            lsu_valid_q    <= 1'b0;
            mult_valid_q   <= 1'b0;
            fpu_valid_q    <= 1'b0;
            csr_valid_q    <= 1'b0;
            branch_valid_q <= 1'b0;
        end
      end
    end
    
    
    
    always_comb begin : issue_scoreboard
        
        issue_ack_o = 1'b0;
        
        
        if (issue_instr_valid_i) begin
            
            if (!stall && !fu_busy) begin
                
                
                
                
                if (is_rd_fpr(issue_instr_i.op) ? (rd_clobber_fpr_i[issue_instr_i.rd] == NONE)
                                                : (rd_clobber_gpr_i[issue_instr_i.rd] == NONE)) begin
                    issue_ack_o = 1'b1;
                end
                
                
                for (int unsigned i = 0; i < NR_COMMIT_PORTS; i++)
                    if (is_rd_fpr(issue_instr_i.op) ? (we_fpr_i[i] && waddr_i[i] == issue_instr_i.rd)
                                                    : (we_gpr_i[i] && waddr_i[i] == issue_instr_i.rd)) begin
                        issue_ack_o = 1'b1;
                    end
            end
            
            
            
            
            
            if (issue_instr_i.ex.valid) begin
                issue_ack_o = 1'b1;
            end
            
            if (issue_instr_i.fu == NONE) begin
                issue_ack_o = 1'b1;
            end
        end
        
        
        if (mult_valid_q && issue_instr_i.fu != MULT) begin
            issue_ack_o = 1'b0;
        end
    end
    
    
    
    logic [1:0][riscv::XLEN-1:0] rdata;
    logic [1:0][4:0]  raddr_pack;
    
    logic [NR_COMMIT_PORTS-1:0][4:0]  waddr_pack;
    logic [NR_COMMIT_PORTS-1:0][riscv::XLEN-1:0] wdata_pack;
    logic [NR_COMMIT_PORTS-1:0]       we_pack;
    assign raddr_pack = {issue_instr_i.rs2[4:0], issue_instr_i.rs1[4:0]};
    for (genvar i = 0; i < NR_COMMIT_PORTS; i++) begin : gen_write_back_port
        assign waddr_pack[i] = waddr_i[i];
        assign wdata_pack[i] = wdata_i[i];
        assign we_pack[i]    = we_gpr_i[i];
    end
    ariane_regfile #(
        .DATA_WIDTH     ( riscv::XLEN     ),
        .NR_READ_PORTS  ( 2               ),
        .NR_WRITE_PORTS ( NR_COMMIT_PORTS ),
        .ZERO_REG_ZERO  ( 1               )
    ) i_ariane_regfile (
        .test_en_i ( 1'b0       ),
        .raddr_i   ( raddr_pack ),
        .rdata_o   ( rdata      ),
        .waddr_i   ( waddr_pack ),
        .wdata_i   ( wdata_pack ),
        .we_i      ( we_pack    ),
        .*
    );
    
    
    
    logic [2:0][FLEN-1:0] fprdata;
    
    logic [2:0][4:0]  fp_raddr_pack;
    logic [NR_COMMIT_PORTS-1:0][riscv::XLEN-1:0] fp_wdata_pack;
    generate
        if (FP_PRESENT) begin : float_regfile_gen
            assign fp_raddr_pack = {issue_instr_i.result[4:0], issue_instr_i.rs2[4:0], issue_instr_i.rs1[4:0]};
            for (genvar i = 0; i < NR_COMMIT_PORTS; i++) begin : gen_fp_wdata_pack
                assign fp_wdata_pack[i] = {wdata_i[i][FLEN-1:0]};
            end
            ariane_regfile #(
                .DATA_WIDTH     ( FLEN            ),
                .NR_READ_PORTS  ( 3               ),
                .NR_WRITE_PORTS ( NR_COMMIT_PORTS ),
                .ZERO_REG_ZERO  ( 0               )
            ) i_ariane_fp_regfile (
                .test_en_i ( 1'b0          ),
                .raddr_i   ( fp_raddr_pack ),
                .rdata_o   ( fprdata       ),
                .waddr_i   ( waddr_pack    ),
                .wdata_i   ( wdata_pack    ),
                .we_i      ( we_fpr_i      ),
                .*
            );
        end else begin : no_fpr_gen
            assign fprdata = '{default: '0};
        end
    endgenerate
    assign operand_a_regfile = is_rs1_fpr(issue_instr_i.op) ? {{riscv::XLEN-FLEN{1'b0}}, fprdata[0]} : rdata[0];
    assign operand_b_regfile = is_rs2_fpr(issue_instr_i.op) ? {{riscv::XLEN-FLEN{1'b0}}, fprdata[1]} : rdata[1];
    assign operand_c_regfile = fprdata[2];
    
    
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (!rst_ni) begin
            operand_a_q           <= '{default: 0};
            operand_b_q           <= '{default: 0};
            imm_q                 <= '0;
            fu_q                  <= NONE;
            operator_q            <= ADD;
            trans_id_q            <= '0;
            pc_o                  <= '0;
            is_compressed_instr_o <= 1'b0;
            branch_predict_o      <= {cf_t'(0), {riscv::VLEN{1'b0}}};
        end else begin
            operand_a_q           <= operand_a_n;
            operand_b_q           <= operand_b_n;
            imm_q                 <= imm_n;
            fu_q                  <= fu_n;
            operator_q            <= operator_n;
            trans_id_q            <= trans_id_n;
            pc_o                  <= issue_instr_i.pc;
            is_compressed_instr_o <= issue_instr_i.is_compressed;
            branch_predict_o      <= issue_instr_i.bp;
        end
    end
    
    
    
    
endmodule
module issue_stage import ariane_pkg::*; #(
    parameter int unsigned NR_ENTRIES = 8,
    parameter int unsigned NR_WB_PORTS = 4,
    parameter int unsigned NR_COMMIT_PORTS = 2
)(
    input  logic                                     clk_i,     
    input  logic                                     rst_ni,    
    output logic                                     sb_full_o,
    input  logic                                     flush_unissued_instr_i,
    input  logic                                     flush_i,
    
    input  scoreboard_entry_t                        decoded_instr_i,
    input  logic                                     decoded_instr_valid_i,
    input  logic                                     is_ctrl_flow_i,
    output logic                                     decoded_instr_ack_o,
    
    output [riscv::VLEN-1:0]                         rs1_forwarding_o,  
    output [riscv::VLEN-1:0]                         rs2_forwarding_o, 
    output fu_data_t                                 fu_data_o,
    output logic [riscv::VLEN-1:0]                   pc_o,
    output logic                                     is_compressed_instr_o,
    input  logic                                     flu_ready_i,
    output logic                                     alu_valid_o,
    
    input  logic                                     resolve_branch_i,
    input  logic                                     lsu_ready_i,
    output logic                                     lsu_valid_o,
    
    output logic                                     branch_valid_o,   
    output branchpredict_sbe_t                       branch_predict_o, 
    output logic                                     mult_valid_o,
    input  logic                                     fpu_ready_i,
    output logic                                     fpu_valid_o,
    output logic [1:0]                               fpu_fmt_o,        
    output logic [2:0]                               fpu_rm_o,         
    output logic                                     csr_valid_o,
    
    input logic [NR_WB_PORTS-1:0][TRANS_ID_BITS-1:0] trans_id_i,
    input bp_resolve_t                               resolved_branch_i,
    input logic [NR_WB_PORTS-1:0][riscv::XLEN-1:0]   wbdata_i,
    input exception_t [NR_WB_PORTS-1:0]              ex_ex_i, 
    input logic [NR_WB_PORTS-1:0]                    wt_valid_i,
    
    input  logic [NR_COMMIT_PORTS-1:0][4:0]          waddr_i,
    input  logic [NR_COMMIT_PORTS-1:0][riscv::XLEN-1:0] wdata_i,
    input  logic [NR_COMMIT_PORTS-1:0]               we_gpr_i,
    input  logic [NR_COMMIT_PORTS-1:0]               we_fpr_i,
    output scoreboard_entry_t [NR_COMMIT_PORTS-1:0]  commit_instr_o,
    input  logic              [NR_COMMIT_PORTS-1:0]  commit_ack_i
);
    
    
    
    fu_t  [2**REG_ADDR_SIZE-1:0] rd_clobber_gpr_sb_iro;
    fu_t  [2**REG_ADDR_SIZE-1:0] rd_clobber_fpr_sb_iro;
    logic [REG_ADDR_SIZE-1:0]  rs1_iro_sb;
    riscv::xlen_t              rs1_sb_iro;
    logic                      rs1_valid_sb_iro;
    logic [REG_ADDR_SIZE-1:0]  rs2_iro_sb;
    riscv::xlen_t              rs2_sb_iro;
    logic                      rs2_valid_iro_sb;
    logic [REG_ADDR_SIZE-1:0]  rs3_iro_sb;
    logic [FLEN-1:0]           rs3_sb_iro;
    logic                      rs3_valid_iro_sb;
    scoreboard_entry_t         issue_instr_rename_sb;
    logic                      issue_instr_valid_rename_sb;
    logic                      issue_ack_sb_rename;
    scoreboard_entry_t         issue_instr_sb_iro;
    logic                      issue_instr_valid_sb_iro;
    logic                      issue_ack_iro_sb;
    
    
    
    re_name i_re_name (
        .clk_i                  ( clk_i                        ),
        .rst_ni                 ( rst_ni                       ),
        .flush_i                ( flush_i                      ),
        .flush_unissied_instr_i ( flush_unissued_instr_i       ),
        .issue_instr_i          ( decoded_instr_i              ),
        .issue_instr_valid_i    ( decoded_instr_valid_i        ),
        .issue_ack_o            ( decoded_instr_ack_o          ),
        .issue_instr_o          ( issue_instr_rename_sb        ),
        .issue_instr_valid_o    ( issue_instr_valid_rename_sb  ),
        .issue_ack_i            ( issue_ack_sb_rename          )
    );
    
    
    
    scoreboard #(
        .NR_ENTRIES (NR_ENTRIES ),
        .NR_WB_PORTS(NR_WB_PORTS),
        .NR_COMMIT_PORTS(NR_COMMIT_PORTS)
    ) i_scoreboard (
        .sb_full_o             ( sb_full_o                                 ),
        .unresolved_branch_i   ( 1'b0                                      ),
        .rd_clobber_gpr_o      ( rd_clobber_gpr_sb_iro                     ),
        .rd_clobber_fpr_o      ( rd_clobber_fpr_sb_iro                     ),
        .rs1_i                 ( rs1_iro_sb                                ),
        .rs1_o                 ( rs1_sb_iro                                ),
        .rs1_valid_o           ( rs1_valid_sb_iro                          ),
        .rs2_i                 ( rs2_iro_sb                                ),
        .rs2_o                 ( rs2_sb_iro                                ),
        .rs2_valid_o           ( rs2_valid_iro_sb                          ),
        .rs3_i                 ( rs3_iro_sb                                ),
        .rs3_o                 ( rs3_sb_iro                                ),
        .rs3_valid_o           ( rs3_valid_iro_sb                          ),
        .decoded_instr_i       ( issue_instr_rename_sb                     ),
        .decoded_instr_valid_i ( issue_instr_valid_rename_sb               ),
        .decoded_instr_ack_o   ( issue_ack_sb_rename                       ),
        .issue_instr_o         ( issue_instr_sb_iro                        ),
        .issue_instr_valid_o   ( issue_instr_valid_sb_iro                  ),
        .issue_ack_i           ( issue_ack_iro_sb                          ),
        .resolved_branch_i     ( resolved_branch_i                         ),
        .trans_id_i            ( trans_id_i                                ),
        .wbdata_i              ( wbdata_i                                  ),
        .ex_i                  ( ex_ex_i                                   ),
        .*
    );
    
    
    
    issue_read_operands #(
      .NR_COMMIT_PORTS ( NR_COMMIT_PORTS )
    )i_issue_read_operands  (
        .flush_i             ( flush_unissued_instr_i          ),
        .issue_instr_i       ( issue_instr_sb_iro              ),
        .issue_instr_valid_i ( issue_instr_valid_sb_iro        ),
        .issue_ack_o         ( issue_ack_iro_sb                ),
        .fu_data_o           ( fu_data_o                       ),
        .flu_ready_i         ( flu_ready_i                     ),
        .rs1_o               ( rs1_iro_sb                      ),
        .rs1_i               ( rs1_sb_iro                      ),
        .rs1_valid_i         ( rs1_valid_sb_iro                ),
        .rs2_o               ( rs2_iro_sb                      ),
        .rs2_i               ( rs2_sb_iro                      ),
        .rs2_valid_i         ( rs2_valid_iro_sb                ),
        .rs3_o               ( rs3_iro_sb                      ),
        .rs3_i               ( rs3_sb_iro                      ),
        .rs3_valid_i         ( rs3_valid_iro_sb                ),
        .rd_clobber_gpr_i    ( rd_clobber_gpr_sb_iro           ),
        .rd_clobber_fpr_i    ( rd_clobber_fpr_sb_iro           ),
        .alu_valid_o         ( alu_valid_o                     ),
        .branch_valid_o      ( branch_valid_o                  ),
        .csr_valid_o         ( csr_valid_o                     ),
        .mult_valid_o        ( mult_valid_o                    ),
        .*
    );
endmodule
module load_unit import ariane_pkg::*; #(
    parameter ariane_pkg::ariane_cfg_t ArianeCfg = ariane_pkg::ArianeDefaultConfig
) (
    input  logic                     clk_i,    
    input  logic                     rst_ni,   
    input  logic                     flush_i,
    
    input  logic                     valid_i,
    input  lsu_ctrl_t                lsu_ctrl_i,
    output logic                     pop_ld_o,
    
    output logic                     valid_o,
    output logic [TRANS_ID_BITS-1:0] trans_id_o,
    output riscv::xlen_t             result_o,
    output exception_t               ex_o,
    
    output logic                     translation_req_o,   
    output logic [riscv::VLEN-1:0]   vaddr_o,             
    input  logic [riscv::PLEN-1:0]   paddr_i,             
    input  exception_t               ex_i,                
    input  logic                     dtlb_hit_i,          
    input  logic [riscv::PPNW-1:0]   dtlb_ppn_i,          
    
    output logic [11:0]              page_offset_o,
    input  logic                     page_offset_matches_i,
    input  logic                     store_buffer_empty_i, 
    input  logic [TRANS_ID_BITS-1:0] commit_tran_id_i,
    
    input dcache_req_o_t             req_port_i,
    output dcache_req_i_t            req_port_o,
    input  logic                     dcache_wbuffer_not_ni_i
);
    enum logic [3:0] { IDLE, WAIT_GNT, SEND_TAG, WAIT_PAGE_OFFSET,
                       ABORT_TRANSACTION, ABORT_TRANSACTION_NI, WAIT_TRANSLATION, WAIT_FLUSH,
                       WAIT_WB_EMPTY
                     } state_d, state_q;
    
    
    struct packed {
        logic [TRANS_ID_BITS-1:0] trans_id;
        logic [2:0]               address_offset;
        fu_op                     operator;
    } load_data_d, load_data_q, in_data;
    
    assign page_offset_o = lsu_ctrl_i.vaddr[11:0];
    
    assign vaddr_o = lsu_ctrl_i.vaddr;
    
    assign req_port_o.data_we = 1'b0;
    assign req_port_o.data_wdata = '0;
    
    assign in_data = {lsu_ctrl_i.trans_id, lsu_ctrl_i.vaddr[2:0], lsu_ctrl_i.operator};
    
    
    assign req_port_o.address_index = lsu_ctrl_i.vaddr[ariane_pkg::DCACHE_INDEX_WIDTH-1:0];
    
    assign req_port_o.address_tag   = paddr_i[ariane_pkg::DCACHE_TAG_WIDTH     +
                                              ariane_pkg::DCACHE_INDEX_WIDTH-1 :
                                              ariane_pkg::DCACHE_INDEX_WIDTH];
    
    assign ex_o.cause = ex_i.cause;
    assign ex_o.tval  = ex_i.tval;
    
    logic paddr_ni;
    logic not_commit_time;
    logic inflight_stores;
    logic stall_ni;
    assign paddr_ni = is_inside_nonidempotent_regions(ArianeCfg, {dtlb_ppn_i,12'd0});
    assign not_commit_time = commit_tran_id_i != lsu_ctrl_i.trans_id;
    assign inflight_stores = (!dcache_wbuffer_not_ni_i || !store_buffer_empty_i);
    assign stall_ni = (inflight_stores || not_commit_time) && paddr_ni;
    
    
    
    always_comb begin : load_control
        
        state_d              = state_q;
        load_data_d          = load_data_q;
        translation_req_o    = 1'b0;
        req_port_o.data_req  = 1'b0;
        
        req_port_o.kill_req  = 1'b0;
        req_port_o.tag_valid = 1'b0;
        req_port_o.data_be   = lsu_ctrl_i.be;
        req_port_o.data_size = extract_transfer_size(lsu_ctrl_i.operator);
        pop_ld_o             = 1'b0;
        case (state_q)
            IDLE: begin
                
                if (valid_i) begin
                    
                    
                    translation_req_o = 1'b1;
                    
                    if (!page_offset_matches_i) begin
                        
                        req_port_o.data_req = 1'b1;
                        
                        if (!req_port_i.data_gnt) begin
                            state_d = WAIT_GNT;
                        end else begin
                            if (dtlb_hit_i && !stall_ni) begin
                                
                                state_d = SEND_TAG;
                                pop_ld_o = 1'b1;
                            
                            end else if (dtlb_hit_i && stall_ni) begin
                                state_d = ABORT_TRANSACTION_NI;
                            end else begin 
                                state_d = ABORT_TRANSACTION;
                            end
                        end
                    end else begin
                        
                        state_d = WAIT_PAGE_OFFSET;
                    end
                end
            end
            
            WAIT_PAGE_OFFSET: begin
                
                if (!page_offset_matches_i) begin
                    state_d = WAIT_GNT;
                end
            end
            
            
            
            ABORT_TRANSACTION, ABORT_TRANSACTION_NI: begin
                req_port_o.kill_req  = 1'b1;
                req_port_o.tag_valid = 1'b1;
                
                state_d = (state_q == ABORT_TRANSACTION_NI) ? WAIT_WB_EMPTY :  WAIT_TRANSLATION;
            end
            
            WAIT_WB_EMPTY: begin
                
                if (dcache_wbuffer_not_ni_i) state_d = WAIT_TRANSLATION;
            end
            WAIT_TRANSLATION: begin
                translation_req_o = 1'b1;
                
                if (dtlb_hit_i)
                    state_d = WAIT_GNT;
            end
            WAIT_GNT: begin
                
                translation_req_o = 1'b1;
                
                req_port_o.data_req = 1'b1;
                
                if (req_port_i.data_gnt) begin
                    
                    if (dtlb_hit_i && !stall_ni) begin
                        state_d = SEND_TAG;
                        pop_ld_o = 1'b1;
                    
                    end else if (dtlb_hit_i && stall_ni) begin
                        state_d = ABORT_TRANSACTION_NI;
                    end else begin
                    
                        state_d = ABORT_TRANSACTION;
                    end
                end
                
            end
            
            SEND_TAG: begin
                req_port_o.tag_valid = 1'b1;
                state_d = IDLE;
                
                if (valid_i) begin
                    
                    
                    translation_req_o = 1'b1;
                    
                    if (!page_offset_matches_i) begin
                        
                        req_port_o.data_req = 1'b1;
                        
                        if (!req_port_i.data_gnt) begin
                            state_d = WAIT_GNT;
                        end else begin
                            
                            if (dtlb_hit_i && !stall_ni) begin
                                
                                state_d = SEND_TAG;
                                pop_ld_o = 1'b1;
                            
                            end else if (dtlb_hit_i && stall_ni) begin
                                state_d = ABORT_TRANSACTION_NI;
                            end else begin
                                state_d = ABORT_TRANSACTION;
                            end
                        end
                    end else begin
                        
                        state_d = WAIT_PAGE_OFFSET;
                    end
                end
                
                
                
                
                if (ex_i.valid) begin
                    req_port_o.kill_req = 1'b1;
                end
            end
            WAIT_FLUSH: begin
                
                
                req_port_o.kill_req  = 1'b1;
                req_port_o.tag_valid = 1'b1;
                
                state_d = IDLE;
            end
        endcase
        
        if (ex_i.valid && valid_i) begin
            
            state_d = IDLE;
            
            if (!req_port_i.data_rvalid)
                pop_ld_o = 1'b1;
        end
        
        if (pop_ld_o && !ex_i.valid) begin
            load_data_d = in_data;
        end
        
        if (flush_i) begin
            state_d = WAIT_FLUSH;
        end
    end
    
    
    
    
    always_comb begin : rvalid_output
        valid_o    = 1'b0;
        ex_o.valid = 1'b0;
        
        trans_id_o = load_data_q.trans_id;
        
        if (req_port_i.data_rvalid && state_q != WAIT_FLUSH) begin
            
            if(!req_port_o.kill_req)
                valid_o = 1'b1;
            
            
            
            if (ex_i.valid && (state_q == SEND_TAG)) begin
                valid_o    = 1'b1;
                ex_o.valid = 1'b1;
            end
        end
        
        
        
        
        
        if (valid_i && ex_i.valid && !req_port_i.data_rvalid) begin
            valid_o    = 1'b1;
            ex_o.valid = 1'b1;
            trans_id_o = lsu_ctrl_i.trans_id;
        
        end else if (state_q == WAIT_TRANSLATION) begin
            valid_o = 1'b0;
        end
    end
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (~rst_ni) begin
            state_q     <= IDLE;
            load_data_q <= '0;
        end else begin
            state_q     <= state_d;
            load_data_q <= load_data_d;
        end
    end
    
    
    
    logic [63:0] shifted_data;
    
    assign shifted_data   = req_port_i.data_rdata >> {load_data_q.address_offset, 3'b000};
    
    logic [7:0]  sign_bits;
    logic [2:0]  idx_d, idx_q;
    logic        sign_bit, signed_d, signed_q, fp_sign_d, fp_sign_q;
    
    assign signed_d  = load_data_d.operator  inside {ariane_pkg::LW,  ariane_pkg::LH,  ariane_pkg::LB};
    assign fp_sign_d = load_data_d.operator  inside {ariane_pkg::FLW, ariane_pkg::FLH, ariane_pkg::FLB};
    assign idx_d     = (load_data_d.operator inside {ariane_pkg::LW,  ariane_pkg::FLW}) ? load_data_d.address_offset + 3 :
                       (load_data_d.operator inside {ariane_pkg::LH,  ariane_pkg::FLH}) ? load_data_d.address_offset + 1 :
                                                                                          load_data_d.address_offset;
    assign sign_bits = { req_port_i.data_rdata[63],
                         req_port_i.data_rdata[55],
                         req_port_i.data_rdata[47],
                         req_port_i.data_rdata[39],
                         req_port_i.data_rdata[31],
                         req_port_i.data_rdata[23],
                         req_port_i.data_rdata[15],
                         req_port_i.data_rdata[7]  };
    
    
    assign sign_bit       = signed_q & sign_bits[idx_q] | fp_sign_q;
    
    always_comb begin
        unique case (load_data_q.operator)
            ariane_pkg::LW, ariane_pkg::LWU, ariane_pkg::FLW:    result_o = {{riscv::XLEN-32{sign_bit}}, shifted_data[31:0]};
            ariane_pkg::LH, ariane_pkg::LHU, ariane_pkg::FLH:    result_o = {{riscv::XLEN-32+16{sign_bit}}, shifted_data[15:0]};
            ariane_pkg::LB, ariane_pkg::LBU, ariane_pkg::FLB:    result_o = {{riscv::XLEN-32+24{sign_bit}}, shifted_data[7:0]};
            default:    result_o = shifted_data[riscv::XLEN-1:0];
        endcase
    end
    always_ff @(posedge clk_i or negedge rst_ni) begin : p_regs
        if (~rst_ni) begin
            idx_q     <= 0;
            signed_q  <= 0;
            fp_sign_q <= 0;
        end else begin
            idx_q     <= idx_d;
            signed_q  <= signed_d;
            fp_sign_q <= fp_sign_d;
        end
    end
    
endmodule
module load_store_unit import ariane_pkg::*; #(
    parameter int unsigned ASID_WIDTH = 1,
    parameter ariane_pkg::ariane_cfg_t ArianeCfg = ariane_pkg::ArianeDefaultConfig
)(
    input  logic                     clk_i,
    input  logic                     rst_ni,
    input  logic                     flush_i,
    output logic                     no_st_pending_o,
    input  logic                     amo_valid_commit_i,
    input  fu_data_t                 fu_data_i,
    output logic                     lsu_ready_o,              
    input  logic                     lsu_valid_i,              
    output logic [TRANS_ID_BITS-1:0] load_trans_id_o,          
    output riscv::xlen_t             load_result_o,
    output logic                     load_valid_o,
    output exception_t               load_exception_o,         
    output logic [TRANS_ID_BITS-1:0] store_trans_id_o,         
    output riscv::xlen_t             store_result_o,
    output logic                     store_valid_o,
    output exception_t               store_exception_o,        
    input  logic                     commit_i,                 
    output logic                     commit_ready_o,           
    input  logic [TRANS_ID_BITS-1:0] commit_tran_id_i,
    input  logic                     enable_translation_i,     
    input  logic                     en_ld_st_translation_i,   
    
    input  icache_areq_o_t           icache_areq_i,
    output icache_areq_i_t           icache_areq_o,
    input  riscv::priv_lvl_t         priv_lvl_i,               
    input  riscv::priv_lvl_t         ld_st_priv_lvl_i,         
    input  logic                     sum_i,                    
    input  logic                     mxr_i,                    
    input  logic [riscv::PPNW-1:0]   satp_ppn_i,               
    input  logic [ASID_WIDTH-1:0]    asid_i,                   
    input  logic [ASID_WIDTH-1:0]    asid_to_be_flushed_i,
    input  logic [riscv::VLEN-1:0]   vaddr_to_be_flushed_i,
    input  logic                     flush_tlb_i,
    
    output logic                     itlb_miss_o,
    output logic                     dtlb_miss_o,
    
    input  dcache_req_o_t [2:0]      dcache_req_ports_i,
    output dcache_req_i_t [2:0]      dcache_req_ports_o,
    input  logic                     dcache_wbuffer_empty_i,
    input  logic                     dcache_wbuffer_not_ni_i,
    
    output amo_req_t                 amo_req_o,
    input  amo_resp_t                amo_resp_i,
    
    input  riscv::pmpcfg_t [15:0]    pmpcfg_i,
    input  logic [15:0][riscv::PLEN-3:0] pmpaddr_i
);
    
    logic data_misaligned;
    
    
    
    
    
    lsu_ctrl_t lsu_ctrl;
    logic      pop_st;
    logic      pop_ld;
    
    
    
    
    logic [riscv::VLEN-1:0]   vaddr_i;
    riscv::xlen_t             vaddr_xlen;
    logic                     overflow;
    logic [7:0]               be_i;
    assign vaddr_xlen = $unsigned($signed(fu_data_i.imm) + $signed(fu_data_i.operand_a));
    assign vaddr_i = vaddr_xlen[riscv::VLEN-1:0];
    
    assign overflow = !((&vaddr_xlen[riscv::XLEN-1:riscv::SV-1]) == 1'b1 || (|vaddr_xlen[riscv::XLEN-1:riscv::SV-1]) == 1'b0);
    logic                     st_valid_i;
    logic                     ld_valid_i;
    logic                     ld_translation_req;
    logic                     st_translation_req;
    logic [riscv::VLEN-1:0]   ld_vaddr;
    logic [riscv::VLEN-1:0]   st_vaddr;
    logic                     translation_req;
    logic                     translation_valid;
    logic [riscv::VLEN-1:0]   mmu_vaddr;
    logic [riscv::PLEN-1:0]   mmu_paddr;
    exception_t               mmu_exception;
    logic                     dtlb_hit;
    logic [riscv::PPNW-1:0]   dtlb_ppn;
    logic                     ld_valid;
    logic [TRANS_ID_BITS-1:0] ld_trans_id;
    riscv::xlen_t             ld_result;
    logic                     st_valid;
    logic [TRANS_ID_BITS-1:0] st_trans_id;
    riscv::xlen_t             st_result;
    logic [11:0]              page_offset;
    logic                     page_offset_matches;
    exception_t               misaligned_exception;
    exception_t               ld_ex;
    exception_t               st_ex;
    
    
    
    if (MMU_PRESENT && (riscv::XLEN == 64)) begin : gen_mmu_sv39
        mmu #(
            .INSTR_TLB_ENTRIES      ( 16                     ),
            .DATA_TLB_ENTRIES       ( 16                     ),
            .ASID_WIDTH             ( ASID_WIDTH             ),
            .ArianeCfg              ( ArianeCfg              )
        ) i_cva6_mmu (
            
            .misaligned_ex_i        ( misaligned_exception   ),
            .lsu_is_store_i         ( st_translation_req     ),
            .lsu_req_i              ( translation_req        ),
            .lsu_vaddr_i            ( mmu_vaddr              ),
            .lsu_valid_o            ( translation_valid      ),
            .lsu_paddr_o            ( mmu_paddr              ),
            .lsu_exception_o        ( mmu_exception          ),
            .lsu_dtlb_hit_o         ( dtlb_hit               ), 
            .lsu_dtlb_ppn_o         ( dtlb_ppn               ), 
            
            .req_port_i             ( dcache_req_ports_i [0] ),
            .req_port_o             ( dcache_req_ports_o [0] ),
            
            .icache_areq_i          ( icache_areq_i          ),
            .asid_to_be_flushed_i,
            .vaddr_to_be_flushed_i,
            .icache_areq_o          ( icache_areq_o          ),
            .pmpcfg_i,
            .pmpaddr_i,
            .*
        );
    end else if (MMU_PRESENT && (riscv::XLEN == 32)) begin : gen_mmu_sv32
        cva6_mmu_sv32 #(
            .INSTR_TLB_ENTRIES      ( 16                     ),
            .DATA_TLB_ENTRIES       ( 16                     ),
            .ASID_WIDTH             ( ASID_WIDTH             ),
            .ArianeCfg              ( ArianeCfg              )
        ) i_cva6_mmu (
            
            .misaligned_ex_i        ( misaligned_exception   ),
            .lsu_is_store_i         ( st_translation_req     ),
            .lsu_req_i              ( translation_req        ),
            .lsu_vaddr_i            ( mmu_vaddr              ),
            .lsu_valid_o            ( translation_valid      ),
            .lsu_paddr_o            ( mmu_paddr              ),
            .lsu_exception_o        ( mmu_exception          ),
            .lsu_dtlb_hit_o         ( dtlb_hit               ), 
            .lsu_dtlb_ppn_o         ( dtlb_ppn               ), 
            
            .req_port_i             ( dcache_req_ports_i [0] ),
            .req_port_o             ( dcache_req_ports_o [0] ),
            
            .icache_areq_i          ( icache_areq_i          ),
            .asid_to_be_flushed_i,
            .vaddr_to_be_flushed_i,
            .icache_areq_o          ( icache_areq_o          ),
            .pmpcfg_i,
            .pmpaddr_i,
            .*
        );
    end else begin : gen_no_mmu
        assign  icache_areq_o.fetch_valid  = icache_areq_i.fetch_req;
        assign  icache_areq_o.fetch_paddr  = icache_areq_i.fetch_vaddr[riscv::PLEN-1:0];
        assign  icache_areq_o.fetch_exception      = '0;
        assign dcache_req_ports_o[0].address_index = '0;
        assign dcache_req_ports_o[0].address_tag   = '0;
        assign dcache_req_ports_o[0].data_wdata    = 64'b0;
        assign dcache_req_ports_o[0].data_req      = 1'b0;
        assign dcache_req_ports_o[0].data_be       = 8'hFF;
        assign dcache_req_ports_o[0].data_size     = 2'b11;
        assign dcache_req_ports_o[0].data_we       = 1'b0;
        assign dcache_req_ports_o[0].kill_req      = '0;
        assign dcache_req_ports_o[0].tag_valid     = 1'b0;
        assign itlb_miss_o = 1'b0;
        assign dtlb_miss_o = 1'b0;
        assign dtlb_ppn    = mmu_vaddr[riscv::PLEN-1:12];
        assign dtlb_hit    = 1'b1;
        assign mmu_exception = '0;
        always_ff @(posedge clk_i or negedge rst_ni) begin
            if (~rst_ni) begin
                mmu_paddr         <= '0;
                translation_valid <= '0;
            end else begin
                mmu_paddr         <=  mmu_vaddr[riscv::PLEN-1:0];
                translation_valid <= translation_req;
            end
        end
    end
    logic store_buffer_empty;
    
    
    
    store_unit i_store_unit (
        .clk_i,
        .rst_ni,
        .flush_i,
        .no_st_pending_o,
        .store_buffer_empty_o  ( store_buffer_empty   ),
        .valid_i               ( st_valid_i           ),
        .lsu_ctrl_i            ( lsu_ctrl             ),
        .pop_st_o              ( pop_st               ),
        .commit_i,
        .commit_ready_o,
        .amo_valid_commit_i,
        .valid_o               ( st_valid             ),
        .trans_id_o            ( st_trans_id          ),
        .result_o              ( st_result            ),
        .ex_o                  ( st_ex                ),
        
        .translation_req_o     ( st_translation_req   ),
        .vaddr_o               ( st_vaddr             ),
        .paddr_i               ( mmu_paddr            ),
        .ex_i                  ( mmu_exception        ),
        .dtlb_hit_i            ( dtlb_hit             ),
        
        .page_offset_i         ( page_offset          ),
        .page_offset_matches_o ( page_offset_matches  ),
        
        .amo_req_o,
        .amo_resp_i,
        
        .req_port_i             ( dcache_req_ports_i [2] ),
        .req_port_o             ( dcache_req_ports_o [2] )
    );
    
    
    
    load_unit #(
        .ArianeCfg ( ArianeCfg )
    ) i_load_unit (
        .valid_i               ( ld_valid_i           ),
        .lsu_ctrl_i            ( lsu_ctrl             ),
        .pop_ld_o              ( pop_ld               ),
        .valid_o               ( ld_valid             ),
        .trans_id_o            ( ld_trans_id          ),
        .result_o              ( ld_result            ),
        .ex_o                  ( ld_ex                ),
        
        .translation_req_o     ( ld_translation_req   ),
        .vaddr_o               ( ld_vaddr             ),
        .paddr_i               ( mmu_paddr            ),
        .ex_i                  ( mmu_exception        ),
        .dtlb_hit_i            ( dtlb_hit             ),
        .dtlb_ppn_i            ( dtlb_ppn             ),
        
        .page_offset_o         ( page_offset          ),
        .page_offset_matches_i ( page_offset_matches  ),
        .store_buffer_empty_i  ( store_buffer_empty   ),
        
        .req_port_i            ( dcache_req_ports_i [1] ),
        .req_port_o            ( dcache_req_ports_o [1] ),
        .dcache_wbuffer_not_ni_i,
        .commit_tran_id_i,
        .*
    );
    
    
    
    shift_reg #(
        .dtype ( logic[$bits(ld_valid) + $bits(ld_trans_id) + $bits(ld_result) + $bits(ld_ex) - 1: 0]),
        .Depth ( NR_LOAD_PIPE_REGS )
    ) i_pipe_reg_load (
        .clk_i,
        .rst_ni,
        .d_i ( {ld_valid, ld_trans_id, ld_result, ld_ex} ),
        .d_o ( {load_valid_o, load_trans_id_o, load_result_o, load_exception_o} )
    );
    shift_reg #(
        .dtype ( logic[$bits(st_valid) + $bits(st_trans_id) + $bits(st_result) + $bits(st_ex) - 1: 0]),
        .Depth ( NR_STORE_PIPE_REGS )
    ) i_pipe_reg_store (
        .clk_i,
        .rst_ni,
        .d_i ( {st_valid, st_trans_id, st_result, st_ex} ),
        .d_o ( {store_valid_o, store_trans_id_o, store_result_o, store_exception_o} )
    );
    
    always_comb begin : which_op
        ld_valid_i = 1'b0;
        st_valid_i = 1'b0;
        translation_req      = 1'b0;
        mmu_vaddr            = {riscv::VLEN{1'b0}};
        
        unique case (lsu_ctrl.fu)
            
            LOAD:  begin
                ld_valid_i           = lsu_ctrl.valid;
                translation_req      = ld_translation_req;
                mmu_vaddr            = ld_vaddr;
            end
            
            STORE: begin
                st_valid_i           = lsu_ctrl.valid;
                translation_req      = st_translation_req;
                mmu_vaddr            = st_vaddr;
            end
            
            default: ;
        endcase
    end
    
    
    
    
    
    
    assign be_i = be_gen(vaddr_i[2:0], extract_transfer_size(fu_data_i.operator));
    
    
    
    
    
    
    always_comb begin : data_misaligned_detection
        misaligned_exception = {
            {riscv::XLEN{1'b0}},
            {riscv::XLEN{1'b0}},
            1'b0
        };
        data_misaligned = 1'b0;
        if (lsu_ctrl.valid) begin
            case (lsu_ctrl.operator)
                
                LD, SD, FLD, FSD,
                AMO_LRD, AMO_SCD,
                AMO_SWAPD, AMO_ADDD, AMO_ANDD, AMO_ORD,
                AMO_XORD, AMO_MAXD, AMO_MAXDU, AMO_MIND,
                AMO_MINDU: begin
                    if (lsu_ctrl.vaddr[2:0] != 3'b000) begin
                        data_misaligned = 1'b1;
                    end
                end
                
                LW, LWU, SW, FLW, FSW,
                AMO_LRW, AMO_SCW,
                AMO_SWAPW, AMO_ADDW, AMO_ANDW, AMO_ORW,
                AMO_XORW, AMO_MAXW, AMO_MAXWU, AMO_MINW,
                AMO_MINWU: begin
                    if (lsu_ctrl.vaddr[1:0] != 2'b00) begin
                        data_misaligned = 1'b1;
                    end
                end
                
                LH, LHU, SH, FLH, FSH: begin
                    if (lsu_ctrl.vaddr[0] != 1'b0) begin
                        data_misaligned = 1'b1;
                    end
                end
                
                default:;
            endcase
        end
        if (data_misaligned) begin
            if (lsu_ctrl.fu == LOAD) begin
                misaligned_exception = {
                    riscv::LD_ADDR_MISALIGNED,
                    {{riscv::XLEN-riscv::VLEN{1'b0}},lsu_ctrl.vaddr},
                    1'b1
                };
            end else if (lsu_ctrl.fu == STORE) begin
                misaligned_exception = {
                    riscv::ST_ADDR_MISALIGNED,
                    {{riscv::XLEN-riscv::VLEN{1'b0}},lsu_ctrl.vaddr},
                    1'b1
                };
            end
        end
        if (en_ld_st_translation_i && lsu_ctrl.overflow) begin
            if (lsu_ctrl.fu == LOAD) begin
                misaligned_exception = {
                    riscv::LD_ACCESS_FAULT,
                    {{riscv::XLEN-riscv::VLEN{1'b0}},lsu_ctrl.vaddr},
                    1'b1
                };
            end else if (lsu_ctrl.fu == STORE) begin
                misaligned_exception = {
                    riscv::ST_ACCESS_FAULT,
                    {{riscv::XLEN-riscv::VLEN{1'b0}},lsu_ctrl.vaddr},
                    1'b1
                };
            end
        end
    end
    
    
    
    
    lsu_ctrl_t lsu_req_i;
    assign lsu_req_i = {lsu_valid_i, vaddr_i, overflow, {{64-riscv::XLEN{1'b0}}, fu_data_i.operand_b}, be_i, fu_data_i.fu, fu_data_i.operator, fu_data_i.trans_id};
    lsu_bypass lsu_bypass_i (
        .lsu_req_i          ( lsu_req_i   ),
        .lsu_req_valid_i    ( lsu_valid_i ),
        .pop_ld_i           ( pop_ld      ),
        .pop_st_i           ( pop_st      ),
        .lsu_ctrl_o         ( lsu_ctrl    ),
        .ready_o            ( lsu_ready_o ),
        .*
    );
endmodule
module lsu_bypass import ariane_pkg::*; (
    input  logic      clk_i,
    input  logic      rst_ni,
    input  logic      flush_i,
    input  lsu_ctrl_t lsu_req_i,
    input  logic      lsu_req_valid_i,
    input  logic      pop_ld_i,
    input  logic      pop_st_i,
    output lsu_ctrl_t lsu_ctrl_o,
    output logic      ready_o
    );
    lsu_ctrl_t [1:0] mem_n, mem_q;
    logic read_pointer_n, read_pointer_q;
    logic write_pointer_n, write_pointer_q;
    logic [1:0] status_cnt_n, status_cnt_q;
    logic  empty;
    assign empty = (status_cnt_q == 0);
    assign ready_o = empty;
    always_comb begin
        automatic logic [1:0] status_cnt;
        automatic logic write_pointer;
        automatic logic read_pointer;
        status_cnt = status_cnt_q;
        write_pointer = write_pointer_q;
        read_pointer = read_pointer_q;
        mem_n = mem_q;
        
        if (lsu_req_valid_i) begin
            mem_n[write_pointer_q] = lsu_req_i;
            write_pointer++;
            status_cnt++;
        end
        if (pop_ld_i) begin
            
            mem_n[read_pointer_q].valid = 1'b0;
            read_pointer++;
            status_cnt--;
        end
        if (pop_st_i) begin
            
            mem_n[read_pointer_q].valid = 1'b0;
            read_pointer++;
            status_cnt--;
        end
        if (pop_st_i && pop_ld_i)
            mem_n = '0;
        if (flush_i) begin
            status_cnt = '0;
            write_pointer = '0;
            read_pointer = '0;
            mem_n = '0;
        end
        
        read_pointer_n  = read_pointer;
        write_pointer_n = write_pointer;
        status_cnt_n    = status_cnt;
    end
    
    always_comb begin : output_assignments
        if (empty) begin
            lsu_ctrl_o = lsu_req_i;
        end else begin
            lsu_ctrl_o = mem_q[read_pointer_q];
        end
    end
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (~rst_ni) begin
            mem_q           <= '0;
            status_cnt_q    <= '0;
            write_pointer_q <= '0;
            read_pointer_q  <= '0;
        end else begin
            mem_q           <= mem_n;
            status_cnt_q    <= status_cnt_n;
            write_pointer_q <= write_pointer_n;
            read_pointer_q  <= read_pointer_n;
        end
    end
endmodule
module mmu import ariane_pkg::*; #(
    parameter int unsigned INSTR_TLB_ENTRIES     = 4,
    parameter int unsigned DATA_TLB_ENTRIES      = 4,
    parameter int unsigned ASID_WIDTH            = 1,
    parameter ariane_pkg::ariane_cfg_t ArianeCfg = ariane_pkg::ArianeDefaultConfig
) (
    input  logic                            clk_i,
    input  logic                            rst_ni,
    input  logic                            flush_i,
    input  logic                            enable_translation_i,
    input  logic                            en_ld_st_translation_i,   
    
    input  icache_areq_o_t                  icache_areq_i,
    output icache_areq_i_t                  icache_areq_o,
    
    
    
    input  exception_t                      misaligned_ex_i,
    input  logic                            lsu_req_i,        
    input  logic [riscv::VLEN-1:0]          lsu_vaddr_i,      
    input  logic                            lsu_is_store_i,   
    
    
    output logic                            lsu_dtlb_hit_o,   
    output logic [riscv::PPNW-1:0]          lsu_dtlb_ppn_o,   
    
    output logic                            lsu_valid_o,      
    output logic [riscv::PLEN-1:0]          lsu_paddr_o,      
    output exception_t                      lsu_exception_o,  
    
    input riscv::priv_lvl_t                 priv_lvl_i,
    input riscv::priv_lvl_t                 ld_st_priv_lvl_i,
    input logic                             sum_i,
    input logic                             mxr_i,
    
    input logic [riscv::PPNW-1:0]           satp_ppn_i,
    input logic [ASID_WIDTH-1:0]            asid_i,
    input logic [ASID_WIDTH-1:0]            asid_to_be_flushed_i,
    input logic [riscv::VLEN-1:0]           vaddr_to_be_flushed_i,
    input logic                             flush_tlb_i,
    
    output logic                            itlb_miss_o,
    output logic                            dtlb_miss_o,
    
    input  dcache_req_o_t                   req_port_i,
    output dcache_req_i_t                   req_port_o,
    
    input  riscv::pmpcfg_t [15:0]           pmpcfg_i,
    input  logic [15:0][riscv::PLEN-3:0]    pmpaddr_i
);
    logic                   iaccess_err;   
    logic                   daccess_err;   
    logic                   ptw_active;    
    logic                   walking_instr; 
    logic                   ptw_error;     
    logic                   ptw_access_exception; 
    logic [riscv::PLEN-1:0] ptw_bad_paddr; 
    logic [riscv::VLEN-1:0] update_vaddr;
    tlb_update_t update_ptw_itlb, update_ptw_dtlb;
    logic        itlb_lu_access;
    riscv::pte_t itlb_content;
    logic        itlb_is_2M;
    logic        itlb_is_1G;
    logic        itlb_lu_hit;
    logic        dtlb_lu_access;
    riscv::pte_t dtlb_content;
    logic        dtlb_is_2M;
    logic        dtlb_is_1G;
    logic        dtlb_lu_hit;
    
    assign itlb_lu_access = icache_areq_i.fetch_req;
    assign dtlb_lu_access = lsu_req_i;
    tlb #(
        .TLB_ENTRIES      ( INSTR_TLB_ENTRIES          ),
        .ASID_WIDTH       ( ASID_WIDTH                 )
    ) i_itlb (
        .clk_i            ( clk_i                      ),
        .rst_ni           ( rst_ni                     ),
        .flush_i          ( flush_tlb_i                ),
        .update_i         ( update_ptw_itlb            ),
        .lu_access_i      ( itlb_lu_access             ),
        .lu_asid_i        ( asid_i                     ),
        .asid_to_be_flushed_i  ( asid_to_be_flushed_i  ),
        .vaddr_to_be_flushed_i ( vaddr_to_be_flushed_i ),
        .lu_vaddr_i       ( icache_areq_i.fetch_vaddr  ),
        .lu_content_o     ( itlb_content               ),
        .lu_is_2M_o       ( itlb_is_2M                 ),
        .lu_is_1G_o       ( itlb_is_1G                 ),
        .lu_hit_o         ( itlb_lu_hit                )
    );
    tlb #(
        .TLB_ENTRIES     ( DATA_TLB_ENTRIES             ),
        .ASID_WIDTH      ( ASID_WIDTH                   )
    ) i_dtlb (
        .clk_i            ( clk_i                       ),
        .rst_ni           ( rst_ni                      ),
        .flush_i          ( flush_tlb_i                 ),
        .update_i         ( update_ptw_dtlb             ),
        .lu_access_i      ( dtlb_lu_access              ),
        .lu_asid_i        ( asid_i                      ),
	      .asid_to_be_flushed_i  ( asid_to_be_flushed_i   ),
	      .vaddr_to_be_flushed_i ( vaddr_to_be_flushed_i  ),
        .lu_vaddr_i       ( lsu_vaddr_i                 ),
        .lu_content_o     ( dtlb_content                ),
        .lu_is_2M_o       ( dtlb_is_2M                  ),
        .lu_is_1G_o       ( dtlb_is_1G                  ),
        .lu_hit_o         ( dtlb_lu_hit                 )
    );
    ptw  #(
        .ASID_WIDTH             ( ASID_WIDTH            ),
        .ArianeCfg              ( ArianeCfg             )
    ) i_ptw (
        .clk_i                  ( clk_i                 ),
        .rst_ni                 ( rst_ni                ),
        .ptw_active_o           ( ptw_active            ),
        .walking_instr_o        ( walking_instr         ),
        .ptw_error_o            ( ptw_error             ),
        .ptw_access_exception_o ( ptw_access_exception  ),
        .enable_translation_i   ( enable_translation_i  ),
        .update_vaddr_o         ( update_vaddr          ),
        .itlb_update_o          ( update_ptw_itlb       ),
        .dtlb_update_o          ( update_ptw_dtlb       ),
        .itlb_access_i          ( itlb_lu_access        ),
        .itlb_hit_i             ( itlb_lu_hit           ),
        .itlb_vaddr_i           ( icache_areq_i.fetch_vaddr ),
        .dtlb_access_i          ( dtlb_lu_access        ),
        .dtlb_hit_i             ( dtlb_lu_hit           ),
        .dtlb_vaddr_i           ( lsu_vaddr_i           ),
        .req_port_i             ( req_port_i            ),
        .req_port_o             ( req_port_o            ),
        .pmpcfg_i,
        .pmpaddr_i,
        .bad_paddr_o            ( ptw_bad_paddr         ),
        .*
    );
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    logic match_any_execute_region;
    logic pmp_instr_allow;
    
    always_comb begin : instr_interface
        
        icache_areq_o.fetch_valid  = icache_areq_i.fetch_req;
        icache_areq_o.fetch_paddr  = icache_areq_i.fetch_vaddr[riscv::PLEN-1:0]; 
        
        
        
        icache_areq_o.fetch_exception      = '0;
        
        iaccess_err   = icache_areq_i.fetch_req && (((priv_lvl_i == riscv::PRIV_LVL_U) && ~itlb_content.u)
                                                 || ((priv_lvl_i == riscv::PRIV_LVL_S) && itlb_content.u));
        
        
        
        
        if (enable_translation_i) begin
            
            if (icache_areq_i.fetch_req && !((&icache_areq_i.fetch_vaddr[riscv::VLEN-1:riscv::SV-1]) == 1'b1 || (|icache_areq_i.fetch_vaddr[riscv::VLEN-1:riscv::SV-1]) == 1'b0)) begin
                icache_areq_o.fetch_exception = {riscv::INSTR_ACCESS_FAULT, {{riscv::XLEN-riscv::VLEN{1'b0}}, icache_areq_i.fetch_vaddr}, 1'b1};
            end
            icache_areq_o.fetch_valid = 1'b0;
            
            icache_areq_o.fetch_paddr = {itlb_content.ppn, icache_areq_i.fetch_vaddr[11:0]};
            
            if (itlb_is_2M) begin
                icache_areq_o.fetch_paddr[20:12] = icache_areq_i.fetch_vaddr[20:12];
            end
            
            if (itlb_is_1G) begin
                icache_areq_o.fetch_paddr[29:12] = icache_areq_i.fetch_vaddr[29:12];
            end
            
            
            
            
            if (itlb_lu_hit) begin
                icache_areq_o.fetch_valid = icache_areq_i.fetch_req;
                
                if (iaccess_err) begin
                    
                    icache_areq_o.fetch_exception = {riscv::INSTR_PAGE_FAULT, {{riscv::XLEN-riscv::VLEN{1'b0}}, icache_areq_i.fetch_vaddr}, 1'b1};
                end else if (!pmp_instr_allow) begin
                    icache_areq_o.fetch_exception = {riscv::INSTR_ACCESS_FAULT, {{riscv::XLEN-riscv::PLEN{1'b0}}, icache_areq_i.fetch_vaddr}, 1'b1};
                end
            end else
            
            
            
            
            if (ptw_active && walking_instr) begin
                icache_areq_o.fetch_valid = ptw_error | ptw_access_exception;
                if (ptw_error) icache_areq_o.fetch_exception = {riscv::INSTR_PAGE_FAULT, {{riscv::XLEN-riscv::VLEN{1'b0}}, update_vaddr}, 1'b1};
                
                else icache_areq_o.fetch_exception = {riscv::INSTR_ACCESS_FAULT, {{riscv::XLEN-riscv::VLEN{1'b0}}, ptw_bad_paddr}, 1'b1};
            end
        end
        
        
        if (!match_any_execute_region || (!enable_translation_i && !pmp_instr_allow)) begin
          icache_areq_o.fetch_exception = {riscv::INSTR_ACCESS_FAULT, {{riscv::XLEN-riscv::PLEN{1'b0}}, icache_areq_o.fetch_paddr}, 1'b1};
        end
    end
    
    assign match_any_execute_region = ariane_pkg::is_inside_execute_regions(ArianeCfg, {{64-riscv::PLEN{1'b0}}, icache_areq_o.fetch_paddr});
    
    pmp #(
        .PLEN       ( riscv::PLEN            ),
        .PMP_LEN    ( riscv::PLEN - 2        ),
        .NR_ENTRIES ( ArianeCfg.NrPMPEntries )
    ) i_pmp_if (
        .addr_i        ( icache_areq_o.fetch_paddr ),
        .priv_lvl_i,
        
        .access_type_i ( riscv::ACCESS_EXEC        ),
        
        .conf_addr_i   ( pmpaddr_i                 ),
        .conf_i        ( pmpcfg_i                  ),
        .allow_o       ( pmp_instr_allow           )
    );
    
    
    
    logic [riscv::VLEN-1:0] lsu_vaddr_n,     lsu_vaddr_q;
    riscv::pte_t dtlb_pte_n,      dtlb_pte_q;
    exception_t  misaligned_ex_n, misaligned_ex_q;
    logic        lsu_req_n,       lsu_req_q;
    logic        lsu_is_store_n,  lsu_is_store_q;
    logic        dtlb_hit_n,      dtlb_hit_q;
    logic        dtlb_is_2M_n,    dtlb_is_2M_q;
    logic        dtlb_is_1G_n,    dtlb_is_1G_q;
    
    assign lsu_dtlb_hit_o = (en_ld_st_translation_i) ? dtlb_lu_hit :  1'b1;
    
    riscv::pmp_access_t pmp_access_type;
    logic        pmp_data_allow;
    localparam   PPNWMin = (riscv::PPNW-1 > 29) ? 29 : riscv::PPNW-1;
    
    always_comb begin : data_interface
        
        lsu_vaddr_n           = lsu_vaddr_i;
        lsu_req_n             = lsu_req_i;
        misaligned_ex_n       = misaligned_ex_i;
        dtlb_pte_n            = dtlb_content;
        dtlb_hit_n            = dtlb_lu_hit;
        lsu_is_store_n        = lsu_is_store_i;
        dtlb_is_2M_n          = dtlb_is_2M;
        dtlb_is_1G_n          = dtlb_is_1G;
        lsu_paddr_o           = lsu_vaddr_q[riscv::PLEN-1:0];
        lsu_dtlb_ppn_o        = lsu_vaddr_n[riscv::PLEN-1:12];
        lsu_valid_o           = lsu_req_q;
        lsu_exception_o       = misaligned_ex_q;
        pmp_access_type       = lsu_is_store_q ? riscv::ACCESS_WRITE : riscv::ACCESS_READ;
        
        misaligned_ex_n.valid = misaligned_ex_i.valid & lsu_req_i;
        
        
        daccess_err = (ld_st_priv_lvl_i == riscv::PRIV_LVL_S && !sum_i && dtlb_pte_q.u) || 
                      (ld_st_priv_lvl_i == riscv::PRIV_LVL_U && !dtlb_pte_q.u);            
        
        if (en_ld_st_translation_i && !misaligned_ex_q.valid) begin
            lsu_valid_o = 1'b0;
            
            lsu_paddr_o = {dtlb_pte_q.ppn, lsu_vaddr_q[11:0]};
            lsu_dtlb_ppn_o = dtlb_content.ppn;
            
            if (dtlb_is_2M_q) begin
              lsu_paddr_o[20:12] = lsu_vaddr_q[20:12];
              lsu_dtlb_ppn_o[20:12] = lsu_vaddr_n[20:12];
            end
            
            if (dtlb_is_1G_q) begin
                lsu_paddr_o[PPNWMin:12] = lsu_vaddr_q[PPNWMin:12];
                lsu_dtlb_ppn_o[PPNWMin:12] = lsu_vaddr_n[PPNWMin:12];
            end
            
            
            
            if (dtlb_hit_q && lsu_req_q) begin
                lsu_valid_o = 1'b1;
                
                
                
                
                
                if (lsu_is_store_q) begin
                    
                    
                    if (!dtlb_pte_q.w || daccess_err || !dtlb_pte_q.d) begin
                        lsu_exception_o = {riscv::STORE_PAGE_FAULT, {{riscv::XLEN-riscv::VLEN{lsu_vaddr_q[riscv::VLEN-1]}},lsu_vaddr_q}, 1'b1};
                    
                    end else if (!pmp_data_allow) begin
                        lsu_exception_o = {riscv::ST_ACCESS_FAULT, {{riscv::XLEN-riscv::PLEN{1'b0}}, lsu_paddr_o}, 1'b1};
                    end
                
                end else begin
                    
                    if (daccess_err) begin
                        lsu_exception_o = {riscv::LOAD_PAGE_FAULT, {{riscv::XLEN-riscv::VLEN{lsu_vaddr_q[riscv::VLEN-1]}},lsu_vaddr_q}, 1'b1};
                    
                    end else if (!pmp_data_allow) begin
                        lsu_exception_o = {riscv::LD_ACCESS_FAULT, {{riscv::XLEN-riscv::PLEN{1'b0}}, lsu_paddr_o}, 1'b1};
                    end
                end
            end else
            
            
            
            
            if (ptw_active && !walking_instr) begin
                
                if (ptw_error) begin
                    
                    lsu_valid_o = 1'b1;
                    
                    if (lsu_is_store_q) begin
                        lsu_exception_o = {riscv::STORE_PAGE_FAULT, {{riscv::XLEN-riscv::VLEN{lsu_vaddr_q[riscv::VLEN-1]}},update_vaddr}, 1'b1};
                    end else begin
                        lsu_exception_o = {riscv::LOAD_PAGE_FAULT, {{riscv::XLEN-riscv::VLEN{lsu_vaddr_q[riscv::VLEN-1]}},update_vaddr}, 1'b1};
                    end
                end
                if (ptw_access_exception) begin
                    
                    lsu_valid_o = 1'b1;
                    
                    lsu_exception_o = {riscv::LD_ACCESS_FAULT, {{riscv::XLEN-riscv::PLEN{1'b0}}, ptw_bad_paddr}, 1'b1};
                end
            end
        end
        
        else if (lsu_req_q && !misaligned_ex_q.valid && !pmp_data_allow) begin
            if (lsu_is_store_q) begin
                lsu_exception_o = {riscv::ST_ACCESS_FAULT, {{riscv::XLEN-riscv::PLEN{1'b0}}, lsu_paddr_o}, 1'b1};
            end else begin
                lsu_exception_o = {riscv::LD_ACCESS_FAULT, {{riscv::XLEN-riscv::PLEN{1'b0}}, lsu_paddr_o}, 1'b1};
            end
        end
    end
    
    pmp #(
        .PLEN       ( riscv::PLEN            ),
        .PMP_LEN    ( riscv::PLEN - 2        ),
        .NR_ENTRIES ( ArianeCfg.NrPMPEntries )
    ) i_pmp_data (
        .addr_i        ( lsu_paddr_o         ),
        .priv_lvl_i    ( ld_st_priv_lvl_i    ),
        .access_type_i ( pmp_access_type     ),
        
        .conf_addr_i   ( pmpaddr_i           ),
        .conf_i        ( pmpcfg_i            ),
        .allow_o       ( pmp_data_allow      )
    );
    
    
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (~rst_ni) begin
            lsu_vaddr_q      <= '0;
            lsu_req_q        <= '0;
            misaligned_ex_q  <= '0;
            dtlb_pte_q       <= '0;
            dtlb_hit_q       <= '0;
            lsu_is_store_q   <= '0;
            dtlb_is_2M_q     <= '0;
            dtlb_is_1G_q     <= '0;
        end else begin
            lsu_vaddr_q      <=  lsu_vaddr_n;
            lsu_req_q        <=  lsu_req_n;
            misaligned_ex_q  <=  misaligned_ex_n;
            dtlb_pte_q       <=  dtlb_pte_n;
            dtlb_hit_q       <=  dtlb_hit_n;
            lsu_is_store_q   <=  lsu_is_store_n;
            dtlb_is_2M_q     <=  dtlb_is_2M_n;
            dtlb_is_1G_q     <=  dtlb_is_1G_n;
        end
    end
endmodule
module cva6_mmu_sv32 import ariane_pkg::*; #(
    parameter int unsigned INSTR_TLB_ENTRIES     = 4,
    parameter int unsigned DATA_TLB_ENTRIES      = 4,
    parameter int unsigned ASID_WIDTH            = 1,
    parameter ariane_pkg::ariane_cfg_t ArianeCfg = ariane_pkg::ArianeDefaultConfig
) (
    input  logic                            clk_i,
    input  logic                            rst_ni,
    input  logic                            flush_i,
    input  logic                            enable_translation_i,
    input  logic                            en_ld_st_translation_i,   
    
    input  icache_areq_o_t                  icache_areq_i,
    output icache_areq_i_t                  icache_areq_o,
    
    
    
    input  exception_t                      misaligned_ex_i,
    input  logic                            lsu_req_i,        
    input  logic [riscv::VLEN-1:0]          lsu_vaddr_i,      
    input  logic                            lsu_is_store_i,   
    
    
    output logic                            lsu_dtlb_hit_o,   
    output logic [riscv::PPNW-1:0]          lsu_dtlb_ppn_o,   
    
    output logic                            lsu_valid_o,      
    output logic [riscv::PLEN-1:0]          lsu_paddr_o,      
    output exception_t                      lsu_exception_o,  
    
    input riscv::priv_lvl_t                 priv_lvl_i,
    input riscv::priv_lvl_t                 ld_st_priv_lvl_i,
    input logic                             sum_i,
    input logic                             mxr_i,
    
    input logic [riscv::PPNW-1:0]           satp_ppn_i,
    input logic [ASID_WIDTH-1:0]            asid_i,
    input logic [ASID_WIDTH-1:0]            asid_to_be_flushed_i,
    input logic [riscv::VLEN-1:0]           vaddr_to_be_flushed_i,
    input logic                             flush_tlb_i,
    
    output logic                            itlb_miss_o,
    output logic                            dtlb_miss_o,
    
    input  dcache_req_o_t                   req_port_i,
    output dcache_req_i_t                   req_port_o,
    
    input  riscv::pmpcfg_t [15:0]           pmpcfg_i,
    input  logic [15:0][riscv::PLEN-3:0]    pmpaddr_i
);
    logic                   iaccess_err;   
    logic                   daccess_err;   
    logic                   ptw_active;    
    logic                   walking_instr; 
    logic                   ptw_error;     
    logic                   ptw_access_exception; 
    logic [riscv::PLEN-1:0] ptw_bad_paddr; 
    logic [riscv::VLEN-1:0] update_vaddr;
    tlb_update_sv32_t update_ptw_itlb, update_ptw_dtlb;
    logic             itlb_lu_access;
    riscv::pte_sv32_t itlb_content;
    logic             itlb_is_4M;
    logic             itlb_lu_hit;
    logic             dtlb_lu_access;
    riscv::pte_sv32_t dtlb_content;
    logic             dtlb_is_4M;
    logic             dtlb_lu_hit;
    
    assign itlb_lu_access = icache_areq_i.fetch_req;
    assign dtlb_lu_access = lsu_req_i;
    cva6_tlb_sv32 #(
        .TLB_ENTRIES      ( INSTR_TLB_ENTRIES          ),
        .ASID_WIDTH       ( ASID_WIDTH                 )
    ) i_itlb (
        .clk_i            ( clk_i                      ),
        .rst_ni           ( rst_ni                     ),
        .flush_i          ( flush_tlb_i                ),
        .update_i         ( update_ptw_itlb            ),
        .lu_access_i      ( itlb_lu_access             ),
        .lu_asid_i        ( asid_i                     ),
        .asid_to_be_flushed_i  ( asid_to_be_flushed_i  ),
        .vaddr_to_be_flushed_i ( vaddr_to_be_flushed_i ),
        .lu_vaddr_i       ( icache_areq_i.fetch_vaddr  ),
        .lu_content_o     ( itlb_content               ),
        .lu_is_4M_o       ( itlb_is_4M                 ),
        .lu_hit_o         ( itlb_lu_hit                )
    );
    cva6_tlb_sv32 #(
        .TLB_ENTRIES     ( DATA_TLB_ENTRIES             ),
        .ASID_WIDTH      ( ASID_WIDTH                   )
    ) i_dtlb (
        .clk_i            ( clk_i                       ),
        .rst_ni           ( rst_ni                      ),
        .flush_i          ( flush_tlb_i                 ),
        .update_i         ( update_ptw_dtlb             ),
        .lu_access_i      ( dtlb_lu_access              ),
        .lu_asid_i        ( asid_i                      ),
        .asid_to_be_flushed_i  ( asid_to_be_flushed_i   ),
        .vaddr_to_be_flushed_i ( vaddr_to_be_flushed_i  ),
        .lu_vaddr_i       ( lsu_vaddr_i                 ),
        .lu_content_o     ( dtlb_content                ),
        .lu_is_4M_o       ( dtlb_is_4M                  ),
        .lu_hit_o         ( dtlb_lu_hit                 )
    );
    cva6_ptw_sv32  #(
        .ASID_WIDTH             ( ASID_WIDTH            ),
        .ArianeCfg              ( ArianeCfg             )
    ) i_ptw (
        .clk_i                  ( clk_i                 ),
        .rst_ni                 ( rst_ni                ),
        .ptw_active_o           ( ptw_active            ),
        .walking_instr_o        ( walking_instr         ),
        .ptw_error_o            ( ptw_error             ),
        .ptw_access_exception_o ( ptw_access_exception  ),
        .enable_translation_i   ( enable_translation_i  ),
        .update_vaddr_o         ( update_vaddr          ),
        .itlb_update_o          ( update_ptw_itlb       ),
        .dtlb_update_o          ( update_ptw_dtlb       ),
        .itlb_access_i          ( itlb_lu_access        ),
        .itlb_hit_i             ( itlb_lu_hit           ),
        .itlb_vaddr_i           ( icache_areq_i.fetch_vaddr ),
        .dtlb_access_i          ( dtlb_lu_access        ),
        .dtlb_hit_i             ( dtlb_lu_hit           ),
        .dtlb_vaddr_i           ( lsu_vaddr_i           ),
        .req_port_i             ( req_port_i            ),
        .req_port_o             ( req_port_o            ),
        .pmpcfg_i,
        .pmpaddr_i,
        .bad_paddr_o            ( ptw_bad_paddr         ),
        .*
    );
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    logic match_any_execute_region;
    logic pmp_instr_allow;
    
    always_comb begin : instr_interface
        
        icache_areq_o.fetch_valid  = icache_areq_i.fetch_req;
        icache_areq_o.fetch_paddr  = {{riscv::PLEN-riscv::VLEN{1'b0}}, icache_areq_i.fetch_vaddr};
        
        
        
        icache_areq_o.fetch_exception      = '0;
        
        iaccess_err   = icache_areq_i.fetch_req && (((priv_lvl_i == riscv::PRIV_LVL_U) && ~itlb_content.u)
                                                 || ((priv_lvl_i == riscv::PRIV_LVL_S) && itlb_content.u));
        
        
        
        
        if (enable_translation_i) begin
            
            if (icache_areq_i.fetch_req && !((&icache_areq_i.fetch_vaddr[riscv::VLEN-1:riscv::SV-1]) == 1'b1 || (|icache_areq_i.fetch_vaddr[riscv::VLEN-1:riscv::SV-1]) == 1'b0)) begin
                icache_areq_o.fetch_exception = {riscv::INSTR_ACCESS_FAULT, {{riscv::XLEN-riscv::VLEN{1'b0}}, icache_areq_i.fetch_vaddr}, 1'b1};
            end
            icache_areq_o.fetch_valid = 1'b0;
            
            icache_areq_o.fetch_paddr = {itlb_content.ppn, icache_areq_i.fetch_vaddr[11:0]};
            
            if (itlb_is_4M) begin
                icache_areq_o.fetch_paddr[21:12] = icache_areq_i.fetch_vaddr[21:12];
            end
            
            
            
            
            if (itlb_lu_hit) begin
                icache_areq_o.fetch_valid = icache_areq_i.fetch_req;
                
                if (iaccess_err) begin
                    
                    icache_areq_o.fetch_exception = {riscv::INSTR_PAGE_FAULT, {{riscv::XLEN-riscv::VLEN{1'b0}}, icache_areq_i.fetch_vaddr}, 1'b1};
                end else if (!pmp_instr_allow) begin
                    icache_areq_o.fetch_exception = {riscv::INSTR_ACCESS_FAULT, icache_areq_i.fetch_vaddr, 1'b1};
                end
            end else
            
            
            
            
            if (ptw_active && walking_instr) begin
                icache_areq_o.fetch_valid = ptw_error | ptw_access_exception;
                if (ptw_error) icache_areq_o.fetch_exception = {riscv::INSTR_PAGE_FAULT, {{riscv::XLEN-riscv::VLEN{1'b0}}, update_vaddr}, 1'b1};
                
                else icache_areq_o.fetch_exception = {riscv::INSTR_ACCESS_FAULT, ptw_bad_paddr[riscv::PLEN-1:2], 1'b1};
            end
        end
        
        
        if (!match_any_execute_region || (!enable_translation_i && !pmp_instr_allow)) begin
          icache_areq_o.fetch_exception = {riscv::INSTR_ACCESS_FAULT, icache_areq_o.fetch_paddr[riscv::PLEN-1:2], 1'b1};
        end
    end
    
    assign match_any_execute_region = ariane_pkg::is_inside_execute_regions(ArianeCfg, {{64-riscv::PLEN{1'b0}}, icache_areq_o.fetch_paddr});
    
    pmp #(
        .PLEN       ( riscv::PLEN            ),
        .PMP_LEN    ( riscv::PLEN - 2        ),
        .NR_ENTRIES ( ArianeCfg.NrPMPEntries )
    ) i_pmp_if (
        .addr_i        ( icache_areq_o.fetch_paddr ),
        .priv_lvl_i,
        
        .access_type_i ( riscv::ACCESS_EXEC        ),
        
        .conf_addr_i   ( pmpaddr_i                 ),
        .conf_i        ( pmpcfg_i                  ),
        .allow_o       ( pmp_instr_allow           )
    );
    
    
    
    logic [riscv::VLEN-1:0] lsu_vaddr_n,     lsu_vaddr_q;
    riscv::pte_sv32_t dtlb_pte_n,      dtlb_pte_q;
    exception_t  misaligned_ex_n, misaligned_ex_q;
    logic        lsu_req_n,       lsu_req_q;
    logic        lsu_is_store_n,  lsu_is_store_q;
    logic        dtlb_hit_n,      dtlb_hit_q;
    logic        dtlb_is_4M_n,    dtlb_is_4M_q;
    
    assign lsu_dtlb_hit_o = (en_ld_st_translation_i) ? dtlb_lu_hit :  1'b1;
    
    riscv::pmp_access_t pmp_access_type;
    logic        pmp_data_allow;
    localparam   PPNWMin = (riscv::PPNW-1 > 29) ? 29 : riscv::PPNW-1;
    
    always_comb begin : data_interface
        
        lsu_vaddr_n           = lsu_vaddr_i;
        lsu_req_n             = lsu_req_i;
        misaligned_ex_n       = misaligned_ex_i;
        dtlb_pte_n            = dtlb_content;
        dtlb_hit_n            = dtlb_lu_hit;
        lsu_is_store_n        = lsu_is_store_i;
        dtlb_is_4M_n          = dtlb_is_4M;
        lsu_paddr_o           = {{riscv::PLEN-riscv::VLEN{1'b0}}, lsu_vaddr_q};
        lsu_dtlb_ppn_o        = {{riscv::PLEN-riscv::VLEN{1'b0}},lsu_vaddr_n[riscv::VLEN-1:12]};
        lsu_valid_o           = lsu_req_q;
        lsu_exception_o       = misaligned_ex_q;
        pmp_access_type       = lsu_is_store_q ? riscv::ACCESS_WRITE : riscv::ACCESS_READ;
        
        misaligned_ex_n.valid = misaligned_ex_i.valid & lsu_req_i;
        
        
        daccess_err = (ld_st_priv_lvl_i == riscv::PRIV_LVL_S && !sum_i && dtlb_pte_q.u) || 
                      (ld_st_priv_lvl_i == riscv::PRIV_LVL_U && !dtlb_pte_q.u);            
        
        if (en_ld_st_translation_i && !misaligned_ex_q.valid) begin
            lsu_valid_o = 1'b0;
            
            lsu_paddr_o = {dtlb_pte_q.ppn, lsu_vaddr_q[11:0]};
            lsu_dtlb_ppn_o = dtlb_content.ppn;
            
            if (dtlb_is_4M_q) begin
              lsu_paddr_o[21:12] = lsu_vaddr_q[21:12];
              lsu_dtlb_ppn_o[21:12] = lsu_vaddr_n[21:12];
            end
            
            
            
            if (dtlb_hit_q && lsu_req_q) begin
                lsu_valid_o = 1'b1;
                
                
                
                
                
                if (lsu_is_store_q) begin
                    
                    
                    if (!dtlb_pte_q.w || daccess_err || !dtlb_pte_q.d) begin
                        lsu_exception_o = {riscv::STORE_PAGE_FAULT, {{riscv::XLEN-riscv::VLEN{lsu_vaddr_q[riscv::VLEN-1]}},lsu_vaddr_q}, 1'b1}; 
                    
                    end else if (!pmp_data_allow) begin
                        lsu_exception_o = {riscv::ST_ACCESS_FAULT, lsu_paddr_o[riscv::PLEN-1:2], 1'b1}; 
                    end
                
                end else begin
                    
                    if (daccess_err) begin
                        lsu_exception_o = {riscv::LOAD_PAGE_FAULT, {{riscv::XLEN-riscv::VLEN{lsu_vaddr_q[riscv::VLEN-1]}},lsu_vaddr_q}, 1'b1};
                    
                    end else if (!pmp_data_allow) begin
                        lsu_exception_o = {riscv::LD_ACCESS_FAULT, lsu_paddr_o[riscv::PLEN-1:2], 1'b1}; 
                    end
                end
            end else
            
            
            
            
            if (ptw_active && !walking_instr) begin
                
                if (ptw_error) begin
                    
                    lsu_valid_o = 1'b1;
                    
                    if (lsu_is_store_q) begin
                        lsu_exception_o = {riscv::STORE_PAGE_FAULT, {{riscv::XLEN-riscv::VLEN{lsu_vaddr_q[riscv::VLEN-1]}},update_vaddr}, 1'b1};
                    end else begin
                        lsu_exception_o = {riscv::LOAD_PAGE_FAULT, {{riscv::XLEN-riscv::VLEN{lsu_vaddr_q[riscv::VLEN-1]}},update_vaddr}, 1'b1};
                    end
                end
                if (ptw_access_exception) begin
                    
                    lsu_valid_o = 1'b1;
                    
                    lsu_exception_o = {riscv::LD_ACCESS_FAULT, ptw_bad_paddr[riscv::PLEN-1:2], 1'b1};
                end
            end
        end
        
        else if (lsu_req_q && !misaligned_ex_q.valid && !pmp_data_allow) begin
            if (lsu_is_store_q) begin
                lsu_exception_o = {riscv::ST_ACCESS_FAULT, lsu_paddr_o[riscv::PLEN-1:2], 1'b1};
            end else begin
                lsu_exception_o = {riscv::LD_ACCESS_FAULT, lsu_paddr_o[riscv::PLEN-1:2], 1'b1};
            end
        end
    end
    
    pmp #(
        .PLEN       ( riscv::PLEN            ),
        .PMP_LEN    ( riscv::PLEN - 2        ),
        .NR_ENTRIES ( ArianeCfg.NrPMPEntries )
    ) i_pmp_data (
        .addr_i        ( lsu_paddr_o         ),
        .priv_lvl_i    ( ld_st_priv_lvl_i    ),
        .access_type_i ( pmp_access_type     ),
        
        .conf_addr_i   ( pmpaddr_i           ),
        .conf_i        ( pmpcfg_i            ),
        .allow_o       ( pmp_data_allow      )
    );
    
    
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (~rst_ni) begin
            lsu_vaddr_q      <= '0;
            lsu_req_q        <= '0;
            misaligned_ex_q  <= '0;
            dtlb_pte_q       <= '0;
            dtlb_hit_q       <= '0;
            lsu_is_store_q   <= '0;
            dtlb_is_4M_q     <= '0;
        end else begin
            lsu_vaddr_q      <=  lsu_vaddr_n;
            lsu_req_q        <=  lsu_req_n;
            misaligned_ex_q  <=  misaligned_ex_n;
            dtlb_pte_q       <=  dtlb_pte_n;
            dtlb_hit_q       <=  dtlb_hit_n;
            lsu_is_store_q   <=  lsu_is_store_n;
            dtlb_is_4M_q     <=  dtlb_is_4M_n;
        end
    end
endmodule
module mult import ariane_pkg::*; (
    input  logic                     clk_i,
    input  logic                     rst_ni,
    input  logic                     flush_i,
    input  fu_data_t                 fu_data_i,
    input  logic                     mult_valid_i,
    output riscv::xlen_t             result_o,
    output logic                     mult_valid_o,
    output logic                     mult_ready_o,
    output logic [TRANS_ID_BITS-1:0] mult_trans_id_o
);
    logic                     mul_valid;
    logic                     div_valid;
    logic                     div_ready_i; 
    logic [TRANS_ID_BITS-1:0] mul_trans_id;
    logic [TRANS_ID_BITS-1:0] div_trans_id;
    riscv::xlen_t             mul_result;
    riscv::xlen_t             div_result;
    logic                     div_valid_op;
    logic                     mul_valid_op;
    
    assign mul_valid_op = ~flush_i && mult_valid_i && (fu_data_i.operator inside { MUL, MULH, MULHU, MULHSU, MULW });
    assign div_valid_op = ~flush_i && mult_valid_i && (fu_data_i.operator inside { DIV, DIVU, DIVW, DIVUW, REM, REMU, REMW, REMUW });
    
    
    
    
    
    assign div_ready_i      = (mul_valid) ? 1'b0         : 1'b1;
    assign mult_trans_id_o  = (mul_valid) ? mul_trans_id : div_trans_id;
    assign result_o         = (mul_valid) ? mul_result   : div_result;
    assign mult_valid_o     = div_valid | mul_valid;
    
    
    
    
    multiplier i_multiplier (
        .clk_i,
        .rst_ni,
        .trans_id_i        ( fu_data_i.trans_id  ),
        .operator_i        ( fu_data_i.operator  ),
        .operand_a_i       ( fu_data_i.operand_a ),
        .operand_b_i       ( fu_data_i.operand_b ),
        .result_o          ( mul_result   ),
        .mult_valid_i      ( mul_valid_op ),
        .mult_valid_o      ( mul_valid    ),
        .mult_trans_id_o   ( mul_trans_id ),
        .mult_ready_o      (              ) 
    );
    
    
    
    riscv::xlen_t           operand_b, operand_a;  
    riscv::xlen_t           result;                
    logic        div_signed;            
    logic        rem;                   
    logic        word_op_d, word_op_q;  
    
    assign div_signed = fu_data_i.operator inside {DIV, DIVW, REM, REMW};
    
    assign rem        = fu_data_i.operator inside {REM, REMU, REMW, REMUW};
    
    always_comb begin
        
        operand_a   = '0;
        operand_b   = '0;
        
        word_op_d   = word_op_q;
        
        if (mult_valid_i && fu_data_i.operator inside {DIV, DIVU, DIVW, DIVUW, REM, REMU, REMW, REMUW}) begin
            
            if (fu_data_i.operator inside {DIVW, DIVUW, REMW, REMUW}) begin
                
                if (div_signed) begin
                    operand_a = sext32(fu_data_i.operand_a[31:0]);
                    operand_b = sext32(fu_data_i.operand_b[31:0]);
                end else begin
                    operand_a = fu_data_i.operand_a[31:0];
                    operand_b = fu_data_i.operand_b[31:0];
                end
                
                word_op_d = 1'b1;
            end else begin
                
                operand_a = fu_data_i.operand_a;
                operand_b = fu_data_i.operand_b;
                word_op_d = 1'b0;
            end
        end
    end
    
    
    
    serdiv #(
        .WIDTH       ( riscv::XLEN )
    ) i_div (
        .clk_i       ( clk_i                ),
        .rst_ni      ( rst_ni               ),
        .id_i        ( fu_data_i.trans_id   ),
        .op_a_i      ( operand_a            ),
        .op_b_i      ( operand_b            ),
        .opcode_i    ( {rem, div_signed}    ), 
        .in_vld_i    ( div_valid_op         ),
        .in_rdy_o    ( mult_ready_o         ),
        .flush_i     ( flush_i              ),
        .out_vld_o   ( div_valid            ),
        .out_rdy_i   ( div_ready_i          ),
        .id_o        ( div_trans_id         ),
        .res_o       ( result               )
    );
    
    
    assign div_result = (word_op_q) ? sext32(result) : result;
    
    
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if(~rst_ni) begin
            word_op_q <= '0;
        end else begin
            word_op_q <= word_op_d;
        end
    end
endmodule
module multiplier import ariane_pkg::*; (
    input  logic                     clk_i,
    input  logic                     rst_ni,
    input  logic [TRANS_ID_BITS-1:0] trans_id_i,
    input  logic                     mult_valid_i,
    input  fu_op                     operator_i,
    input  riscv::xlen_t             operand_a_i,
    input  riscv::xlen_t             operand_b_i,
    output riscv::xlen_t             result_o,
    output logic                     mult_valid_o,
    output logic                     mult_ready_o,
    output logic [TRANS_ID_BITS-1:0] mult_trans_id_o
);
    
    logic [TRANS_ID_BITS-1:0]    trans_id_q;
    logic                        mult_valid_q;
    fu_op                        operator_d, operator_q;
    logic [riscv::XLEN*2-1:0] mult_result_d, mult_result_q;
    
    logic                       sign_a, sign_b;
    logic                       mult_valid;
    
    assign mult_valid_o    = mult_valid_q;
    assign mult_trans_id_o = trans_id_q;
    assign mult_ready_o    = 1'b1;
    assign mult_valid      = mult_valid_i && (operator_i inside {MUL, MULH, MULHU, MULHSU, MULW});
    
    logic [riscv::XLEN*2-1:0] mult_result;
    assign mult_result   = $signed({operand_a_i[riscv::XLEN-1] & sign_a, operand_a_i}) * $signed({operand_b_i[riscv::XLEN-1] & sign_b, operand_b_i});
    
    always_comb begin
        sign_a = 1'b0;
        sign_b = 1'b0;
        
        if (operator_i == MULH) begin
            sign_a   = 1'b1;
            sign_b   = 1'b1;
        
        end else if (operator_i == MULHSU) begin
            sign_a   = 1'b1;
        
        end else begin
            sign_a   = 1'b0;
            sign_b   = 1'b0;
        end
    end
    
    assign mult_result_d   = $signed({operand_a_i[riscv::XLEN-1] & sign_a, operand_a_i}) *
                             $signed({operand_b_i[riscv::XLEN-1] & sign_b, operand_b_i});
    assign operator_d = operator_i;
    always_comb begin : p_selmux
        unique case (operator_q)
            MULH, MULHU, MULHSU: result_o = mult_result_q[riscv::XLEN*2-1:riscv::XLEN];
            MULW:                result_o = sext32(mult_result_q[31:0]);
            
            default:             result_o = mult_result_q[riscv::XLEN-1:0];
        endcase
    end
    
    
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (~rst_ni) begin
            mult_valid_q    <= '0;
            trans_id_q      <= '0;
            operator_q      <=  MUL;
            mult_result_q   <= '0;
         end else begin
            
            trans_id_q   <= trans_id_i;
            
            mult_valid_q    <= mult_valid;
            operator_q      <= operator_d;
            mult_result_q   <= mult_result_d;
         end
    end
endmodule
module serdiv import ariane_pkg::*; #(
  parameter WIDTH       = 64
) (
  input  logic                      clk_i,
  input  logic                      rst_ni,
  
  input  logic [TRANS_ID_BITS-1:0]  id_i,
  input  logic [WIDTH-1:0]          op_a_i,
  input  logic [WIDTH-1:0]          op_b_i,
  input  logic [1:0]                opcode_i, 
  
  input  logic                      in_vld_i, 
  output logic                      in_rdy_o,
  input  logic                      flush_i,
  
  output logic                      out_vld_o,
  input  logic                      out_rdy_i,
  output logic [TRANS_ID_BITS-1:0]  id_o,
  output logic [WIDTH-1:0]          res_o
);
  enum logic [1:0] {IDLE, DIVIDE, FINISH} state_d, state_q;
  logic [WIDTH-1:0]       res_q, res_d;
  logic [WIDTH-1:0]       op_a_q, op_a_d;
  logic [WIDTH-1:0]       op_b_q, op_b_d;
  logic                   op_a_sign, op_b_sign;
  logic                   op_b_zero, op_b_zero_q, op_b_zero_d;
  logic [TRANS_ID_BITS-1:0] id_q, id_d;
  logic rem_sel_d, rem_sel_q;
  logic comp_inv_d, comp_inv_q;
  logic res_inv_d, res_inv_q;
  logic [WIDTH-1:0] add_mux;
  logic [WIDTH-1:0] add_out;
  logic [WIDTH-1:0] add_tmp;
  logic [WIDTH-1:0] b_mux;
  logic [WIDTH-1:0] out_mux;
  logic [$clog2(WIDTH+1)-1:0] cnt_q, cnt_d;
  logic cnt_zero;
  logic [WIDTH-1:0] lzc_a_input, lzc_b_input, op_b;
  logic [$clog2(WIDTH)-1:0] lzc_a_result, lzc_b_result;
  logic [$clog2(WIDTH+1)-1:0] shift_a;
  logic [$clog2(WIDTH+1):0] div_shift;
  logic a_reg_en, b_reg_en, res_reg_en, ab_comp, pm_sel, load_en;
  logic lzc_a_no_one, lzc_b_no_one;
  logic div_res_zero_d, div_res_zero_q;
  assign op_b_zero = (op_b_i == 0);
  assign op_a_sign = op_a_i[$high(op_a_i)];
  assign op_b_sign = op_b_i[$high(op_b_i)];
  assign lzc_a_input = (opcode_i[0] & op_a_sign) ? {~op_a_i, 1'b0} : op_a_i;
  assign lzc_b_input = (opcode_i[0] & op_b_sign) ? ~op_b_i         : op_b_i;
  lzc #(
    .MODE    ( 1          ), 
    .WIDTH   ( WIDTH      )
  ) i_lzc_a (
    .in_i    ( lzc_a_input  ),
    .cnt_o   ( lzc_a_result ),
    .empty_o ( lzc_a_no_one )
  );
  lzc #(
    .MODE    ( 1          ), 
    .WIDTH   ( WIDTH      )
  ) i_lzc_b (
    .in_i    ( lzc_b_input  ),
    .cnt_o   ( lzc_b_result ),
    .empty_o ( lzc_b_no_one )
  );
  assign shift_a      = (lzc_a_no_one) ? WIDTH : lzc_a_result;
  assign div_shift    = (lzc_b_no_one) ? WIDTH : lzc_b_result-shift_a;
  assign op_b         = op_b_i <<< $unsigned(div_shift);
  
  assign div_res_zero_d = (load_en) ? ($signed(div_shift) < 0) : div_res_zero_q;
  assign pm_sel      = load_en & ~(opcode_i[0] & (op_a_sign ^ op_b_sign));
  
  assign add_mux     = (load_en)   ? op_a_i  : op_b_q;
  
  assign b_mux       = (load_en)   ? op_b : {comp_inv_q, (op_b_q[$high(op_b_q):1])};
  
  assign out_mux     = (rem_sel_q) ? op_a_q : res_q;
  
  
  assign res_o       = (res_inv_q) ? -$signed(out_mux) : out_mux;
  
  assign ab_comp     = ((op_a_q == op_b_q) | ((op_a_q > op_b_q) ^ comp_inv_q)) & ((|op_a_q) | op_b_zero_q);
  
  assign add_tmp     = (load_en) ? 0 : op_a_q;
  assign add_out     = (pm_sel)  ? add_tmp + add_mux : add_tmp - $signed(add_mux);
  assign cnt_zero = (cnt_q == 0);
  assign cnt_d    = (load_en)   ? div_shift  :
                    (~cnt_zero) ? cnt_q - 1  : cnt_q;
  always_comb begin : p_fsm
    
    state_d        = state_q;
    in_rdy_o       = 1'b0;
    out_vld_o      = 1'b0;
    load_en        = 1'b0;
    a_reg_en       = 1'b0;
    b_reg_en       = 1'b0;
    res_reg_en     = 1'b0;
    unique case (state_q)
      IDLE: begin
        in_rdy_o    = 1'b1;
        if (in_vld_i) begin
          in_rdy_o  = 1'b0;
          a_reg_en  = 1'b1;
          b_reg_en  = 1'b1;
          load_en   = 1'b1;
          state_d   = DIVIDE;
        end
      end
      DIVIDE: begin
        if(~div_res_zero_q) begin
          a_reg_en     = ab_comp;
          b_reg_en     = 1'b1;
          res_reg_en   = 1'b1;
        end
        
        if(div_res_zero_q) begin
          out_vld_o = 1'b1;
          state_d   = FINISH;
          if(out_rdy_i) begin
            
            state_d  = IDLE;
          end
        end else if (cnt_zero) begin
          state_d   = FINISH;
        end
      end
      FINISH: begin
        out_vld_o = 1'b1;
        if (out_rdy_i) begin
          
          state_d  = IDLE;
        end
      end
      default : state_d = IDLE;
    endcase
    if (flush_i) begin
        in_rdy_o   = 1'b0;
        out_vld_o  = 1'b0;
        a_reg_en   = 1'b0;
        b_reg_en   = 1'b0;
        load_en    = 1'b0;
        state_d    = IDLE;
    end
  end
  
  assign rem_sel_d    = (load_en) ? opcode_i[1]               : rem_sel_q;
  assign comp_inv_d   = (load_en) ? opcode_i[0] & op_b_sign   : comp_inv_q;
  assign op_b_zero_d  = (load_en) ? op_b_zero                 : op_b_zero_q;
  assign res_inv_d    = (load_en) ? (~op_b_zero | opcode_i[1]) & opcode_i[0] & (op_a_sign ^ op_b_sign) : res_inv_q;
  
  assign id_d = (load_en) ? id_i : id_q;
  assign id_o = id_q;
  assign op_a_d   = (a_reg_en)   ? add_out : op_a_q;
  assign op_b_d   = (b_reg_en)   ? b_mux   : op_b_q;
  assign res_d    = (load_en)   ? '0       :
                    (res_reg_en) ? {res_q[$high(res_q)-1:0], ab_comp} : res_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin : p_regs
    if (~rst_ni) begin
      state_q        <= IDLE;
      op_a_q         <= '0;
      op_b_q         <= '0;
      res_q          <= '0;
      cnt_q          <= '0;
      id_q           <= '0;
      rem_sel_q      <= 1'b0;
      comp_inv_q     <= 1'b0;
      res_inv_q      <= 1'b0;
      op_b_zero_q    <= 1'b0;
      div_res_zero_q <= 1'b0;
    end else begin
      state_q        <= state_d;
      op_a_q         <= op_a_d;
      op_b_q         <= op_b_d;
      res_q          <= res_d;
      cnt_q          <= cnt_d;
      id_q           <= id_d;
      rem_sel_q      <= rem_sel_d;
      comp_inv_q     <= comp_inv_d;
      res_inv_q      <= res_inv_d;
      op_b_zero_q    <= op_b_zero_d;
      div_res_zero_q <= div_res_zero_d;
    end
  end
endmodule
module perf_counters import ariane_pkg::*; (
  input  logic                                    clk_i,
  input  logic                                    rst_ni,
  input  logic                                    debug_mode_i, 
  
  input  logic [4:0]                              addr_i,   
  input  logic                                    we_i,     
  input  riscv::xlen_t                            data_i,   
  output riscv::xlen_t                            data_o,   
  
  input  scoreboard_entry_t [NR_COMMIT_PORTS-1:0] commit_instr_i,     
  input  logic [NR_COMMIT_PORTS-1:0]              commit_ack_i,       
  
  input  logic                                    l1_icache_miss_i,
  input  logic                                    l1_dcache_miss_i,
  
  input  logic                                    itlb_miss_i,
  input  logic                                    dtlb_miss_i,
  
  input  logic                                    sb_full_i,
  
  input  logic                                    if_empty_i,
  
  input  exception_t                              ex_i,
  input  logic                                    eret_i,
  input  bp_resolve_t                             resolved_branch_i
);
  localparam logic [6:0] RegOffset = riscv::CSR_ML1_ICACHE_MISS >> 5;
  logic [riscv::CSR_MIF_EMPTY : riscv::CSR_ML1_ICACHE_MISS][riscv::XLEN-1:0] perf_counter_d, perf_counter_q;
  always_comb begin : perf_counters
    perf_counter_d = perf_counter_q;
    data_o = 'b0;
    
    if (!debug_mode_i) begin
      
      
      
      if (l1_icache_miss_i)
        perf_counter_d[riscv::CSR_ML1_ICACHE_MISS] = perf_counter_q[riscv::CSR_ML1_ICACHE_MISS] + 1'b1;
      if (l1_dcache_miss_i)
        perf_counter_d[riscv::CSR_ML1_DCACHE_MISS] = perf_counter_q[riscv::CSR_ML1_DCACHE_MISS] + 1'b1;
      if (itlb_miss_i)
        perf_counter_d[riscv::CSR_MITLB_MISS] = perf_counter_q[riscv::CSR_MITLB_MISS] + 1'b1;
      if (dtlb_miss_i)
        perf_counter_d[riscv::CSR_MDTLB_MISS] = perf_counter_q[riscv::CSR_MDTLB_MISS] + 1'b1;
      
      for (int unsigned i = 0; i < NR_COMMIT_PORTS-1; i++) begin
        if (commit_ack_i[i]) begin
          if (commit_instr_i[i].fu == LOAD)
            perf_counter_d[riscv::CSR_MLOAD] = perf_counter_q[riscv::CSR_MLOAD] + 1'b1;
          if (commit_instr_i[i].fu == STORE)
            perf_counter_d[riscv::CSR_MSTORE] = perf_counter_q[riscv::CSR_MSTORE] + 1'b1;
          if (commit_instr_i[i].fu == CTRL_FLOW)
            perf_counter_d[riscv::CSR_MBRANCH_JUMP] = perf_counter_q[riscv::CSR_MBRANCH_JUMP] + 1'b1;
          
          
          if (commit_instr_i[i].fu == CTRL_FLOW && commit_instr_i[i].op == '0
                                                && (commit_instr_i[i].rd == 'd1 || commit_instr_i[i].rd == 'd1))
            perf_counter_d[riscv::CSR_MCALL] = perf_counter_q[riscv::CSR_MCALL] + 1'b1;
          
          if (commit_instr_i[i].op == JALR && (commit_instr_i[i].rd == 'd1 || commit_instr_i[i].rd == 'd1))
            perf_counter_d[riscv::CSR_MRET] = perf_counter_q[riscv::CSR_MRET] + 1'b1;
        end
      end
      if (ex_i.valid)
        perf_counter_d[riscv::CSR_MEXCEPTION] = perf_counter_q[riscv::CSR_MEXCEPTION] + 1'b1;
      if (eret_i)
        perf_counter_d[riscv::CSR_MEXCEPTION_RET] = perf_counter_q[riscv::CSR_MEXCEPTION_RET] + 1'b1;
      if (resolved_branch_i.valid && resolved_branch_i.is_mispredict)
        perf_counter_d[riscv::CSR_MMIS_PREDICT] = perf_counter_q[riscv::CSR_MMIS_PREDICT] + 1'b1;
      if (sb_full_i) begin
        perf_counter_d[riscv::CSR_MSB_FULL] = perf_counter_q[riscv::CSR_MSB_FULL] + 1'b1;
      end
      if (if_empty_i) begin
        perf_counter_d[riscv::CSR_MIF_EMPTY] = perf_counter_q[riscv::CSR_MIF_EMPTY] + 1'b1;
      end
    end
    
    data_o = perf_counter_q[{RegOffset,addr_i}];
    if (we_i) begin
      perf_counter_d[{RegOffset,addr_i}] = data_i;
    end
  end
  
  
  
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      perf_counter_q <= '0;
    end else begin
      perf_counter_q <= perf_counter_d;
    end
  end
endmodule
module ptw import ariane_pkg::*; #(
        parameter int ASID_WIDTH = 1,
        parameter ariane_pkg::ariane_cfg_t ArianeCfg = ariane_pkg::ArianeDefaultConfig
) (
    input  logic                    clk_i,                  
    input  logic                    rst_ni,                 
    input  logic                    flush_i,                
                                                            
                                                            
    output logic                    ptw_active_o,
    output logic                    walking_instr_o,        
    output logic                    ptw_error_o,            
    output logic                    ptw_access_exception_o, 
    input  logic                    enable_translation_i,   
    input  logic                    en_ld_st_translation_i, 
    input  logic                    lsu_is_store_i,         
    
    input  dcache_req_o_t           req_port_i,
    output dcache_req_i_t           req_port_o,
    
    output tlb_update_t             itlb_update_o,
    output tlb_update_t             dtlb_update_o,
    output logic [riscv::VLEN-1:0]  update_vaddr_o,
    input  logic [ASID_WIDTH-1:0]   asid_i,
    
    
    input  logic                    itlb_access_i,
    input  logic                    itlb_hit_i,
    input  logic [riscv::VLEN-1:0]  itlb_vaddr_i,
    input  logic                    dtlb_access_i,
    input  logic                    dtlb_hit_i,
    input  logic [riscv::VLEN-1:0]  dtlb_vaddr_i,
    
    input  logic [riscv::PPNW-1:0]  satp_ppn_i, 
    input  logic                    mxr_i,
    
    output logic                    itlb_miss_o,
    output logic                    dtlb_miss_o,
    
    input  riscv::pmpcfg_t [15:0]   pmpcfg_i,
    input  logic [15:0][riscv::PLEN-3:0] pmpaddr_i,
    output logic [riscv::PLEN-1:0]  bad_paddr_o
);
    
    logic data_rvalid_q;
    logic [63:0] data_rdata_q;
    riscv::pte_t pte;
    assign pte = riscv::pte_t'(data_rdata_q);
    enum logic[2:0] {
      IDLE,
      WAIT_GRANT,
      PTE_LOOKUP,
      WAIT_RVALID,
      PROPAGATE_ERROR,
      PROPAGATE_ACCESS_ERROR
    } state_q, state_d;
    
    enum logic [1:0] {
        LVL1, LVL2, LVL3
    } ptw_lvl_q, ptw_lvl_n;
    
    logic is_instr_ptw_q,   is_instr_ptw_n;
    logic global_mapping_q, global_mapping_n;
    
    logic tag_valid_n,      tag_valid_q;
    
    logic [ASID_WIDTH-1:0]  tlb_update_asid_q, tlb_update_asid_n;
    
    logic [riscv::VLEN-1:0] vaddr_q,   vaddr_n;
    
    logic [riscv::PLEN-1:0] ptw_pptr_q, ptw_pptr_n;
    
    assign update_vaddr_o  = vaddr_q;
    assign ptw_active_o    = (state_q != IDLE);
    assign walking_instr_o = is_instr_ptw_q;
    
    assign req_port_o.address_index = ptw_pptr_q[DCACHE_INDEX_WIDTH-1:0];
    assign req_port_o.address_tag   = ptw_pptr_q[DCACHE_INDEX_WIDTH+DCACHE_TAG_WIDTH-1:DCACHE_INDEX_WIDTH];
    
    assign req_port_o.kill_req      = '0;
    
    assign req_port_o.data_wdata    = 64'b0;
    
    
    
    assign itlb_update_o.vpn = {{39-riscv::SV{1'b0}}, vaddr_q[riscv::SV-1:12]};
    assign dtlb_update_o.vpn = {{39-riscv::SV{1'b0}}, vaddr_q[riscv::SV-1:12]};
    
    assign itlb_update_o.is_2M = (ptw_lvl_q == LVL2);
    assign itlb_update_o.is_1G = (ptw_lvl_q == LVL1);
    assign dtlb_update_o.is_2M = (ptw_lvl_q == LVL2);
    assign dtlb_update_o.is_1G = (ptw_lvl_q == LVL1);
    
    assign itlb_update_o.asid = tlb_update_asid_q;
    assign dtlb_update_o.asid = tlb_update_asid_q;
    
    assign itlb_update_o.content = pte | (global_mapping_q << 5);
    assign dtlb_update_o.content = pte | (global_mapping_q << 5);
    assign req_port_o.tag_valid      = tag_valid_q;
    logic allow_access;
    assign bad_paddr_o = ptw_access_exception_o ? ptw_pptr_q : 'b0;
    pmp #(
        .PLEN       ( riscv::PLEN            ),
        .PMP_LEN    ( riscv::PLEN - 2        ),
        .NR_ENTRIES ( ArianeCfg.NrPMPEntries )
    ) i_pmp_ptw (
        .addr_i        ( ptw_pptr_q         ),
        
        .priv_lvl_i    ( riscv::PRIV_LVL_S  ),
        
        .access_type_i ( riscv::ACCESS_READ ),
        
        .conf_addr_i   ( pmpaddr_i          ),
        .conf_i        ( pmpcfg_i           ),
        .allow_o       ( allow_access       )
    );
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    always_comb begin : ptw
        
        
        tag_valid_n            = 1'b0;
        req_port_o.data_req    = 1'b0;
        req_port_o.data_be     = 8'hFF;
        req_port_o.data_size   = 2'b11;
        req_port_o.data_we     = 1'b0;
        ptw_error_o            = 1'b0;
        ptw_access_exception_o = 1'b0;
        itlb_update_o.valid    = 1'b0;
        dtlb_update_o.valid    = 1'b0;
        is_instr_ptw_n         = is_instr_ptw_q;
        ptw_lvl_n              = ptw_lvl_q;
        ptw_pptr_n             = ptw_pptr_q;
        state_d                = state_q;
        global_mapping_n       = global_mapping_q;
        
        tlb_update_asid_n     = tlb_update_asid_q;
        vaddr_n               = vaddr_q;
        itlb_miss_o           = 1'b0;
        dtlb_miss_o           = 1'b0;
        case (state_q)
            IDLE: begin
                
                ptw_lvl_n        = LVL1;
                global_mapping_n = 1'b0;
                is_instr_ptw_n   = 1'b0;
                
                if (enable_translation_i & itlb_access_i & ~itlb_hit_i & ~dtlb_access_i) begin
                    ptw_pptr_n          = {satp_ppn_i, itlb_vaddr_i[riscv::SV-1:30], 3'b0};
                    is_instr_ptw_n      = 1'b1;
                    tlb_update_asid_n   = asid_i;
                    vaddr_n             = itlb_vaddr_i;
                    state_d             = WAIT_GRANT;
                    itlb_miss_o         = 1'b1;
                
                end else if (en_ld_st_translation_i & dtlb_access_i & ~dtlb_hit_i) begin
                    ptw_pptr_n          = {satp_ppn_i, dtlb_vaddr_i[riscv::SV-1:30], 3'b0};
                    tlb_update_asid_n   = asid_i;
                    vaddr_n             = dtlb_vaddr_i;
                    state_d             = WAIT_GRANT;
                    dtlb_miss_o         = 1'b1;
                end
            end
            WAIT_GRANT: begin
                
                req_port_o.data_req = 1'b1;
                
                if (req_port_i.data_gnt) begin
                    
                    tag_valid_n = 1'b1;
                    state_d     = PTE_LOOKUP;
                end
            end
            PTE_LOOKUP: begin
                
                if (data_rvalid_q) begin
                    
                    if (pte.g)
                        global_mapping_n = 1'b1;
                    
                    
                    
                    
                    if (!pte.v || (!pte.r && pte.w))
                        state_d = PROPAGATE_ERROR;
                    
                    
                    
                    else begin
                        state_d = IDLE;
                        
                        
                        if (pte.r || pte.x) begin
                            
                            if (is_instr_ptw_q) begin
                                
                                
                                
                                
                                
                                
                                if (!pte.x || !pte.a)
                                  state_d = PROPAGATE_ERROR;
                                else
                                  itlb_update_o.valid = 1'b1;
                            end else begin
                                
                                
                                
                                
                                
                                
                                
                                
                                if (pte.a && (pte.r || (pte.x && mxr_i))) begin
                                  dtlb_update_o.valid = 1'b1;
                                end else begin
                                  state_d   = PROPAGATE_ERROR;
                                end
                                
                                
                                
                                if (lsu_is_store_i && (!pte.w || !pte.d)) begin
                                    dtlb_update_o.valid = 1'b0;
                                    state_d   = PROPAGATE_ERROR;
                                end
                            end
                            
                            
                            
                            if (ptw_lvl_q == LVL1 && pte.ppn[17:0] != '0) begin
                                state_d             = PROPAGATE_ERROR;
                                dtlb_update_o.valid = 1'b0;
                                itlb_update_o.valid = 1'b0;
                            end else if (ptw_lvl_q == LVL2 && pte.ppn[8:0] != '0) begin
                                state_d             = PROPAGATE_ERROR;
                                dtlb_update_o.valid = 1'b0;
                                itlb_update_o.valid = 1'b0;
                            end
                        
                        end else begin
                            
                            if (ptw_lvl_q == LVL1) begin
                                
                                ptw_lvl_n  = LVL2;
                                ptw_pptr_n = {pte.ppn, vaddr_q[29:21], 3'b0};
                            end
                            if (ptw_lvl_q == LVL2) begin
                                
                                ptw_lvl_n  = LVL3;
                                ptw_pptr_n = {pte.ppn, vaddr_q[20:12], 3'b0};
                            end
                            state_d = WAIT_GRANT;
                            if (ptw_lvl_q == LVL3) begin
                              
                              ptw_lvl_n   = LVL3;
                              state_d = PROPAGATE_ERROR;
                            end
                        end
                    end
                    
                    if (!allow_access) begin
                        itlb_update_o.valid = 1'b0;
                        dtlb_update_o.valid = 1'b0;
                        
                        ptw_pptr_n = ptw_pptr_q;
                        state_d = PROPAGATE_ACCESS_ERROR;
                    end
                end
                
            end
            
            PROPAGATE_ERROR: begin
                state_d     = IDLE;
                ptw_error_o = 1'b1;
            end
            PROPAGATE_ACCESS_ERROR: begin
                state_d     = IDLE;
                ptw_access_exception_o = 1'b1;
            end
            
            WAIT_RVALID: begin
                if (data_rvalid_q)
                    state_d = IDLE;
            end
            default: begin
                state_d = IDLE;
            end
        endcase
        
        
        
        
        if (flush_i) begin
            
            
            
            
            if ((state_q == PTE_LOOKUP && !data_rvalid_q) || ((state_q == WAIT_GRANT) && req_port_i.data_gnt))
                state_d = WAIT_RVALID;
            else
                state_d = IDLE;
        end
    end
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (~rst_ni) begin
            state_q            <= IDLE;
            is_instr_ptw_q     <= 1'b0;
            ptw_lvl_q          <= LVL1;
            tag_valid_q        <= 1'b0;
            tlb_update_asid_q  <= '0;
            vaddr_q            <= '0;
            ptw_pptr_q         <= '0;
            global_mapping_q   <= 1'b0;
            data_rdata_q       <= '0;
            data_rvalid_q      <= 1'b0;
        end else begin
            state_q            <= state_d;
            ptw_pptr_q         <= ptw_pptr_n;
            is_instr_ptw_q     <= is_instr_ptw_n;
            ptw_lvl_q          <= ptw_lvl_n;
            tag_valid_q        <= tag_valid_n;
            tlb_update_asid_q  <= tlb_update_asid_n;
            vaddr_q            <= vaddr_n;
            global_mapping_q   <= global_mapping_n;
            data_rdata_q       <= req_port_i.data_rdata;
            data_rvalid_q      <= req_port_i.data_rvalid;
        end
    end
endmodule
module tlb import ariane_pkg::*; #(
      parameter int unsigned TLB_ENTRIES = 4,
      parameter int unsigned ASID_WIDTH  = 1
  )(
    input  logic                    clk_i,    
    input  logic                    rst_ni,   
    input  logic                    flush_i,  
    
    input  tlb_update_t             update_i,
    
    input  logic                    lu_access_i,
    input  logic [ASID_WIDTH-1:0]   lu_asid_i,
    input  logic [riscv::VLEN-1:0]  lu_vaddr_i,
    output riscv::pte_t             lu_content_o,
    input  logic [ASID_WIDTH-1:0]   asid_to_be_flushed_i,
    input  logic [riscv::VLEN-1:0]  vaddr_to_be_flushed_i,
    output logic                    lu_is_2M_o,
    output logic                    lu_is_1G_o,
    output logic                    lu_hit_o
);
    
    struct packed {
      logic [ASID_WIDTH-1:0] asid;
      logic [riscv::VPN2:0]  vpn2;
      logic [8:0]            vpn1;
      logic [8:0]            vpn0;
      logic                  is_2M;
      logic                  is_1G;
      logic                  valid;
    } [TLB_ENTRIES-1:0] tags_q, tags_n;
    riscv::pte_t [TLB_ENTRIES-1:0] content_q, content_n;
    logic [8:0] vpn0, vpn1;
    logic [riscv::VPN2:0] vpn2;
    logic [TLB_ENTRIES-1:0] lu_hit;     
    logic [TLB_ENTRIES-1:0] replace_en; 
    
    
    
    always_comb begin : translation
        vpn0 = lu_vaddr_i[20:12];
        vpn1 = lu_vaddr_i[29:21];
        vpn2 = lu_vaddr_i[30+riscv::VPN2:30];
        
        lu_hit       = '{default: 0};
        lu_hit_o     = 1'b0;
        lu_content_o = '{default: 0};
        lu_is_1G_o   = 1'b0;
        lu_is_2M_o   = 1'b0;
        for (int unsigned i = 0; i < TLB_ENTRIES; i++) begin
            
            
            if (tags_q[i].valid && ((lu_asid_i == tags_q[i].asid) || content_q[i].g)  && vpn2 == tags_q[i].vpn2) begin
                
                if (tags_q[i].is_1G) begin
                    lu_is_1G_o = 1'b1;
                    lu_content_o = content_q[i];
                    lu_hit_o   = 1'b1;
                    lu_hit[i]  = 1'b1;
                
                end else if (vpn1 == tags_q[i].vpn1) begin
                    
                    
                    if (tags_q[i].is_2M || vpn0 == tags_q[i].vpn0) begin
                        lu_is_2M_o   = tags_q[i].is_2M;
                        lu_content_o = content_q[i];
                        lu_hit_o     = 1'b1;
                        lu_hit[i]    = 1'b1;
                    end
                end
            end
        end
    end
    logic asid_to_be_flushed_is0;  
    logic vaddr_to_be_flushed_is0;  
    logic  [TLB_ENTRIES-1:0] vaddr_vpn0_match;
    logic  [TLB_ENTRIES-1:0] vaddr_vpn1_match;
    logic  [TLB_ENTRIES-1:0] vaddr_vpn2_match;
    assign asid_to_be_flushed_is0 =  ~(|asid_to_be_flushed_i);
    assign vaddr_to_be_flushed_is0 = ~(|vaddr_to_be_flushed_i);
	  
    
    
    always_comb begin : update_flush
        tags_n    = tags_q;
        content_n = content_q;
        for (int unsigned i = 0; i < TLB_ENTRIES; i++) begin
            vaddr_vpn0_match[i] = (vaddr_to_be_flushed_i[20:12] == tags_q[i].vpn0);
            vaddr_vpn1_match[i] = (vaddr_to_be_flushed_i[29:21] == tags_q[i].vpn1);
            vaddr_vpn2_match[i] = (vaddr_to_be_flushed_i[30+riscv::VPN2:30] == tags_q[i].vpn2);
            if (flush_i) begin
                
                
        				if (asid_to_be_flushed_is0 && vaddr_to_be_flushed_is0 )
                    tags_n[i].valid = 1'b0;
                
                else if (asid_to_be_flushed_is0 && ((vaddr_vpn0_match[i] && vaddr_vpn1_match[i] && vaddr_vpn2_match[i]) || (vaddr_vpn2_match[i] && tags_q[i].is_1G) || (vaddr_vpn1_match[i] && vaddr_vpn2_match[i] && tags_q[i].is_2M) ) && (~vaddr_to_be_flushed_is0))
                    tags_n[i].valid = 1'b0;
                
                else if ((!content_q[i].g) && ((vaddr_vpn0_match[i] && vaddr_vpn1_match[i] && vaddr_vpn2_match[i]) || (vaddr_vpn2_match[i] && tags_q[i].is_1G) || (vaddr_vpn1_match[i] && vaddr_vpn2_match[i] && tags_q[i].is_2M)) && (asid_to_be_flushed_i == tags_q[i].asid) && (!vaddr_to_be_flushed_is0) && (!asid_to_be_flushed_is0))
				          	tags_n[i].valid = 1'b0;
                
				        else if ((!content_q[i].g) && (vaddr_to_be_flushed_is0) && (asid_to_be_flushed_i == tags_q[i].asid) && (!asid_to_be_flushed_is0))
				        	  tags_n[i].valid = 1'b0;
            
            end else if (update_i.valid & replace_en[i]) begin
                
                tags_n[i] = '{
                    asid:  update_i.asid,
                    vpn2:  update_i.vpn [18+riscv::VPN2:18],
                    vpn1:  update_i.vpn [17:9],
                    vpn0:  update_i.vpn [8:0],
                    is_1G: update_i.is_1G,
                    is_2M: update_i.is_2M,
                    valid: 1'b1
                };
                
                content_n[i] = update_i.content;
            end
        end
    end
    
    
    
    logic[2*(TLB_ENTRIES-1)-1:0] plru_tree_q, plru_tree_n;
    always_comb begin : plru_replacement
        plru_tree_n = plru_tree_q;
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        for (int unsigned i = 0; i < TLB_ENTRIES; i++) begin
            automatic int unsigned idx_base, shift, new_index;
            
            if (lu_hit[i] & lu_access_i) begin
                
                for (int unsigned lvl = 0; lvl < $clog2(TLB_ENTRIES); lvl++) begin
                  idx_base = $unsigned((2**lvl)-1);
                  
                  shift = $clog2(TLB_ENTRIES) - lvl;
                  
                  new_index =  ~((i >> (shift-1)) & 32'b1);
                  plru_tree_n[idx_base + (i >> shift)] = new_index[0];
                end
            end
        end
        
        
        
        
        
        
        
        
        
        
        
        
        
        
        for (int unsigned i = 0; i < TLB_ENTRIES; i += 1) begin
            automatic logic en;
            automatic int unsigned idx_base, shift, new_index;
            en = 1'b1;
            for (int unsigned lvl = 0; lvl < $clog2(TLB_ENTRIES); lvl++) begin
                idx_base = $unsigned((2**lvl)-1);
                
                shift = $clog2(TLB_ENTRIES) - lvl;
                
                new_index =  (i >> (shift-1)) & 32'b1;
                if (new_index[0]) begin
                  en &= plru_tree_q[idx_base + (i>>shift)];
                end else begin
                  en &= ~plru_tree_q[idx_base + (i>>shift)];
                end
            end
            replace_en[i] = en;
        end
    end
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if(~rst_ni) begin
            tags_q      <= '{default: 0};
            content_q   <= '{default: 0};
            plru_tree_q <= '{default: 0};
        end else begin
            tags_q      <= tags_n;
            content_q   <= content_n;
            plru_tree_q <= plru_tree_n;
        end
    end
    
    
    
    
    
    
    
endmodule
module ariane_regfile #(
  parameter int unsigned DATA_WIDTH     = 32,
  parameter int unsigned NR_READ_PORTS  = 2,
  parameter int unsigned NR_WRITE_PORTS = 2,
  parameter bit          ZERO_REG_ZERO  = 0
)(
  
  input  logic                                      clk_i,
  input  logic                                      rst_ni,
  
  input  logic                                      test_en_i,
  
  input  logic [NR_READ_PORTS-1:0][4:0]             raddr_i,
  output logic [NR_READ_PORTS-1:0][DATA_WIDTH-1:0]  rdata_o,
  
  input  logic [NR_WRITE_PORTS-1:0][4:0]            waddr_i,
  input  logic [NR_WRITE_PORTS-1:0][DATA_WIDTH-1:0] wdata_i,
  input  logic [NR_WRITE_PORTS-1:0]                 we_i
);
  localparam    ADDR_WIDTH = 5;
  localparam    NUM_WORDS  = 2**ADDR_WIDTH;
  logic [NUM_WORDS-1:0][DATA_WIDTH-1:0]     mem;
  logic [NR_WRITE_PORTS-1:0][NUM_WORDS-1:0] we_dec;
    always_comb begin : we_decoder
        for (int unsigned j = 0; j < NR_WRITE_PORTS; j++) begin
            for (int unsigned i = 0; i < NUM_WORDS; i++) begin
                if (waddr_i[j] == i)
                    we_dec[j][i] = we_i[j];
                else
                    we_dec[j][i] = 1'b0;
            end
        end
    end
    
    always_ff @(posedge clk_i, negedge rst_ni) begin : register_write_behavioral
        if (~rst_ni) begin
            mem <= '{default: '0};
        end else begin
            for (int unsigned j = 0; j < NR_WRITE_PORTS; j++) begin
                for (int unsigned i = 0; i < NUM_WORDS; i++) begin
                    if (we_dec[j][i]) begin
                        mem[i] <= wdata_i[j];
                    end
                end
                if (ZERO_REG_ZERO) begin
                  mem[0] <= '0;
                end
            end
        end
    end
  for (genvar i = 0; i < NR_READ_PORTS; i++) begin
    assign rdata_o[i] = mem[raddr_i[i]];
  end
endmodule
module re_name import ariane_pkg::*; (
    input  logic                                   clk_i,    
    input  logic                                   rst_ni,   
    input  logic                                   flush_i,  
    input  logic                                   flush_unissied_instr_i,
    
    input  scoreboard_entry_t                      issue_instr_i,
    input  logic                                   issue_instr_valid_i,
    output logic                                   issue_ack_o,
    
    output scoreboard_entry_t                      issue_instr_o,
    output logic                                   issue_instr_valid_o,
    input  logic                                   issue_ack_i
);
    
    assign issue_instr_valid_o = issue_instr_valid_i;
    assign issue_ack_o         = issue_ack_i;
    
    logic [31:0] re_name_table_gpr_n, re_name_table_gpr_q;
    logic [31:0] re_name_table_fpr_n, re_name_table_fpr_q;
    
    
    
    always_comb begin
        
        logic name_bit_rs1, name_bit_rs2, name_bit_rs3, name_bit_rd;
        
        re_name_table_gpr_n = re_name_table_gpr_q;
        re_name_table_fpr_n = re_name_table_fpr_q;
        issue_instr_o       = issue_instr_i;
        if (issue_ack_i && !flush_unissied_instr_i) begin
            
            if (is_rd_fpr(issue_instr_i.op))
                re_name_table_fpr_n[issue_instr_i.rd] = re_name_table_fpr_q[issue_instr_i.rd] ^ 1'b1;
            else
                re_name_table_gpr_n[issue_instr_i.rd] = re_name_table_gpr_q[issue_instr_i.rd] ^ 1'b1;
        end
        
        name_bit_rs1 = is_rs1_fpr(issue_instr_i.op) ? re_name_table_fpr_q[issue_instr_i.rs1]
                                                    : re_name_table_gpr_q[issue_instr_i.rs1];
        name_bit_rs2 = is_rs2_fpr(issue_instr_i.op) ? re_name_table_fpr_q[issue_instr_i.rs2]
                                                    : re_name_table_gpr_q[issue_instr_i.rs2];
        
        name_bit_rs3 = re_name_table_fpr_q[issue_instr_i.result[4:0]]; 
        
        name_bit_rd = is_rd_fpr(issue_instr_i.op) ? re_name_table_fpr_q[issue_instr_i.rd] ^ 1'b1
                                                  : re_name_table_gpr_q[issue_instr_i.rd] ^ (issue_instr_i.rd != '0); 
        
        issue_instr_o.rs1 = { ENABLE_RENAME & name_bit_rs1, issue_instr_i.rs1[4:0] };
        issue_instr_o.rs2 = { ENABLE_RENAME & name_bit_rs2, issue_instr_i.rs2[4:0] };
        
        if (is_imm_fpr(issue_instr_i.op))
            issue_instr_o.result = { ENABLE_RENAME & name_bit_rs3, issue_instr_i.result[4:0]};
        
        issue_instr_o.rd = { ENABLE_RENAME & name_bit_rd, issue_instr_i.rd[4:0] };
        
        re_name_table_gpr_n[0] = 1'b0;
        
        if (flush_i) begin
            re_name_table_gpr_n = '0;
            re_name_table_fpr_n = '0;
        end
    end
    
    
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (~rst_ni) begin
            re_name_table_gpr_q <= '0;
            re_name_table_fpr_q <= '0;
        end else begin
            re_name_table_gpr_q <= re_name_table_gpr_n;
            re_name_table_fpr_q <= re_name_table_fpr_n;
        end
    end
endmodule
module scoreboard #(
  parameter int unsigned NR_ENTRIES      = 8, 
  parameter int unsigned NR_WB_PORTS     = 1,
  parameter int unsigned NR_COMMIT_PORTS = 2
) (
  input  logic                                                  clk_i,    
  input  logic                                                  rst_ni,   
  output logic                                                  sb_full_o,
  input  logic                                                  flush_unissued_instr_i, 
  input  logic                                                  flush_i,  
  input  logic                                                  unresolved_branch_i, 
  
  output ariane_pkg::fu_t [2**ariane_pkg::REG_ADDR_SIZE-1:0]    rd_clobber_gpr_o,
  output ariane_pkg::fu_t [2**ariane_pkg::REG_ADDR_SIZE-1:0]    rd_clobber_fpr_o,
  
  input  logic [ariane_pkg::REG_ADDR_SIZE-1:0]                  rs1_i,
  output riscv::xlen_t                                          rs1_o,
  output logic                                                  rs1_valid_o,
  input  logic [ariane_pkg::REG_ADDR_SIZE-1:0]                  rs2_i,
  output riscv::xlen_t                                          rs2_o,
  output logic                                                  rs2_valid_o,
  input  logic [ariane_pkg::REG_ADDR_SIZE-1:0]                  rs3_i,
  output logic [ariane_pkg::FLEN-1:0]                           rs3_o,
  output logic                                                  rs3_valid_o,
  
  output ariane_pkg::scoreboard_entry_t [NR_COMMIT_PORTS-1:0]   commit_instr_o,
  input  logic              [NR_COMMIT_PORTS-1:0]               commit_ack_i,
  
  
  input  ariane_pkg::scoreboard_entry_t                         decoded_instr_i,
  input  logic                                                  decoded_instr_valid_i,
  output logic                                                  decoded_instr_ack_o,
  
  output ariane_pkg::scoreboard_entry_t                         issue_instr_o,
  output logic                                                  issue_instr_valid_o,
  input  logic                                                  issue_ack_i,
  
  input ariane_pkg::bp_resolve_t                                resolved_branch_i,
  input logic [NR_WB_PORTS-1:0][ariane_pkg::TRANS_ID_BITS-1:0]  trans_id_i,  
  input logic [NR_WB_PORTS-1:0][riscv::XLEN-1:0]                wbdata_i,    
  input ariane_pkg::exception_t [NR_WB_PORTS-1:0]               ex_i,        
  input logic [NR_WB_PORTS-1:0]                                 wt_valid_i   
);
  localparam int unsigned BITS_ENTRIES = $clog2(NR_ENTRIES);
  
  typedef struct packed {
    logic                          issued;         
    logic                          is_rd_fpr_flag; 
    ariane_pkg::scoreboard_entry_t sbe;            
  } sb_mem_t;
  sb_mem_t [NR_ENTRIES-1:0] mem_q, mem_n;
  logic                    issue_full, issue_en;
  logic [BITS_ENTRIES-1:0] issue_cnt_n,      issue_cnt_q;
  logic [BITS_ENTRIES-1:0] issue_pointer_n,  issue_pointer_q;
  logic [NR_COMMIT_PORTS-1:0][BITS_ENTRIES-1:0] commit_pointer_n, commit_pointer_q;
  logic [$clog2(NR_COMMIT_PORTS):0] num_commit;
  
  
  assign issue_full = &issue_cnt_q;
  assign sb_full_o = issue_full;
  
  always_comb begin : commit_ports
    for (int unsigned i = 0; i < NR_COMMIT_PORTS; i++) begin
      commit_instr_o[i] = mem_q[commit_pointer_q[i]].sbe;
      commit_instr_o[i].trans_id = commit_pointer_q[i];
    end
  end
  
  always_comb begin
    issue_instr_o          = decoded_instr_i;
    
    issue_instr_o.trans_id = issue_pointer_q;
    
    
    issue_instr_valid_o    = decoded_instr_valid_i & ~unresolved_branch_i & ~issue_full;
    decoded_instr_ack_o    = issue_ack_i & ~issue_full;
  end
  
  
  always_comb begin : issue_fifo
    
    mem_n          = mem_q;
    issue_en       = 1'b0;
    
    if (decoded_instr_valid_i && decoded_instr_ack_o && !flush_unissued_instr_i) begin
      
      
      issue_en = 1'b1;
      mem_n[issue_pointer_q] = {1'b1,                                      
                                ariane_pkg::is_rd_fpr(decoded_instr_i.op), 
                                decoded_instr_i                            
                                };
    end
    
    
    
    for (int unsigned i = 0; i < NR_ENTRIES; i++) begin
      
      if (mem_q[i].sbe.fu == ariane_pkg::NONE && mem_q[i].issued)
        mem_n[i].sbe.valid = 1'b1;
    end
    
    
    
    for (int unsigned i = 0; i < NR_WB_PORTS; i++) begin
      
      
      if (wt_valid_i[i] && mem_q[trans_id_i[i]].issued) begin
        mem_n[trans_id_i[i]].sbe.valid  = 1'b1;
        mem_n[trans_id_i[i]].sbe.result = wbdata_i[i];
        
        mem_n[trans_id_i[i]].sbe.bp.predict_address = resolved_branch_i.target_address;
        
        if (ex_i[i].valid)
          mem_n[trans_id_i[i]].sbe.ex = ex_i[i];
        
        else if (mem_q[trans_id_i[i]].sbe.fu inside {ariane_pkg::FPU, ariane_pkg::FPU_VEC})
          mem_n[trans_id_i[i]].sbe.ex.cause = ex_i[i].cause;
      end
    end
    
    
    
    
    for (logic [BITS_ENTRIES-1:0] i = 0; i < NR_COMMIT_PORTS; i++) begin
      if (commit_ack_i[i]) begin
        
        mem_n[commit_pointer_q[i]].issued     = 1'b0;
        mem_n[commit_pointer_q[i]].sbe.valid  = 1'b0;
      end
    end
    
    
    
    if (flush_i) begin
      for (int unsigned i = 0; i < NR_ENTRIES; i++) begin
        
        mem_n[i].issued       = 1'b0;
        mem_n[i].sbe.valid    = 1'b0;
        mem_n[i].sbe.ex.valid = 1'b0;
      end
    end
  end
  
  popcount #(
    .INPUT_WIDTH(NR_COMMIT_PORTS)
  ) i_popcount (
    .data_i(commit_ack_i),
    .popcount_o(num_commit)
  );
  assign issue_cnt_n         = (flush_i) ? '0 : issue_cnt_q         - num_commit + issue_en;
  assign commit_pointer_n[0] = (flush_i) ? '0 : commit_pointer_q[0] + num_commit;
  assign issue_pointer_n     = (flush_i) ? '0 : issue_pointer_q     + issue_en;
  
  for (genvar k=1; k < NR_COMMIT_PORTS; k++) begin : gen_cnt_incr
    assign commit_pointer_n[k] = (flush_i) ? '0 : commit_pointer_n[0] + unsigned'(k);
  end
  
  
  
  
  logic [2**ariane_pkg::REG_ADDR_SIZE-1:0][NR_ENTRIES:0]              gpr_clobber_vld;
  logic [2**ariane_pkg::REG_ADDR_SIZE-1:0][NR_ENTRIES:0]              fpr_clobber_vld;
  ariane_pkg::fu_t [NR_ENTRIES:0]                                     clobber_fu;
  always_comb begin : clobber_assign
    gpr_clobber_vld  = '0;
    fpr_clobber_vld  = '0;
    
    clobber_fu[NR_ENTRIES] = ariane_pkg::NONE;
    for (int unsigned i = 0; i < 2**ariane_pkg::REG_ADDR_SIZE; i++) begin
      gpr_clobber_vld[i][NR_ENTRIES] = 1'b1;
      fpr_clobber_vld[i][NR_ENTRIES] = 1'b1;
    end
    
    for (int unsigned i = 0; i < NR_ENTRIES; i++) begin
      gpr_clobber_vld[mem_q[i].sbe.rd][i] = mem_q[i].issued & ~mem_q[i].is_rd_fpr_flag;
      fpr_clobber_vld[mem_q[i].sbe.rd][i] = mem_q[i].issued & mem_q[i].is_rd_fpr_flag;
      clobber_fu[i]                       = mem_q[i].sbe.fu;
    end
    
    gpr_clobber_vld[0] = '0;
  end
  for (genvar k = 0; k < 2**ariane_pkg::REG_ADDR_SIZE; k++) begin : gen_sel_clobbers
    
    rr_arb_tree #(
      .NumIn(NR_ENTRIES+1),
      .DataType(ariane_pkg::fu_t),
      .ExtPrio(1'b1),
      .AxiVldRdy(1'b1)
    ) i_sel_gpr_clobbers (
      .clk_i   ( clk_i               ),
      .rst_ni  ( rst_ni              ),
      .flush_i ( 1'b0                ),
      .rr_i    ( '0                  ),
      .req_i   ( gpr_clobber_vld[k]  ),
      .gnt_o   (                     ),
      .data_i  ( clobber_fu          ),
      .gnt_i   ( 1'b1                ),
      .req_o   (                     ),
      .data_o  ( rd_clobber_gpr_o[k] ),
      .idx_o   (                     )
    );
    rr_arb_tree #(
      .NumIn(NR_ENTRIES+1),
      .DataType(ariane_pkg::fu_t),
      .ExtPrio(1'b1),
      .AxiVldRdy(1'b1)
    ) i_sel_fpr_clobbers (
      .clk_i   ( clk_i               ),
      .rst_ni  ( rst_ni              ),
      .flush_i ( 1'b0                ),
      .rr_i    ( '0                  ),
      .req_i   ( fpr_clobber_vld[k]  ),
      .gnt_o   (                     ),
      .data_i  ( clobber_fu          ),
      .gnt_i   ( 1'b1                ),
      .req_o   (                     ),
      .data_o  ( rd_clobber_fpr_o[k] ),
      .idx_o   (                     )
    );
  end
  
  
  
  
  logic [NR_ENTRIES+NR_WB_PORTS-1:0] rs1_fwd_req, rs2_fwd_req, rs3_fwd_req;
  logic [NR_ENTRIES+NR_WB_PORTS-1:0][riscv::XLEN-1:0] rs_data;
  logic rs1_valid, rs2_valid;
  
  for (genvar k = 0; unsigned'(k) < NR_WB_PORTS; k++) begin : gen_rs_wb
    assign rs1_fwd_req[k] = (mem_q[trans_id_i[k]].sbe.rd == rs1_i) & wt_valid_i[k] & (~ex_i[k].valid) & (mem_q[trans_id_i[k]].is_rd_fpr_flag == ariane_pkg::is_rs1_fpr(issue_instr_o.op));
    assign rs2_fwd_req[k] = (mem_q[trans_id_i[k]].sbe.rd == rs2_i) & wt_valid_i[k] & (~ex_i[k].valid) & (mem_q[trans_id_i[k]].is_rd_fpr_flag == ariane_pkg::is_rs2_fpr(issue_instr_o.op));
    assign rs3_fwd_req[k] = (mem_q[trans_id_i[k]].sbe.rd == rs3_i) & wt_valid_i[k] & (~ex_i[k].valid) & (mem_q[trans_id_i[k]].is_rd_fpr_flag == ariane_pkg::is_imm_fpr(issue_instr_o.op));
    assign rs_data[k]     = wbdata_i[k];
  end
  for (genvar k = 0; unsigned'(k) < NR_ENTRIES; k++) begin : gen_rs_entries
    assign rs1_fwd_req[k+NR_WB_PORTS] = (mem_q[k].sbe.rd == rs1_i) & mem_q[k].issued & mem_q[k].sbe.valid & (mem_q[k].is_rd_fpr_flag == ariane_pkg::is_rs1_fpr(issue_instr_o.op));
    assign rs2_fwd_req[k+NR_WB_PORTS] = (mem_q[k].sbe.rd == rs2_i) & mem_q[k].issued & mem_q[k].sbe.valid & (mem_q[k].is_rd_fpr_flag == ariane_pkg::is_rs2_fpr(issue_instr_o.op));
    assign rs3_fwd_req[k+NR_WB_PORTS] = (mem_q[k].sbe.rd == rs3_i) & mem_q[k].issued & mem_q[k].sbe.valid & (mem_q[k].is_rd_fpr_flag == ariane_pkg::is_imm_fpr(issue_instr_o.op));
    assign rs_data[k+NR_WB_PORTS]     = mem_q[k].sbe.result;
  end
  
  assign rs1_valid_o = rs1_valid & ((|rs1_i) | ariane_pkg::is_rs1_fpr(issue_instr_o.op));
  assign rs2_valid_o = rs2_valid & ((|rs2_i) | ariane_pkg::is_rs2_fpr(issue_instr_o.op));
  
  
  rr_arb_tree #(
    .NumIn(NR_ENTRIES+NR_WB_PORTS),
    .DataWidth(riscv::XLEN),
    .ExtPrio(1'b1),
    .AxiVldRdy(1'b1)
  ) i_sel_rs1 (
    .clk_i   ( clk_i       ),
    .rst_ni  ( rst_ni      ),
    .flush_i ( 1'b0        ),
    .rr_i    ( '0          ),
    .req_i   ( rs1_fwd_req ),
    .gnt_o   (             ),
    .data_i  ( rs_data     ),
    .gnt_i   ( 1'b1        ),
    .req_o   ( rs1_valid   ),
    .data_o  ( rs1_o       ),
    .idx_o   (             )
  );
  rr_arb_tree #(
    .NumIn(NR_ENTRIES+NR_WB_PORTS),
    .DataWidth(riscv::XLEN),
    .ExtPrio(1'b1),
    .AxiVldRdy(1'b1)
  ) i_sel_rs2 (
    .clk_i   ( clk_i       ),
    .rst_ni  ( rst_ni      ),
    .flush_i ( 1'b0        ),
    .rr_i    ( '0          ),
    .req_i   ( rs2_fwd_req ),
    .gnt_o   (             ),
    .data_i  ( rs_data     ),
    .gnt_i   ( 1'b1        ),
    .req_o   ( rs2_valid   ),
    .data_o  ( rs2_o       ),
    .idx_o   (             )
  );
  riscv::xlen_t           rs3;
  rr_arb_tree #(
    .NumIn(NR_ENTRIES+NR_WB_PORTS),
    .DataWidth(riscv::XLEN),
    .ExtPrio(1'b1),
    .AxiVldRdy(1'b1)
  ) i_sel_rs3 (
    .clk_i   ( clk_i       ),
    .rst_ni  ( rst_ni      ),
    .flush_i ( 1'b0        ),
    .rr_i    ( '0          ),
    .req_i   ( rs3_fwd_req ),
    .gnt_o   (             ),
    .data_i  ( rs_data     ),
    .gnt_i   ( 1'b1        ),
    .req_o   ( rs3_valid_o ),
    .data_o  ( rs3         ),
    .idx_o   (             )
  );
  assign rs3_o = rs3[ariane_pkg::FLEN-1:0];
  
  always_ff @(posedge clk_i or negedge rst_ni) begin : regs
    if(!rst_ni) begin
      mem_q                 <= '{default: sb_mem_t'(0)};
      issue_cnt_q           <= '0;
      commit_pointer_q      <= '0;
      issue_pointer_q       <= '0;
    end else begin
      issue_cnt_q           <= issue_cnt_n;
      issue_pointer_q       <= issue_pointer_n;
      mem_q                 <= mem_n;
      commit_pointer_q      <= commit_pointer_n;
    end
  end
  
  
  
  
endmodule
module store_buffer import ariane_pkg::*; (
    input logic          clk_i,           
    input logic          rst_ni,          
    input logic          flush_i,         
                                          
    output logic         no_st_pending_o, 
    output logic         store_buffer_empty_o, 
    input  logic [11:0]  page_offset_i,         
    output logic         page_offset_matches_o, 
    input  logic         commit_i,        
    output logic         commit_ready_o,  
    output logic         ready_o,         
                                          
                                          
    input  logic         valid_i,         
    input  logic         valid_without_flush_i, 
    input  logic [riscv::PLEN-1:0]  paddr_i,         
    input  riscv::xlen_t            data_i,          
    input  logic [7:0]   be_i,            
    input  logic [1:0]   data_size_i,     
    
    input  dcache_req_o_t req_port_i,
    output dcache_req_i_t req_port_o
);
    
    
    
    struct packed {
        logic [riscv::PLEN-1:0] address;
        riscv::xlen_t           data;
        logic [7:0]             be;
        logic [1:0]             data_size;
        logic                   valid;     
    } speculative_queue_n [DEPTH_SPEC-1:0], speculative_queue_q [DEPTH_SPEC-1:0],
      commit_queue_n [DEPTH_COMMIT-1:0],    commit_queue_q [DEPTH_COMMIT-1:0];
    
    logic [$clog2(DEPTH_SPEC):0] speculative_status_cnt_n, speculative_status_cnt_q;
    logic [$clog2(DEPTH_COMMIT):0] commit_status_cnt_n, commit_status_cnt_q;
    
    logic [$clog2(DEPTH_SPEC)-1:0] speculative_read_pointer_n,  speculative_read_pointer_q;
    logic [$clog2(DEPTH_SPEC)-1:0] speculative_write_pointer_n, speculative_write_pointer_q;
    
    logic [$clog2(DEPTH_COMMIT)-1:0] commit_read_pointer_n,  commit_read_pointer_q;
    logic [$clog2(DEPTH_COMMIT)-1:0] commit_write_pointer_n, commit_write_pointer_q;
    assign store_buffer_empty_o = (speculative_status_cnt_q == 0) & no_st_pending_o;
    
    
    
    always_comb begin : core_if
        automatic logic [DEPTH_SPEC:0] speculative_status_cnt;
        speculative_status_cnt = speculative_status_cnt_q;
        
        ready_o = (speculative_status_cnt_q < (DEPTH_SPEC - 1)) || commit_i;
        
        speculative_status_cnt_n    = speculative_status_cnt_q;
        speculative_read_pointer_n  = speculative_read_pointer_q;
        speculative_write_pointer_n = speculative_write_pointer_q;
        speculative_queue_n         = speculative_queue_q;
        
        
        if (valid_i) begin
            speculative_queue_n[speculative_write_pointer_q].address   = paddr_i;
            speculative_queue_n[speculative_write_pointer_q].data      = data_i;
            speculative_queue_n[speculative_write_pointer_q].be        = be_i;
            speculative_queue_n[speculative_write_pointer_q].data_size = data_size_i;
            speculative_queue_n[speculative_write_pointer_q].valid   = 1'b1;
            
            speculative_write_pointer_n = speculative_write_pointer_q + 1'b1;
            speculative_status_cnt++;
        end
        
        
        if (commit_i) begin
            
            speculative_queue_n[speculative_read_pointer_q].valid = 1'b0;
            
            speculative_read_pointer_n = speculative_read_pointer_q + 1'b1;
            speculative_status_cnt--;
        end
        speculative_status_cnt_n = speculative_status_cnt;
        
        if (flush_i) begin
            
            for (int unsigned i = 0; i < DEPTH_SPEC; i++)
                speculative_queue_n[i].valid = 1'b0;
            speculative_write_pointer_n = speculative_read_pointer_q;
            
            speculative_status_cnt_n = 'b0;
        end
    end
    
    
    
    
    
    assign req_port_o.kill_req  = 1'b0;
    assign req_port_o.data_we   = 1'b1; 
    assign req_port_o.tag_valid = 1'b0;
    
    assign req_port_o.address_index = commit_queue_q[commit_read_pointer_q].address[ariane_pkg::DCACHE_INDEX_WIDTH-1:0];
    
    assign req_port_o.address_tag   = commit_queue_q[commit_read_pointer_q].address[ariane_pkg::DCACHE_TAG_WIDTH     +
                                                                                    ariane_pkg::DCACHE_INDEX_WIDTH-1 :
                                                                                    ariane_pkg::DCACHE_INDEX_WIDTH];
    assign req_port_o.data_wdata    = (req_port_o.address_index[2] == 1'b0) ? {{64-riscv::XLEN{1'b0}}, commit_queue_q[commit_read_pointer_q].data} :
                                                                              {commit_queue_q[commit_read_pointer_q].data, {64-riscv::XLEN{1'b0}}};
    assign req_port_o.data_be       = commit_queue_q[commit_read_pointer_q].be;
    assign req_port_o.data_size     = commit_queue_q[commit_read_pointer_q].data_size;
    always_comb begin : store_if
        automatic logic [DEPTH_COMMIT:0] commit_status_cnt;
        commit_status_cnt = commit_status_cnt_q;
        commit_ready_o = (commit_status_cnt_q < DEPTH_COMMIT);
        
        no_st_pending_o         = (commit_status_cnt_q == 0);
        
        commit_read_pointer_n   = commit_read_pointer_q;
        commit_write_pointer_n  = commit_write_pointer_q;
        commit_queue_n = commit_queue_q;
        req_port_o.data_req     = 1'b0;
        
        
        if (commit_queue_q[commit_read_pointer_q].valid) begin
            req_port_o.data_req = 1'b1;
            if (req_port_i.data_gnt) begin
                
                commit_queue_n[commit_read_pointer_q].valid = 1'b0;
                
                commit_read_pointer_n = commit_read_pointer_q + 1'b1;
                commit_status_cnt--;
            end
        end
        
        
        
        if (commit_i) begin
            commit_queue_n[commit_write_pointer_q] = speculative_queue_q[speculative_read_pointer_q];
            commit_write_pointer_n = commit_write_pointer_n + 1'b1;
            commit_status_cnt++;
        end
        commit_status_cnt_n     = commit_status_cnt;
    end
    
    
    
    
    
    
    
    
    
    
    
    
    
    
    always_comb begin : address_checker
        page_offset_matches_o = 1'b0;
        
        for (int unsigned i = 0; i < DEPTH_COMMIT; i++) begin
            
            if ((page_offset_i[11:3] == commit_queue_q[i].address[11:3]) && commit_queue_q[i].valid) begin
                page_offset_matches_o = 1'b1;
                break;
            end
        end
        for (int unsigned i = 0; i < DEPTH_SPEC; i++) begin
            
            if ((page_offset_i[11:3] == speculative_queue_q[i].address[11:3]) && speculative_queue_q[i].valid) begin
                page_offset_matches_o = 1'b1;
                break;
            end
        end
        
        if ((page_offset_i[11:3] == paddr_i[11:3]) && valid_without_flush_i) begin
            page_offset_matches_o = 1'b1;
        end
    end
    
    always_ff @(posedge clk_i or negedge rst_ni) begin : p_spec
        if (~rst_ni) begin
            speculative_queue_q         <= '{default: 0};
            speculative_read_pointer_q  <= '0;
            speculative_write_pointer_q <= '0;
            speculative_status_cnt_q    <= '0;
        end else begin
            speculative_queue_q         <= speculative_queue_n;
            speculative_read_pointer_q  <= speculative_read_pointer_n;
            speculative_write_pointer_q <= speculative_write_pointer_n;
            speculative_status_cnt_q    <= speculative_status_cnt_n;
        end
     end
    
    always_ff @(posedge clk_i or negedge rst_ni) begin : p_commit
        if (~rst_ni) begin
            commit_queue_q              <= '{default: 0};
            commit_read_pointer_q       <= '0;
            commit_write_pointer_q      <= '0;
            commit_status_cnt_q         <= '0;
        end else begin
            commit_queue_q              <= commit_queue_n;
            commit_read_pointer_q       <= commit_read_pointer_n;
            commit_write_pointer_q      <= commit_write_pointer_n;
            commit_status_cnt_q         <= commit_status_cnt_n;
        end
     end
    
    
    
    
endmodule
module amo_buffer (
    input  logic clk_i,              
    input  logic rst_ni,             
    input  logic flush_i,            
    input  logic             valid_i,            
    output logic             ready_o,            
    input  ariane_pkg::amo_t amo_op_i,           
    input  logic [riscv::PLEN-1:0]      paddr_i,            
    input  riscv::xlen_t     data_i,             
    input  logic [1:0]       data_size_i,        
    
    output ariane_pkg::amo_req_t  amo_req_o,          
    input  ariane_pkg::amo_resp_t amo_resp_i,         
    
    input  logic amo_valid_commit_i, 
    input  logic no_st_pending_i     
);
    logic flush_amo_buffer;
    logic amo_valid;
    typedef struct packed {
        ariane_pkg::amo_t        op;
        logic [riscv::PLEN-1:0] paddr;
        riscv::xlen_t data;
        logic [1:0]  size;
    } amo_op_t ;
    amo_op_t amo_data_in, amo_data_out;
    
    assign amo_req_o.req = no_st_pending_i & amo_valid_commit_i & amo_valid;
    assign amo_req_o.amo_op = amo_data_out.op;
    assign amo_req_o.size = amo_data_out.size;
    assign amo_req_o.operand_a = {{64-riscv::PLEN{1'b0}}, amo_data_out.paddr};
    assign amo_req_o.operand_b = {{64-riscv::XLEN{1'b0}}, amo_data_out.data};
    assign amo_data_in.op = amo_op_i;
    assign amo_data_in.data = data_i;
    assign amo_data_in.paddr = paddr_i;
    assign amo_data_in.size = data_size_i;
    
    
    assign flush_amo_buffer = flush_i & !amo_valid_commit_i;
    fifo_v3 #(
        .DEPTH        ( 1                ),
        .dtype        ( amo_op_t         )
    ) i_amo_fifo (
        .clk_i        ( clk_i            ),
        .rst_ni       ( rst_ni           ),
        .flush_i      ( flush_amo_buffer ),
        .testmode_i   ( 1'b0             ),
        .full_o       ( amo_valid        ),
        .empty_o      ( ready_o          ),
        .usage_o      (  ), 
        .data_i       ( amo_data_in      ),
        .push_i       ( valid_i          ),
        .data_o       ( amo_data_out     ),
        .pop_i        ( amo_resp_i.ack   )
    );
endmodule
module store_unit import ariane_pkg::*; (
    input  logic                     clk_i,    
    input  logic                     rst_ni,  
    input  logic                     flush_i,
    output logic                     no_st_pending_o,
    output logic                     store_buffer_empty_o,
    
    input  logic                     valid_i,
    input  lsu_ctrl_t                lsu_ctrl_i,
    output logic                     pop_st_o,
    input  logic                     commit_i,
    output logic                     commit_ready_o,
    input  logic                     amo_valid_commit_i,
    
    output logic                     valid_o,
    output logic [TRANS_ID_BITS-1:0] trans_id_o,
    output riscv::xlen_t             result_o,
    output exception_t               ex_o,
    
    output logic                     translation_req_o, 
    output logic [riscv::VLEN-1:0]   vaddr_o,           
    input  logic [riscv::PLEN-1:0]   paddr_i,           
    input  exception_t               ex_i,
    input  logic                     dtlb_hit_i,       
    
    input  logic [11:0]              page_offset_i,
    output logic                     page_offset_matches_o,
    
    output amo_req_t                 amo_req_o,
    input  amo_resp_t                amo_resp_i,
    input  dcache_req_o_t            req_port_i,
    output dcache_req_i_t            req_port_o
);
    
    assign result_o = '0;
    enum logic [1:0] {
        IDLE,
        VALID_STORE,
        WAIT_TRANSLATION,
        WAIT_STORE_READY
    } state_d, state_q;
    
    logic st_ready;
    logic st_valid;
    logic st_valid_without_flush;
    logic instr_is_amo;
    assign instr_is_amo = is_amo(lsu_ctrl_i.operator);
    
    riscv::xlen_t st_data_n, st_data_q;
    logic [7:0]   st_be_n,        st_be_q;
    logic [1:0]   st_data_size_n, st_data_size_q;
    amo_t         amo_op_d,       amo_op_q;
    logic [TRANS_ID_BITS-1:0] trans_id_n, trans_id_q;
    
    assign vaddr_o    = lsu_ctrl_i.vaddr; 
    assign trans_id_o = trans_id_q; 
    always_comb begin : store_control
        translation_req_o      = 1'b0;
        valid_o                = 1'b0;
        st_valid               = 1'b0;
        st_valid_without_flush = 1'b0;
        pop_st_o               = 1'b0;
        ex_o                   = ex_i;
        trans_id_n             = lsu_ctrl_i.trans_id;
        state_d                     = state_q;
        case (state_q)
            
            IDLE: begin
                if (valid_i) begin
                    state_d = VALID_STORE;
                    translation_req_o = 1'b1;
                    pop_st_o = 1'b1;
                    
                    
                    if (!dtlb_hit_i) begin
                        state_d = WAIT_TRANSLATION;
                        pop_st_o = 1'b0;
                    end
                    if (!st_ready) begin
                        state_d = WAIT_STORE_READY;
                        pop_st_o = 1'b0;
                    end
                end
            end
            VALID_STORE: begin
                valid_o  = 1'b1;
                
                if (!flush_i)
                    st_valid = 1'b1;
                st_valid_without_flush = 1'b1;
                
                if (valid_i && !instr_is_amo) begin
                    translation_req_o = 1'b1;
                    state_d = VALID_STORE;
                    pop_st_o = 1'b1;
                    if (!dtlb_hit_i) begin
                        state_d = WAIT_TRANSLATION;
                        pop_st_o = 1'b0;
                    end
                    if (!st_ready) begin
                        state_d = WAIT_STORE_READY;
                        pop_st_o = 1'b0;
                    end
                
                end else begin
                    state_d = IDLE;
                end
            end
            
            WAIT_STORE_READY: begin
                
                translation_req_o = 1'b1;
                if (st_ready && dtlb_hit_i) begin
                    state_d = IDLE;
                end
            end
            
            
            
            WAIT_TRANSLATION: begin
                translation_req_o = 1'b1;
                if (dtlb_hit_i) begin
                    state_d = IDLE;
                end
            end
        endcase
        
        
        
        
        if (ex_i.valid && (state_q != IDLE)) begin
            
            pop_st_o = 1'b1;
            st_valid = 1'b0;
            state_d  = IDLE;
            valid_o  = 1'b1;
        end
        if (flush_i)
            state_d = IDLE;
    end
    
    
    
    
    always_comb begin
        st_be_n   = lsu_ctrl_i.be;
        
        st_data_n = instr_is_amo ? lsu_ctrl_i.data[riscv::XLEN-1:0]
                                 : data_align(lsu_ctrl_i.vaddr[2:0], {{64-riscv::XLEN{1'b0}}, lsu_ctrl_i.data[riscv::XLEN-1:0]});
        st_data_size_n = extract_transfer_size(lsu_ctrl_i.operator);
        
        case (lsu_ctrl_i.operator)
            AMO_LRW, AMO_LRD:     amo_op_d = AMO_LR;
            AMO_SCW, AMO_SCD:     amo_op_d = AMO_SC;
            AMO_SWAPW, AMO_SWAPD: amo_op_d = AMO_SWAP;
            AMO_ADDW, AMO_ADDD:   amo_op_d = AMO_ADD;
            AMO_ANDW, AMO_ANDD:   amo_op_d = AMO_AND;
            AMO_ORW, AMO_ORD:     amo_op_d = AMO_OR;
            AMO_XORW, AMO_XORD:   amo_op_d = AMO_XOR;
            AMO_MAXW, AMO_MAXD:   amo_op_d = AMO_MAX;
            AMO_MAXWU, AMO_MAXDU: amo_op_d = AMO_MAXU;
            AMO_MINW, AMO_MIND:   amo_op_d = AMO_MIN;
            AMO_MINWU, AMO_MINDU: amo_op_d = AMO_MINU;
            default: amo_op_d = AMO_NONE;
        endcase
    end
    logic store_buffer_valid, amo_buffer_valid;
    logic store_buffer_ready, amo_buffer_ready;
    
    assign store_buffer_valid = st_valid & (amo_op_q == AMO_NONE);
    assign amo_buffer_valid = st_valid & (amo_op_q != AMO_NONE);
    assign st_ready = store_buffer_ready & amo_buffer_ready;
    
    
    
    store_buffer store_buffer_i (
        .clk_i,
        .rst_ni,
        .flush_i,
        .no_st_pending_o,
        .store_buffer_empty_o,
        .page_offset_i,
        .page_offset_matches_o,
        .commit_i,
        .commit_ready_o,
        .ready_o               ( store_buffer_ready     ),
        .valid_i               ( store_buffer_valid     ),
        
        
        
        
        
        .valid_without_flush_i ( st_valid_without_flush ),
        .paddr_i,
        .data_i                ( st_data_q              ),
        .be_i                  ( st_be_q                ),
        .data_size_i           ( st_data_size_q         ),
        .req_port_i            ( req_port_i             ),
        .req_port_o            ( req_port_o             )
    );
    amo_buffer i_amo_buffer (
        .clk_i,
        .rst_ni,
        .flush_i,
        .valid_i            ( amo_buffer_valid   ),
        .ready_o            ( amo_buffer_ready   ),
        .paddr_i            ( paddr_i            ),
        .amo_op_i           ( amo_op_q           ),
        .data_i             ( st_data_q          ),
        .data_size_i        ( st_data_size_q     ),
        .amo_req_o          ( amo_req_o          ),
        .amo_resp_i         ( amo_resp_i         ),
        .amo_valid_commit_i ( amo_valid_commit_i ),
        .no_st_pending_i    ( no_st_pending_o    )
    );
    
    
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (~rst_ni) begin
            state_q             <= IDLE;
            st_be_q        <= '0;
            st_data_q      <= '0;
            st_data_size_q <= '0;
            trans_id_q     <= '0;
            amo_op_q       <= AMO_NONE;
        end else begin
            state_q        <= state_d;
            st_be_q        <= st_be_n;
            st_data_q      <= st_data_n;
            trans_id_q     <= trans_id_n;
            st_data_size_q <= st_data_size_n;
            amo_op_q       <= amo_op_d;
        end
    end
endmodule
module commit_stage import ariane_pkg::*; #(
    parameter int unsigned NR_COMMIT_PORTS = 2
)(
    input  logic                                    clk_i,
    input  logic                                    rst_ni,
    input  logic                                    halt_i,             
    input  logic                                    flush_dcache_i,     
    output exception_t                              exception_o,        
    output logic                                    dirty_fp_state_o,   
    input  logic                                    single_step_i,      
    
    input  scoreboard_entry_t [NR_COMMIT_PORTS-1:0] commit_instr_i,     
    output logic [NR_COMMIT_PORTS-1:0]              commit_ack_o,       
    
    output  logic [NR_COMMIT_PORTS-1:0][4:0]        waddr_o,            
    output  logic [NR_COMMIT_PORTS-1:0][riscv::XLEN-1:0] wdata_o,       
    output  logic [NR_COMMIT_PORTS-1:0]             we_gpr_o,           
    output  logic [NR_COMMIT_PORTS-1:0]             we_fpr_o,           
    
    input  amo_resp_t                               amo_resp_i,         
    
    output logic [riscv::VLEN-1:0]                  pc_o,
    
    output fu_op                                    csr_op_o,           
    output riscv::xlen_t                            csr_wdata_o,        
    input  riscv::xlen_t                            csr_rdata_i,        
    input  exception_t                              csr_exception_i,    
    output logic                                    csr_write_fflags_o, 
    
    output logic                                    commit_lsu_o,       
    input  logic                                    commit_lsu_ready_i, 
    output logic [TRANS_ID_BITS-1:0]                commit_tran_id_o,   
    output logic                                    amo_valid_commit_o, 
    input  logic                                    no_st_pending_i,    
    output logic                                    commit_csr_o,       
    output logic                                    fence_i_o,          
    output logic                                    fence_o,            
    output logic                                    flush_commit_o,     
    output logic                                    sfence_vma_o        
);
    for (genvar i = 0; i < NR_COMMIT_PORTS; i++) begin : gen_waddr
      assign waddr_o[i] = commit_instr_i[i].rd[4:0];
    end
    assign pc_o       = commit_instr_i[0].pc;
    
    always_comb begin : dirty_fp_state
      dirty_fp_state_o = 1'b0;
      for (int i = 0; i < NR_COMMIT_PORTS; i++) begin
        dirty_fp_state_o |= commit_ack_o[i] & (commit_instr_i[i].fu inside {FPU, FPU_VEC} || is_rd_fpr(commit_instr_i[i].op));
      end
    end
    assign commit_tran_id_o = commit_instr_i[0].trans_id;
    logic instr_0_is_amo;
    assign instr_0_is_amo = is_amo(commit_instr_i[0].op);
    
    
    
    
    always_comb begin : commit
        
        commit_ack_o[0]    = 1'b0;
        commit_ack_o[1]    = 1'b0;
        amo_valid_commit_o = 1'b0;
        we_gpr_o[0]        = 1'b0;
        we_gpr_o[1]        = 1'b0;
        we_fpr_o           = '{default: 1'b0};
        commit_lsu_o       = 1'b0;
        commit_csr_o       = 1'b0;
        
        wdata_o[0]      = (amo_resp_i.ack) ? amo_resp_i.result[riscv::XLEN-1:0] : commit_instr_i[0].result;
        wdata_o[1]      = commit_instr_i[1].result;
        csr_op_o        = ADD; 
        csr_wdata_o        = {riscv::XLEN{1'b0}};
        fence_i_o          = 1'b0;
        fence_o            = 1'b0;
        sfence_vma_o       = 1'b0;
        csr_write_fflags_o = 1'b0;
        flush_commit_o  = 1'b0;
        
        
        if (commit_instr_i[0].valid && !commit_instr_i[0].ex.valid && !halt_i) begin
            
            
            commit_ack_o[0] = 1'b1;
            if (is_rd_fpr(commit_instr_i[0].op)) begin
                we_fpr_o[0] = 1'b1;
            end else begin
                we_gpr_o[0] = 1'b1;
            end
            
            if (commit_instr_i[0].fu == STORE && !instr_0_is_amo) begin
                
                if (commit_lsu_ready_i) begin
                    commit_ack_o[0] = 1'b1;
                    commit_lsu_o = 1'b1;
                
                end else begin
                    commit_ack_o[0] = 1'b0;
                end
            end
            
            
            
            if (commit_instr_i[0].fu inside {FPU, FPU_VEC}) begin
                
                csr_wdata_o = {{riscv::XLEN-5{1'b0}}, commit_instr_i[0].ex.cause[4:0]};
                csr_write_fflags_o = 1'b1;
                commit_ack_o[0] = 1'b1;
            end
            
            
            
            
            
            if (commit_instr_i[0].fu == CSR) begin
                
                csr_op_o     = commit_instr_i[0].op;
                csr_wdata_o  = commit_instr_i[0].result;
                if (!csr_exception_i.valid) begin
                  commit_csr_o = 1'b1;
                  wdata_o[0]   = csr_rdata_i;
                  commit_ack_o[0] = 1'b1;
                end else begin
                  commit_ack_o[0] = 1'b0;
                  we_gpr_o[0] = 1'b0;
                end
            end
            
            
            
            
            
            
            if (commit_instr_i[0].op == SFENCE_VMA) begin
                
                sfence_vma_o = no_st_pending_i;
                
                commit_ack_o[0] = no_st_pending_i;
            end
            
            
            
            
            
            
            
            if (commit_instr_i[0].op == FENCE_I || (flush_dcache_i && commit_instr_i[0].fu != STORE)) begin
                commit_ack_o[0] = no_st_pending_i;
                
                fence_i_o = no_st_pending_i;
            end
            
            
            
            
            
            if (commit_instr_i[0].op == FENCE) begin
                commit_ack_o[0] = no_st_pending_i;
                
                fence_o = no_st_pending_i;
            end
            
            
            
            if (RVA && instr_0_is_amo) begin
                
                commit_ack_o[0] = amo_resp_i.ack;
                
                flush_commit_o = amo_resp_i.ack;
                amo_valid_commit_o = 1'b1;
                we_gpr_o[0] = amo_resp_i.ack;
            end
        end
        if (NR_COMMIT_PORTS > 1) begin
            
            
            
            
            
            if (commit_ack_o[0] && commit_instr_i[1].valid
                                && !halt_i
                                && !(commit_instr_i[0].fu inside {CSR})
                                && !flush_dcache_i
                                && !instr_0_is_amo
                                && !single_step_i) begin
                
                
                if (!exception_o.valid && !commit_instr_i[1].ex.valid
                                       && (commit_instr_i[1].fu inside {ALU, LOAD, CTRL_FLOW, MULT, FPU, FPU_VEC})) begin
                    if (is_rd_fpr(commit_instr_i[1].op))
                        we_fpr_o[1] = 1'b1;
                    else
                        we_gpr_o[1] = 1'b1;
                    commit_ack_o[1] = 1'b1;
                    
                    
                    if (commit_instr_i[1].fu inside {FPU, FPU_VEC}) begin
                        if (csr_write_fflags_o)
                            csr_wdata_o = {{riscv::XLEN-5{1'b0}}, (commit_instr_i[0].ex.cause[4:0] | commit_instr_i[1].ex.cause[4:0])};
                        else
                            csr_wdata_o = {{riscv::XLEN-5{1'b0}}, commit_instr_i[1].ex.cause[4:0]};
                        csr_write_fflags_o = 1'b1;
                    end
                end
            end
        end
    end
    
    
    
    
    always_comb begin : exception_handling
        
        
        
        exception_o.valid = 1'b0;
        exception_o.cause = '0;
        exception_o.tval  = '0;
        
        if (commit_instr_i[0].valid) begin
            
            
            
            if (csr_exception_i.valid) begin
                exception_o      = csr_exception_i;
                
                
                
                exception_o.tval = commit_instr_i[0].ex.tval;
            end
            
            
            
            
            
            if (commit_instr_i[0].ex.valid) begin
                exception_o = commit_instr_i[0].ex;
            end
        end
        
        
        if (halt_i) begin
            exception_o.valid = 1'b0;
        end
    end
endmodule
module wt_dcache_ctrl import ariane_pkg::*; import wt_cache_pkg::*; #(
  parameter logic [CACHE_ID_WIDTH-1:0]  RdTxId    = 1,                              
  parameter ariane_pkg::ariane_cfg_t    ArianeCfg = ariane_pkg::ArianeDefaultConfig 
) (
  input  logic                            clk_i,          
  input  logic                            rst_ni,         
  input  logic                            cache_en_i,
  
  input  dcache_req_i_t                   req_port_i,
  output dcache_req_o_t                   req_port_o,
  
  output logic                            miss_req_o,
  input  logic                            miss_ack_i,
  output logic                            miss_we_o,       
  output logic [63:0]                     miss_wdata_o,    
  output logic [DCACHE_SET_ASSOC-1:0]     miss_vld_bits_o, 
  output logic [riscv::PLEN-1:0]          miss_paddr_o,
  output logic                            miss_nc_o,       
  output logic [2:0]                      miss_size_o,     
  output logic [CACHE_ID_WIDTH-1:0]       miss_id_o,       
  input  logic                            miss_replay_i,   
  input  logic                            miss_rtrn_vld_i, 
  
  input  logic                            wr_cl_vld_i,
  
  output logic [DCACHE_TAG_WIDTH-1:0]     rd_tag_o,        
  output logic [DCACHE_CL_IDX_WIDTH-1:0]  rd_idx_o,
  output logic [DCACHE_OFFSET_WIDTH-1:0]  rd_off_o,
  output logic                            rd_req_o,        
  output logic                            rd_tag_only_o,   
  input  logic                            rd_ack_i,
  input  logic [63:0]                     rd_data_i,
  input  logic [DCACHE_SET_ASSOC-1:0]     rd_vld_bits_i,
  input  logic [DCACHE_SET_ASSOC-1:0]     rd_hit_oh_i
);
  
  typedef enum logic[2:0] {IDLE, READ, MISS_REQ, MISS_WAIT, KILL_MISS, KILL_MISS_ACK, REPLAY_REQ, REPLAY_READ} state_e;
  state_e state_d, state_q;
  logic [DCACHE_TAG_WIDTH-1:0]    address_tag_d, address_tag_q;
  logic [DCACHE_CL_IDX_WIDTH-1:0] address_idx_d, address_idx_q;
  logic [DCACHE_OFFSET_WIDTH-1:0] address_off_d, address_off_q;
  logic [DCACHE_SET_ASSOC-1:0]    vld_data_d,    vld_data_q;
  logic save_tag, rd_req_d, rd_req_q, rd_ack_d, rd_ack_q;
  logic [1:0] data_size_d, data_size_q;
  
  assign vld_data_d    = (rd_req_q)            ? rd_vld_bits_i                                                      : vld_data_q;
  assign address_tag_d = (save_tag)            ? req_port_i.address_tag                                             : address_tag_q;
  assign address_idx_d = (req_port_o.data_gnt) ? req_port_i.address_index[DCACHE_INDEX_WIDTH-1:DCACHE_OFFSET_WIDTH] : address_idx_q;
  assign address_off_d = (req_port_o.data_gnt) ? req_port_i.address_index[DCACHE_OFFSET_WIDTH-1:0]                  : address_off_q;
  assign data_size_d   = (req_port_o.data_gnt) ? req_port_i.data_size                                               : data_size_q;
  assign rd_tag_o      = address_tag_d;
  assign rd_idx_o      = address_idx_d;
  assign rd_off_o      = address_off_d;
  assign req_port_o.data_rdata = rd_data_i;
  
  assign miss_vld_bits_o       = vld_data_q;
  assign miss_paddr_o          = {address_tag_q, address_idx_q, address_off_q};
  assign miss_size_o           = (miss_nc_o) ? data_size_q : 3'b111;
  
  assign miss_nc_o = (~cache_en_i) | (~ariane_pkg::is_inside_cacheable_regions(ArianeCfg, {{{64-DCACHE_TAG_WIDTH}{1'b0}}, address_tag_q, {DCACHE_INDEX_WIDTH{1'b0}}}));
  assign miss_we_o    = '0;
  assign miss_wdata_o = '0;
  assign miss_id_o    = RdTxId;
  assign rd_req_d     = rd_req_o;
  assign rd_ack_d     = rd_ack_i;
  assign rd_tag_only_o = '0;
  always_comb begin : p_fsm
    
    state_d                = state_q;
    save_tag               = 1'b0;
    rd_req_o               = 1'b0;
    miss_req_o             = 1'b0;
    req_port_o.data_rvalid = 1'b0;
    req_port_o.data_gnt    = 1'b0;
    
    unique case (state_q)
        
        
        IDLE: begin
          if (req_port_i.data_req) begin
            rd_req_o = 1'b1;
            
            if (rd_ack_i) begin
              state_d = READ;
              req_port_o.data_gnt = 1'b1;
            end
          end
        end
        
        
        
        
        
        
        READ, REPLAY_READ: begin
          
          rd_req_o = 1'b1;
          
          if(req_port_i.kill_req) begin
            state_d = IDLE;
            req_port_o.data_rvalid = 1'b1;
          end else if(req_port_i.tag_valid | state_q==REPLAY_READ) begin
            save_tag = (state_q!=REPLAY_READ);
            if(wr_cl_vld_i || !rd_ack_q) begin
              state_d = REPLAY_REQ;
            
            end else if((|rd_hit_oh_i) && cache_en_i) begin
              state_d = IDLE;
              req_port_o.data_rvalid = 1'b1;
              
              if (rd_ack_i && req_port_i.data_req) begin
                state_d = READ;
                req_port_o.data_gnt = 1'b1;
              end
            
            end else begin
              state_d = MISS_REQ;
            end
          end
        end
        
        
        MISS_REQ: begin
          miss_req_o = 1'b1;
          if(req_port_i.kill_req) begin
            req_port_o.data_rvalid = 1'b1;
            if(miss_ack_i) begin
              state_d = KILL_MISS;
            end else begin
              state_d = KILL_MISS_ACK;
            end
          end else if(miss_replay_i) begin
            state_d  = REPLAY_REQ;
          end else if(miss_ack_i) begin
            state_d  = MISS_WAIT;
          end
        end
        
        
        
        MISS_WAIT: begin
          if(req_port_i.kill_req) begin
            req_port_o.data_rvalid = 1'b1;
            if(miss_rtrn_vld_i) begin
              state_d = IDLE;
            end else begin
              state_d = KILL_MISS;
            end
          end else if(miss_rtrn_vld_i) begin
            state_d = IDLE;
            req_port_o.data_rvalid = 1'b1;
          end
        end
        
        
        REPLAY_REQ: begin
          rd_req_o = 1'b1;
          if (req_port_i.kill_req) begin
            req_port_o.data_rvalid = 1'b1;
            state_d = IDLE;
          end else if(rd_ack_i) begin
            state_d = REPLAY_READ;
          end
        end
        
        KILL_MISS_ACK: begin
          miss_req_o = 1'b1;
          
          
          if(miss_replay_i) begin
            state_d = IDLE;
          end else if(miss_ack_i) begin
            state_d = KILL_MISS;
          end
        end
        
        
        
        
        KILL_MISS: begin
          if (miss_rtrn_vld_i) begin
            state_d = IDLE;
          end
        end
        default: begin
          
          state_d = IDLE;
        end
    endcase 
  end
  always_ff @(posedge clk_i or negedge rst_ni) begin : p_regs
    if(!rst_ni) begin
      state_q          <= IDLE;
      address_tag_q    <= '0;
      address_idx_q    <= '0;
      address_off_q    <= '0;
      vld_data_q       <= '0;
      data_size_q      <= '0;
      rd_req_q         <= '0;
      rd_ack_q         <= '0;
    end else begin
      state_q          <= state_d;
      address_tag_q    <= address_tag_d;
      address_idx_q    <= address_idx_d;
      address_off_q    <= address_off_d;
      vld_data_q       <= vld_data_d;
      data_size_q      <= data_size_d;
      rd_req_q         <= rd_req_d;
      rd_ack_q         <= rd_ack_d;
    end
  end
endmodule 
module wt_dcache_mem import ariane_pkg::*; import wt_cache_pkg::*; #(
  parameter bit          Axi64BitCompliant  = 1'b0, 
  parameter int unsigned NumPorts           = 3
) (
  input  logic                                              clk_i,
  input  logic                                              rst_ni,
  
  input  logic  [NumPorts-1:0][DCACHE_TAG_WIDTH-1:0]        rd_tag_i,           
  input  logic  [NumPorts-1:0][DCACHE_CL_IDX_WIDTH-1:0]     rd_idx_i,
  input  logic  [NumPorts-1:0][DCACHE_OFFSET_WIDTH-1:0]     rd_off_i,
  input  logic  [NumPorts-1:0]                              rd_req_i,           
  input  logic  [NumPorts-1:0]                              rd_tag_only_i,      
  input  logic  [NumPorts-1:0]                              rd_prio_i,          
  output logic  [NumPorts-1:0]                              rd_ack_o,
  output logic                [DCACHE_SET_ASSOC-1:0]        rd_vld_bits_o,
  output logic                [DCACHE_SET_ASSOC-1:0]        rd_hit_oh_o,
  output logic                [63:0]                        rd_data_o,
  
  input  logic                                              wr_cl_vld_i,
  input  logic                                              wr_cl_nc_i,         
  input  logic                [DCACHE_SET_ASSOC-1:0]        wr_cl_we_i,         
  input  logic                [DCACHE_TAG_WIDTH-1:0]        wr_cl_tag_i,
  input  logic                [DCACHE_CL_IDX_WIDTH-1:0]     wr_cl_idx_i,
  input  logic                [DCACHE_OFFSET_WIDTH-1:0]     wr_cl_off_i,
  input  logic                [DCACHE_LINE_WIDTH-1:0]       wr_cl_data_i,
  input  logic                [DCACHE_LINE_WIDTH/8-1:0]     wr_cl_data_be_i,
  input  logic                [DCACHE_SET_ASSOC-1:0]        wr_vld_bits_i,
  
  input  logic                [DCACHE_SET_ASSOC-1:0]        wr_req_i,           
  output logic                                              wr_ack_o,
  input  logic                [DCACHE_CL_IDX_WIDTH-1:0]     wr_idx_i,
  input  logic                [DCACHE_OFFSET_WIDTH-1:0]     wr_off_i,
  input  logic                [63:0]                        wr_data_i,
  input  logic                [7:0]                         wr_data_be_i,
  
  input wbuffer_t             [DCACHE_WBUF_DEPTH-1:0]       wbuffer_data_i
);
  logic [DCACHE_NUM_BANKS-1:0]                                  bank_req;
  logic [DCACHE_NUM_BANKS-1:0]                                  bank_we;
  logic [DCACHE_NUM_BANKS-1:0][DCACHE_SET_ASSOC-1:0][7:0]       bank_be;
  logic [DCACHE_NUM_BANKS-1:0][DCACHE_CL_IDX_WIDTH-1:0]         bank_idx;
  logic [DCACHE_CL_IDX_WIDTH-1:0]                               bank_idx_d, bank_idx_q;
  logic [DCACHE_OFFSET_WIDTH-1:0]                               bank_off_d, bank_off_q;
  logic [DCACHE_NUM_BANKS-1:0][DCACHE_SET_ASSOC-1:0][63:0]      bank_wdata;                   
  logic [DCACHE_NUM_BANKS-1:0][DCACHE_SET_ASSOC-1:0][63:0]      bank_rdata;                   
  logic [DCACHE_SET_ASSOC-1:0][63:0]                            rdata_cl;                     
  logic [DCACHE_TAG_WIDTH-1:0]                                  rd_tag;
  logic [DCACHE_SET_ASSOC-1:0]                                  vld_req;                      
  logic                                                         vld_we;                       
  logic [DCACHE_SET_ASSOC-1:0]                                  vld_wdata;                    
  logic [DCACHE_SET_ASSOC-1:0][DCACHE_TAG_WIDTH-1:0]            tag_rdata;                    
  logic                       [DCACHE_CL_IDX_WIDTH-1:0]         vld_addr;                     
  logic [$clog2(NumPorts)-1:0]                                  vld_sel_d, vld_sel_q;
  logic [DCACHE_WBUF_DEPTH-1:0]                                 wbuffer_hit_oh;
  logic [7:0]                                                   wbuffer_be;
  logic [63:0]                                                  wbuffer_rdata, rdata;
  logic [63:0]                                                  wbuffer_cmp_addr;
  logic                                                         cmp_en_d, cmp_en_q;
  logic                                                         rd_acked;
  logic [NumPorts-1:0]                                          bank_collision, rd_req_masked, rd_req_prio;
  
  
  
  
  
  
  
  for (genvar k=0;k<DCACHE_NUM_BANKS;k++) begin : gen_bank
    for (genvar j=0;j<DCACHE_SET_ASSOC;j++) begin : gen_bank_way
      assign bank_be[k][j]   = (wr_cl_we_i[j] & wr_cl_vld_i)  ? wr_cl_data_be_i[k*8 +: 8] :
                               (wr_req_i[j]   & wr_ack_o)     ? wr_data_be_i              :
                                                                '0;
      assign bank_wdata[k][j] = (wr_cl_we_i[j] & wr_cl_vld_i) ?  wr_cl_data_i[k*64 +: 64] :
                                                                 wr_data_i;
    end
  end
  assign vld_wdata  = wr_vld_bits_i;
  assign vld_addr   = (wr_cl_vld_i) ? wr_cl_idx_i   : rd_idx_i[vld_sel_d];
  assign rd_tag     = rd_tag_i[vld_sel_q]; 
  assign bank_off_d = (wr_cl_vld_i) ? wr_cl_off_i   : rd_off_i[vld_sel_d];
  assign bank_idx_d = (wr_cl_vld_i) ? wr_cl_idx_i   : rd_idx_i[vld_sel_d];
  assign vld_req    = (wr_cl_vld_i) ? wr_cl_we_i    : (rd_acked) ? '1 : '0;
  
  
  assign rd_req_prio   = rd_req_i & rd_prio_i;
  assign rd_req_masked = (|rd_req_prio) ? rd_req_prio : rd_req_i;
  logic rd_req;
  rr_arb_tree #(
    .NumIn     (NumPorts),
    .DataWidth (1)
  ) i_rr_arb_tree (
    .clk_i  (clk_i   ),
    .rst_ni (rst_ni  ),
    .flush_i('0      ),
    .rr_i   ('0      ),
    .req_i  (rd_req_masked ),
    .gnt_o  (rd_ack_o      ),
    .data_i ('0            ),
    .gnt_i  (~wr_cl_vld_i  ),
    .req_o  (rd_req        ),
    .data_o (              ),
    .idx_o  (vld_sel_d     )
  );
  assign rd_acked = rd_req & ~wr_cl_vld_i;
  always_comb begin : p_bank_req
    vld_we   = wr_cl_vld_i;
    bank_req = '0;
    wr_ack_o = '0;
    bank_we  = '0;
    bank_idx = '{default:wr_idx_i};
    for(int k=0; k<NumPorts; k++) begin
      bank_collision[k] = rd_off_i[k][DCACHE_OFFSET_WIDTH-1:3] == wr_off_i[DCACHE_OFFSET_WIDTH-1:3];
    end
    if(wr_cl_vld_i & |wr_cl_we_i) begin
      bank_req = '1;
      bank_we  = '1;
      bank_idx = '{default:wr_cl_idx_i};
    end else begin
      if(rd_acked) begin
        if(!rd_tag_only_i[vld_sel_d]) begin
          bank_req                                               = dcache_cl_bin2oh(rd_off_i[vld_sel_d][DCACHE_OFFSET_WIDTH-1:3]);
          bank_idx[rd_off_i[vld_sel_d][DCACHE_OFFSET_WIDTH-1:3]] = rd_idx_i[vld_sel_d];
        end
      end
      if(|wr_req_i) begin
        if(rd_tag_only_i[vld_sel_d] || !(rd_ack_o[vld_sel_d] && bank_collision[vld_sel_d])) begin
          wr_ack_o = 1'b1;
          bank_req |= dcache_cl_bin2oh(wr_off_i[DCACHE_OFFSET_WIDTH-1:3]);
          bank_we   = dcache_cl_bin2oh(wr_off_i[DCACHE_OFFSET_WIDTH-1:3]);
        end
      end
    end
  end
  logic [DCACHE_OFFSET_WIDTH-1:0]       wr_cl_off;
  logic [$clog2(DCACHE_WBUF_DEPTH)-1:0] wbuffer_hit_idx;
  logic [$clog2(DCACHE_SET_ASSOC)-1:0]  rd_hit_idx;
  assign cmp_en_d = (|vld_req) & ~vld_we;
  
  assign wbuffer_cmp_addr = (wr_cl_vld_i) ? {wr_cl_tag_i, wr_cl_idx_i, wr_cl_off_i} :
                                            {rd_tag, bank_idx_q, bank_off_q};
  
  for (genvar i=0;i<DCACHE_SET_ASSOC;i++) begin : gen_tag_cmpsel
    
    assign rd_hit_oh_o[i] = (rd_tag == tag_rdata[i]) & rd_vld_bits_o[i]  & cmp_en_q;
    
    assign rdata_cl[i] = bank_rdata[bank_off_q[DCACHE_OFFSET_WIDTH-1:3]][i];
  end
  for(genvar k=0; k<DCACHE_WBUF_DEPTH; k++) begin : gen_wbuffer_hit
    assign wbuffer_hit_oh[k] = (|wbuffer_data_i[k].valid) & (wbuffer_data_i[k].wtag == (wbuffer_cmp_addr >> 3));
  end
  lzc #(
    .WIDTH ( DCACHE_WBUF_DEPTH )
  ) i_lzc_wbuffer_hit (
    .in_i    ( wbuffer_hit_oh   ),
    .cnt_o   ( wbuffer_hit_idx  ),
    .empty_o (                  )
  );
  lzc #(
    .WIDTH ( DCACHE_SET_ASSOC )
  ) i_lzc_rd_hit (
    .in_i    ( rd_hit_oh_o  ),
    .cnt_o   ( rd_hit_idx   ),
    .empty_o (              )
  );
  assign wbuffer_rdata = wbuffer_data_i[wbuffer_hit_idx].data;
  assign wbuffer_be    = (|wbuffer_hit_oh) ? wbuffer_data_i[wbuffer_hit_idx].valid : '0;
  if (Axi64BitCompliant) begin : gen_axi_off
      assign wr_cl_off     = (wr_cl_nc_i) ? '0 : wr_cl_off_i[DCACHE_OFFSET_WIDTH-1:3];
  end else begin  : gen_piton_off
      assign wr_cl_off     = wr_cl_off_i[DCACHE_OFFSET_WIDTH-1:3];
  end
  assign rdata         = (wr_cl_vld_i)  ? wr_cl_data_i[wr_cl_off*64 +: 64] :
                                          rdata_cl[rd_hit_idx];
  
  for(genvar k=0; k<8; k++) begin : gen_rd_data
    assign rd_data_o[8*k +: 8] = (wbuffer_be[k]) ? wbuffer_rdata[8*k +: 8] : rdata[8*k +: 8];
  end
  logic [DCACHE_TAG_WIDTH:0] vld_tag_rdata [DCACHE_SET_ASSOC-1:0];
  for (genvar k = 0; k < DCACHE_NUM_BANKS; k++) begin : gen_data_banks
    
    sram #(
      .DATA_WIDTH ( ariane_pkg::DCACHE_SET_ASSOC * 64 ),
      .NUM_WORDS  ( wt_cache_pkg::DCACHE_NUM_WORDS    )
    ) i_data_sram (
      .clk_i      ( clk_i               ),
      .rst_ni     ( rst_ni              ),
      .req_i      ( bank_req   [k]      ),
      .we_i       ( bank_we    [k]      ),
      .addr_i     ( bank_idx   [k]      ),
      .wdata_i    ( bank_wdata [k]      ),
      .be_i       ( bank_be    [k]      ),
      .rdata_o    ( bank_rdata [k]      )
    );
  end
  for (genvar i = 0; i < DCACHE_SET_ASSOC; i++) begin : gen_tag_srams
    assign tag_rdata[i]     = vld_tag_rdata[i][DCACHE_TAG_WIDTH-1:0];
    assign rd_vld_bits_o[i] = vld_tag_rdata[i][DCACHE_TAG_WIDTH];
    
    sram #(
      
      .DATA_WIDTH ( ariane_pkg::DCACHE_TAG_WIDTH + 1 ),
      .NUM_WORDS  ( wt_cache_pkg::DCACHE_NUM_WORDS   )
    ) i_tag_sram (
      .clk_i     ( clk_i               ),
      .rst_ni    ( rst_ni              ),
      .req_i     ( vld_req[i]          ),
      .we_i      ( vld_we              ),
      .addr_i    ( vld_addr            ),
      .wdata_i   ( {vld_wdata[i], wr_cl_tag_i} ),
      .be_i      ( '1                  ),
      .rdata_o   ( vld_tag_rdata[i]    )
    );
  end
  always_ff @(posedge clk_i or negedge rst_ni) begin : p_regs
    if(!rst_ni) begin
      bank_idx_q <= '0;
      bank_off_q <= '0;
      vld_sel_q  <= '0;
      cmp_en_q   <= '0;
    end else begin
      bank_idx_q <= bank_idx_d;
      bank_off_q <= bank_off_d;
      vld_sel_q  <= vld_sel_d ;
      cmp_en_q   <= cmp_en_d;
    end
  end
endmodule 
module wt_dcache_missunit import ariane_pkg::*; import wt_cache_pkg::*; #(
  parameter bit                         Axi64BitCompliant  = 1'b0, 
  parameter logic [CACHE_ID_WIDTH-1:0]  AmoTxId            = 1,    
  parameter int unsigned                NumPorts           = 3     
) (
  input  logic                                       clk_i,       
  input  logic                                       rst_ni,      
  
  input  logic                                       enable_i,    
  input  logic                                       flush_i,     
  output logic                                       flush_ack_o, 
  output logic                                       miss_o,      
  
  input  logic                                       wbuffer_empty_i,
  output logic                                       cache_en_o,  
  
  input  amo_req_t                                   amo_req_i,
  output amo_resp_t                                  amo_resp_o,
  
  input  logic [NumPorts-1:0]                        miss_req_i,
  output logic [NumPorts-1:0]                        miss_ack_o,
  input  logic [NumPorts-1:0]                        miss_nc_i,
  input  logic [NumPorts-1:0]                        miss_we_i,
  input  logic [NumPorts-1:0][63:0]                  miss_wdata_i,
  input  logic [NumPorts-1:0][riscv::PLEN-1:0]       miss_paddr_i,
  input  logic [NumPorts-1:0][DCACHE_SET_ASSOC-1:0]  miss_vld_bits_i,
  input  logic [NumPorts-1:0][2:0]                   miss_size_i,
  input  logic [NumPorts-1:0][CACHE_ID_WIDTH-1:0]    miss_id_i,          
  
  output logic [NumPorts-1:0]                        miss_replay_o,
  
  output logic [NumPorts-1:0]                        miss_rtrn_vld_o,
  output logic [CACHE_ID_WIDTH-1:0]                  miss_rtrn_id_o,     
  
  input  logic [DCACHE_MAX_TX-1:0][riscv::PLEN-1:0]  tx_paddr_i,         
  input  logic [DCACHE_MAX_TX-1:0]                   tx_vld_i,           
  
  output logic                                       wr_cl_vld_o,        
  output logic                                       wr_cl_nc_o,         
  output logic [DCACHE_SET_ASSOC-1:0]                wr_cl_we_o,         
  output logic [DCACHE_TAG_WIDTH-1:0]                wr_cl_tag_o,
  output logic [DCACHE_CL_IDX_WIDTH-1:0]             wr_cl_idx_o,
  output logic [DCACHE_OFFSET_WIDTH-1:0]             wr_cl_off_o,
  output logic [DCACHE_LINE_WIDTH-1:0]               wr_cl_data_o,
  output logic [DCACHE_LINE_WIDTH/8-1:0]             wr_cl_data_be_o,
  output logic [DCACHE_SET_ASSOC-1:0]                wr_vld_bits_o,
  
  input  logic                                       mem_rtrn_vld_i,
  input  dcache_rtrn_t                               mem_rtrn_i,
  output logic                                       mem_data_req_o,
  input  logic                                       mem_data_ack_i,
  output dcache_req_t                                mem_data_o
);
  
  typedef enum logic[2:0] {IDLE, DRAIN, AMO,  FLUSH, STORE_WAIT, LOAD_WAIT, AMO_WAIT} state_e;
  state_e state_d, state_q;
  
  typedef struct packed {
    logic [riscv::PLEN-1:0]              paddr   ;
    logic [2:0]                          size    ;
    logic [DCACHE_SET_ASSOC-1:0]         vld_bits;
    logic [CACHE_ID_WIDTH-1:0]          id      ;
    logic                                nc      ;
    logic [$clog2(DCACHE_SET_ASSOC)-1:0] repl_way;
    logic [$clog2(NumPorts)-1:0]        miss_port_idx;
  } mshr_t;
  mshr_t mshr_d, mshr_q;
  logic [$clog2(DCACHE_SET_ASSOC)-1:0] repl_way, inv_way, rnd_way;
  logic mshr_vld_d, mshr_vld_q, mshr_vld_q1;
  logic mshr_allocate;
  logic update_lfsr, all_ways_valid;
  logic enable_d, enable_q;
  logic flush_ack_d, flush_ack_q;
  logic flush_en, flush_done;
  logic mask_reads, lock_reqs;
  logic amo_sel, miss_is_write;
  logic amo_req_d, amo_req_q;
  logic [63:0] amo_data, amo_rtrn_mux;
  logic [riscv::PLEN-1:0] tmp_paddr;
  logic [$clog2(NumPorts)-1:0] miss_port_idx;
  logic [DCACHE_CL_IDX_WIDTH-1:0] cnt_d, cnt_q;
  logic [NumPorts-1:0] miss_req_masked_d, miss_req_masked_q;
  logic inv_vld, inv_vld_all, cl_write_en;
  logic load_ack, store_ack, amo_ack;
  logic [NumPorts-1:0] mshr_rdrd_collision_d, mshr_rdrd_collision_q;
  logic [NumPorts-1:0] mshr_rdrd_collision;
  logic tx_rdwr_collision, mshr_rdwr_collision;
  assign cache_en_o      = enable_q;
  assign cnt_d           = (flush_en) ? cnt_q + 1 : '0;
  assign flush_done      = (cnt_q == wt_cache_pkg::DCACHE_NUM_WORDS-1);
  assign miss_req_masked_d = (lock_reqs)  ? miss_req_masked_q      :
                             (mask_reads) ? miss_we_i & miss_req_i : miss_req_i;
  assign miss_is_write     = miss_we_i[miss_port_idx];
  
  lzc #(
    .WIDTH ( NumPorts )
  ) i_lzc_reqs (
    .in_i    ( miss_req_masked_d ),
    .cnt_o   ( miss_port_idx     ),
    .empty_o (                   )
  );
  always_comb begin : p_ack
    miss_ack_o = '0;
    if (!amo_sel) begin
      miss_ack_o[miss_port_idx] = mem_data_ack_i & mem_data_req_o;
    end
  end
  
  lzc #(
    .WIDTH ( ariane_pkg::DCACHE_SET_ASSOC )
  ) i_lzc_inv (
    .in_i    ( ~miss_vld_bits_i[miss_port_idx] ),
    .cnt_o   ( inv_way                         ),
    .empty_o ( all_ways_valid                  )
  );
  
  lfsr #(
    .LfsrWidth  ( ariane_pkg::DCACHE_SET_ASSOC        ),
    .OutWidth   ( $clog2(ariane_pkg::DCACHE_SET_ASSOC))
  ) i_lfsr_inv (
    .clk_i          ( clk_i       ),
    .rst_ni         ( rst_ni      ),
    .en_i           ( update_lfsr ),
    .out_o          ( rnd_way     )
  );
  assign repl_way               = (all_ways_valid) ? rnd_way : inv_way;
  assign mshr_d.size            = (mshr_allocate)  ? miss_size_i    [miss_port_idx] : mshr_q.size;
  assign mshr_d.paddr           = (mshr_allocate)  ? miss_paddr_i   [miss_port_idx] : mshr_q.paddr;
  assign mshr_d.vld_bits        = (mshr_allocate)  ? miss_vld_bits_i[miss_port_idx] : mshr_q.vld_bits;
  assign mshr_d.id              = (mshr_allocate)  ? miss_id_i      [miss_port_idx] : mshr_q.id;
  assign mshr_d.nc              = (mshr_allocate)  ? miss_nc_i      [miss_port_idx] : mshr_q.nc;
  assign mshr_d.repl_way        = (mshr_allocate)  ? repl_way                       : mshr_q.repl_way;
  assign mshr_d.miss_port_idx   = (mshr_allocate)  ? miss_port_idx                  : mshr_q.miss_port_idx;
  
  assign mshr_vld_d = (mshr_allocate) ? 1'b1 :
                      (load_ack)      ? 1'b0 :
                                        mshr_vld_q;
  assign miss_o     = (mshr_allocate) ? ~miss_nc_i[miss_port_idx] : 1'b0;
  for(genvar k=0; k<NumPorts; k++) begin : gen_rdrd_collision
    assign mshr_rdrd_collision[k]   = (mshr_q.paddr[riscv::PLEN-1:DCACHE_OFFSET_WIDTH] == miss_paddr_i[k][riscv::PLEN-1:DCACHE_OFFSET_WIDTH]) && (mshr_vld_q | mshr_vld_q1);
    assign mshr_rdrd_collision_d[k] = (!miss_req_i[k]) ? 1'b0 : mshr_rdrd_collision_q[k] | mshr_rdrd_collision[k];
  end
  
  
  assign mshr_rdwr_collision = (mshr_q.paddr[riscv::PLEN-1:DCACHE_OFFSET_WIDTH] == miss_paddr_i[NumPorts-1][riscv::PLEN-1:DCACHE_OFFSET_WIDTH]) && mshr_vld_q;
  
  always_comb begin : p_tx_coll
    tx_rdwr_collision = 1'b0;
    for(int k=0; k<DCACHE_MAX_TX; k++) begin
      tx_rdwr_collision |= (miss_paddr_i[miss_port_idx][riscv::PLEN-1:DCACHE_OFFSET_WIDTH] == tx_paddr_i[k][riscv::PLEN-1:DCACHE_OFFSET_WIDTH]) && tx_vld_i[k];
    end
  end
  
  assign amo_data = (amo_req_i.size==2'b10) ? {amo_req_i.operand_b[0 +: 32],
                                               amo_req_i.operand_b[0 +: 32]} :
                                               amo_req_i.operand_b;
  
  if (Axi64BitCompliant) begin : gen_axi_rtrn_mux
    assign amo_rtrn_mux = mem_rtrn_i.data[0 +: 64];
  end else begin : gen_piton_rtrn_mux
    assign amo_rtrn_mux = mem_rtrn_i.data[amo_req_i.operand_a[DCACHE_OFFSET_WIDTH-1:3]*64 +: 64];
  end
  
  assign amo_resp_o.result = (amo_req_i.size==2'b10) ? {{32{amo_rtrn_mux[amo_req_i.operand_a[2]*32 + 31]}},
                                                            amo_rtrn_mux[amo_req_i.operand_a[2]*32 +: 32]} :
                                                       amo_rtrn_mux;
  assign amo_req_d = amo_req_i.req;
  
  assign mem_data_o.tid    = (amo_sel) ? AmoTxId             : miss_id_i[miss_port_idx];
  assign mem_data_o.nc     = (amo_sel) ? 1'b1                : miss_nc_i[miss_port_idx];
  assign mem_data_o.way    = (amo_sel) ? '0                  : repl_way;
  assign mem_data_o.data   = (amo_sel) ? amo_data            : miss_wdata_i[miss_port_idx];
  assign mem_data_o.size   = (amo_sel) ? amo_req_i.size      : miss_size_i [miss_port_idx];
  assign mem_data_o.amo_op = (amo_sel) ? amo_req_i.amo_op    : AMO_NONE;
  assign tmp_paddr         = (amo_sel) ? amo_req_i.operand_a[riscv::PLEN-1:0] : miss_paddr_i[miss_port_idx];
  assign mem_data_o.paddr  = wt_cache_pkg::paddrSizeAlign(tmp_paddr, mem_data_o.size);
  logic sc_fail, sc_pass, sc_backoff_over;
  exp_backoff #(
    .Seed(3),
    .MaxExp(16)
  ) i_exp_backoff (
    .clk_i,
    .rst_ni,
    .set_i     ( sc_fail         ),
    .clr_i     ( sc_pass         ),
    .is_zero_o ( sc_backoff_over )
  );
  
  logic store_sent;
  logic [$clog2(wt_cache_pkg::DCACHE_MAX_TX + 1)-1:0] stores_inflight_d, stores_inflight_q;
  assign store_sent = mem_data_req_o   & mem_data_ack_i & (mem_data_o.rtype == DCACHE_STORE_REQ);
  assign stores_inflight_d = (store_ack && store_sent) ? stores_inflight_q     :
                             (store_ack)               ? stores_inflight_q - 1 :
                             (store_sent)              ? stores_inflight_q + 1 :
                                                         stores_inflight_q;
  
  always_comb begin : p_rtrn_logic
    load_ack        = 1'b0;
    store_ack       = 1'b0;
    amo_ack         = 1'b0;
    inv_vld         = 1'b0;
    inv_vld_all     = 1'b0;
    sc_fail         = 1'b0;
    sc_pass         = 1'b0;
    miss_rtrn_vld_o ='0;
    if (mem_rtrn_vld_i) begin
      unique case (mem_rtrn_i.rtype)
        DCACHE_LOAD_ACK: begin
          if (mshr_vld_q) begin
            load_ack = 1'b1;
            miss_rtrn_vld_o[mshr_q.miss_port_idx] = 1'b1;
          end
        end
        DCACHE_STORE_ACK: begin
          if (stores_inflight_q) begin
            store_ack = 1'b1;
            miss_rtrn_vld_o[NumPorts-1] = 1'b1;
          end
        end
        DCACHE_ATOMIC_ACK: begin
          if (amo_req_q) begin
            amo_ack = 1'b1;
            
            
            if (amo_req_i.amo_op == AMO_SC) begin
              if (amo_resp_o.result) begin
                sc_fail = 1'b1;
              end else begin
                sc_pass = 1'b1;
              end
            end
          end
        end
        DCACHE_INV_REQ: begin
          inv_vld     = mem_rtrn_i.inv.vld | mem_rtrn_i.inv.all;
          inv_vld_all = mem_rtrn_i.inv.all;
        end
        
        
        
        default : begin
        end
      endcase
    end
  end
  
  assign miss_rtrn_id_o           = mem_rtrn_i.tid;
  
  assign wr_cl_nc_o      = mshr_q.nc;
  assign wr_cl_vld_o     = load_ack | (| wr_cl_we_o);
  assign wr_cl_we_o      = (flush_en   )  ? '1                                    :
                           (inv_vld_all)   ? '1                                    :
                           (inv_vld    )   ? dcache_way_bin2oh(mem_rtrn_i.inv.way) :
                           (cl_write_en)   ? dcache_way_bin2oh(mshr_q.repl_way)    :
                                             '0;
  assign wr_vld_bits_o   = (flush_en   )   ? '0                                    :
                           (inv_vld    )   ? '0                                    :
                           (cl_write_en)   ? dcache_way_bin2oh(mshr_q.repl_way)    :
                                              '0;
  assign wr_cl_idx_o     = (flush_en) ? cnt_q                                                        :
                           (inv_vld)  ? mem_rtrn_i.inv.idx[DCACHE_INDEX_WIDTH-1:DCACHE_OFFSET_WIDTH] :
                                        mshr_q.paddr[DCACHE_INDEX_WIDTH-1:DCACHE_OFFSET_WIDTH];
  assign wr_cl_tag_o     = mshr_q.paddr[DCACHE_TAG_WIDTH+DCACHE_INDEX_WIDTH-1:DCACHE_INDEX_WIDTH];
  assign wr_cl_off_o     = mshr_q.paddr[DCACHE_OFFSET_WIDTH-1:0];
  assign wr_cl_data_o    = mem_rtrn_i.data;
  assign wr_cl_data_be_o = (cl_write_en) ? '1 : '0;
  
  assign cl_write_en     = load_ack & ~mshr_q.nc;
  always_comb begin : p_fsm
    
    state_d          = state_q;
    flush_ack_o      = 1'b0;
    mem_data_o.rtype = DCACHE_LOAD_REQ;
    mem_data_req_o   = 1'b0;
    amo_resp_o.ack   = 1'b0;
    miss_replay_o    = '0;
    
    enable_d         = enable_q & enable_i;
    flush_ack_d      = flush_ack_q;
    flush_en         = 1'b0;
    amo_sel          = 1'b0;
    update_lfsr      = 1'b0;
    mshr_allocate    = 1'b0;
    lock_reqs        = 1'b0;
    mask_reads       = mshr_vld_q;
    
    unique case (state_q)
      
      
      IDLE: begin
        if (flush_i || (enable_i && !enable_q)) begin
          if (wbuffer_empty_i && !mshr_vld_q) begin
            flush_ack_d = flush_i;
            state_d     = FLUSH;
          end else begin
            state_d     = DRAIN;
          end
        end else if (amo_req_i.req) begin
          if (wbuffer_empty_i && !mshr_vld_q) begin
            state_d     = AMO;
          end else begin
            state_d     = DRAIN;
          end
        
        end else if (|miss_req_masked_d) begin
          
          if (miss_is_write) begin
            
            if (!mshr_rdwr_collision) begin
              mem_data_req_o            = 1'b1;
              mem_data_o.rtype          = DCACHE_STORE_REQ;
              if (!mem_data_ack_i) begin
                state_d = STORE_WAIT;
              end
            end
          
          
          end else if (!mshr_vld_q || load_ack) begin
            
            
            if (mshr_rdrd_collision_d[miss_port_idx]) begin
              miss_replay_o[miss_port_idx] = 1'b1;
            
            end else if (!tx_rdwr_collision) begin
              mem_data_req_o            = 1'b1;
              mem_data_o.rtype          = DCACHE_LOAD_REQ;
              update_lfsr               = all_ways_valid & mem_data_ack_i;
              mshr_allocate             = mem_data_ack_i;
              if (!mem_data_ack_i) begin
                state_d = LOAD_WAIT;
              end
            end
          end
        end
      end
      
      
      STORE_WAIT: begin
        lock_reqs                 = 1'b1;
        mem_data_req_o            = 1'b1;
        mem_data_o.rtype          = DCACHE_STORE_REQ;
        if (mem_data_ack_i) begin
          state_d = IDLE;
        end
      end
      
      
      LOAD_WAIT: begin
        lock_reqs                 = 1'b1;
        mem_data_req_o            = 1'b1;
        mem_data_o.rtype          = DCACHE_LOAD_REQ;
        if (mem_data_ack_i) begin
          update_lfsr   = all_ways_valid;
          mshr_allocate = 1'b1;
          state_d       = IDLE;
        end
      end
      
      
      
      DRAIN: begin
        mask_reads = 1'b1;
        
        if (|miss_req_masked_d && !mshr_rdwr_collision) begin
          mem_data_req_o            = 1'b1;
          mem_data_o.rtype          = DCACHE_STORE_REQ;
        end
        if (wbuffer_empty_i && !mshr_vld_q) begin
          state_d = IDLE;
        end
      end
      
      
      FLUSH: begin
        
        flush_en   = 1'b1;
        if (flush_done) begin
          state_d     = IDLE;
          flush_ack_o = flush_ack_q;
          flush_ack_d = 1'b0;
          enable_d    = enable_i;
        end
      end
      
      
      AMO: begin
        mem_data_o.rtype = DCACHE_ATOMIC_REQ;
        amo_sel          = 1'b1;
        
        if ((amo_req_i.amo_op != AMO_LR) || sc_backoff_over) begin
          mem_data_req_o   = 1'b1;
          if (mem_data_ack_i) begin
            state_d = AMO_WAIT;
          end
        end
      end
      
      
      AMO_WAIT: begin
        amo_sel = 1'b1;
        if (amo_ack) begin
          amo_resp_o.ack = 1'b1;
          state_d        = IDLE;
        end
      end
      
      default: begin
        
        state_d = IDLE;
      end
    endcase 
  end
always_ff @(posedge clk_i or negedge rst_ni) begin : p_regs
  if (!rst_ni) begin
    state_q               <= FLUSH;
    cnt_q                 <= '0;
    enable_q              <= '0;
    flush_ack_q           <= '0;
    mshr_vld_q            <= '0;
    mshr_vld_q1           <= '0;
    mshr_q                <= '0;
    mshr_rdrd_collision_q <= '0;
    miss_req_masked_q     <= '0;
    amo_req_q             <= '0;
    stores_inflight_q     <= '0;
  end else begin
    state_q               <= state_d;
    cnt_q                 <= cnt_d;
    enable_q              <= enable_d;
    flush_ack_q           <= flush_ack_d;
    mshr_vld_q            <= mshr_vld_d;
    mshr_vld_q1           <= mshr_vld_q;
    mshr_q                <= mshr_d;
    mshr_rdrd_collision_q <= mshr_rdrd_collision_d;
    miss_req_masked_q     <= miss_req_masked_d;
    amo_req_q             <= amo_req_d;
    stores_inflight_q     <= stores_inflight_d;
  end
end
endmodule 
module wt_dcache_wbuffer import ariane_pkg::*; import wt_cache_pkg::*; #(
  parameter ariane_pkg::ariane_cfg_t    ArianeCfg          = ariane_pkg::ArianeDefaultConfig     
) (
  input  logic                               clk_i,          
  input  logic                               rst_ni,         
  input  logic                               cache_en_i,     
  output logic                               empty_o,        
  output logic                               not_ni_o,    
   
  input  dcache_req_i_t                      req_port_i,
  output dcache_req_o_t                      req_port_o,
  
  input  logic                               miss_ack_i,
  output logic [riscv::PLEN-1:0]             miss_paddr_o,
  output logic                               miss_req_o,
  output logic                               miss_we_o,       
  output logic [63:0]                        miss_wdata_o,
  output logic [DCACHE_SET_ASSOC-1:0]        miss_vld_bits_o, 
  output logic                               miss_nc_o,       
  output logic [2:0]                         miss_size_o,     
  output logic [CACHE_ID_WIDTH-1:0]          miss_id_o,       
  
  input  logic                               miss_rtrn_vld_i,
  input  logic [CACHE_ID_WIDTH-1:0]          miss_rtrn_id_i,  
  
  output logic [DCACHE_TAG_WIDTH-1:0]        rd_tag_o,        
  output logic [DCACHE_CL_IDX_WIDTH-1:0]     rd_idx_o,
  output logic [DCACHE_OFFSET_WIDTH-1:0]     rd_off_o,
  output logic                               rd_req_o,        
  output logic                               rd_tag_only_o,   
  input  logic                               rd_ack_i,
  input logic  [63:0]                        rd_data_i,       
  input logic  [DCACHE_SET_ASSOC-1:0]        rd_vld_bits_i,   
  input logic  [DCACHE_SET_ASSOC-1:0]        rd_hit_oh_i,
  
  input logic                                wr_cl_vld_i,
  input logic [DCACHE_CL_IDX_WIDTH-1:0]      wr_cl_idx_i,
  
  output logic [DCACHE_SET_ASSOC-1:0]        wr_req_o,
  input  logic                               wr_ack_i,
  output logic [DCACHE_CL_IDX_WIDTH-1:0]     wr_idx_o,
  output logic [DCACHE_OFFSET_WIDTH-1:0]     wr_off_o,
  output logic [63:0]                        wr_data_o,
  output logic [7:0]                         wr_data_be_o,
  
  output wbuffer_t  [DCACHE_WBUF_DEPTH-1:0]  wbuffer_data_o,
  output logic [DCACHE_MAX_TX-1:0][riscv::PLEN-1:0]     tx_paddr_o,      
  output logic [DCACHE_MAX_TX-1:0]           tx_vld_o
);
  tx_stat_t [DCACHE_MAX_TX-1:0]             tx_stat_d, tx_stat_q;
  wbuffer_t [DCACHE_WBUF_DEPTH-1:0]         wbuffer_d, wbuffer_q;
  logic     [DCACHE_WBUF_DEPTH-1:0]         valid;
  logic     [DCACHE_WBUF_DEPTH-1:0]         dirty;
  logic     [DCACHE_WBUF_DEPTH-1:0]         tocheck;
  logic     [DCACHE_WBUF_DEPTH-1:0]         wbuffer_hit_oh, inval_hit;
  logic     [DCACHE_WBUF_DEPTH-1:0][7:0]    bdirty;
  logic [$clog2(DCACHE_WBUF_DEPTH)-1:0] next_ptr, dirty_ptr, hit_ptr, wr_ptr, check_ptr_d, check_ptr_q, check_ptr_q1, rtrn_ptr;
  logic [CACHE_ID_WIDTH-1:0] tx_id, rtrn_id;
  logic [2:0] bdirty_off;
  logic [7:0] tx_be;
  logic [riscv::PLEN-1:0] wr_paddr, rd_paddr;
  logic [DCACHE_TAG_WIDTH-1:0] rd_tag_d, rd_tag_q;
  logic [DCACHE_SET_ASSOC-1:0] rd_hit_oh_d, rd_hit_oh_q;
  logic check_en_d, check_en_q, check_en_q1;
  logic full, dirty_rd_en, rdy;
  logic rtrn_empty, evict;
  logic [DCACHE_WBUF_DEPTH-1:0] ni_pending_d, ni_pending_q;
  logic wbuffer_wren;
  logic free_tx_slots;
  logic wr_cl_vld_q, wr_cl_vld_d;
  logic [DCACHE_CL_IDX_WIDTH-1:0] wr_cl_idx_q, wr_cl_idx_d;
  logic [riscv::PLEN-1:0] debug_paddr [DCACHE_WBUF_DEPTH-1:0];
  wbuffer_t wbuffer_check_mux, wbuffer_dirty_mux;
  logic [ariane_pkg::DCACHE_TAG_WIDTH-1:0] miss_tag;
  logic is_nc_miss;
  logic is_ni;
  assign miss_tag = miss_paddr_o[ariane_pkg::DCACHE_INDEX_WIDTH+:ariane_pkg::DCACHE_TAG_WIDTH];
  assign is_nc_miss = !ariane_pkg::is_inside_cacheable_regions(ArianeCfg, {{64-DCACHE_TAG_WIDTH{1'b0}}, miss_tag, {DCACHE_INDEX_WIDTH{1'b0}}});
  assign miss_nc_o = !cache_en_i || is_nc_miss; 
  
  assign is_ni = ariane_pkg::is_inside_nonidempotent_regions(ArianeCfg, {{64-DCACHE_TAG_WIDTH{1'b0}}, req_port_i.address_tag, {DCACHE_INDEX_WIDTH{1'b0}}});
  assign miss_we_o       = 1'b1;
  assign miss_vld_bits_o = '0;
  assign wbuffer_data_o  = wbuffer_q;
  for (genvar k=0; k<DCACHE_MAX_TX;k++) begin : gen_tx_vld
    assign tx_vld_o[k]   = tx_stat_q[k].vld;
    assign tx_paddr_o[k] = wbuffer_q[tx_stat_q[k].ptr].wtag<<3;
  end
  
  lzc #(
    .WIDTH ( 8 )
  ) i_vld_bdirty (
    .in_i    ( bdirty[dirty_ptr] ),
    .cnt_o   ( bdirty_off        ),
    .empty_o (                   )
  );
  
  assign miss_paddr_o = {wbuffer_dirty_mux.wtag, bdirty_off};
  assign miss_id_o    = tx_id;
  
  assign miss_req_o = (|dirty) && free_tx_slots;
  
  
  
  
  assign miss_size_o  = toSize64(bdirty[dirty_ptr]);
  
  assign miss_wdata_o = repData64(wbuffer_dirty_mux.data,
                                  bdirty_off,
                                  miss_size_o[1:0]);
  assign tx_be        = toByteEnable8(bdirty_off,
                                      miss_size_o[1:0]);
  
  fifo_v3 #(
    .FALL_THROUGH ( 1'b0                  ),
    .DATA_WIDTH   ( $clog2(DCACHE_MAX_TX) ),
    .DEPTH        ( DCACHE_MAX_TX         )
  ) i_rtrn_id_fifo (
    .clk_i      ( clk_i            ),
    .rst_ni     ( rst_ni           ),
    .flush_i    ( 1'b0             ),
    .testmode_i ( 1'b0             ),
    .full_o     (                  ),
    .empty_o    ( rtrn_empty       ),
    .usage_o    (                  ),
    .data_i     ( miss_rtrn_id_i   ),
    .push_i     ( miss_rtrn_vld_i  ),
    .data_o     ( rtrn_id          ),
    .pop_i      ( evict            )
  );
  always_comb begin : p_tx_stat
    tx_stat_d = tx_stat_q;
    evict     = 1'b0;
    wr_req_o  = '0;
    
    if ((!rtrn_empty) && wbuffer_q[rtrn_ptr].checked) begin
      
      
      if ((|wr_data_be_o) && (|wbuffer_q[rtrn_ptr].hit_oh)) begin
        wr_req_o = wbuffer_q[rtrn_ptr].hit_oh;
        if (wr_ack_i) begin
          evict    = 1'b1;
          tx_stat_d[rtrn_id].vld = 1'b0;
        end
      end else begin
        evict = 1'b1;
        tx_stat_d[rtrn_id].vld = 1'b0;
      end
    end
    
    if (dirty_rd_en) begin
      tx_stat_d[tx_id].vld = 1'b1;
      tx_stat_d[tx_id].ptr = dirty_ptr;
      tx_stat_d[tx_id].be  = tx_be;
    end
  end
  assign free_tx_slots = |(~tx_vld_o);
  
  rr_arb_tree #(
    .NumIn     (DCACHE_MAX_TX),
    .LockIn    (1'b1),
    .DataWidth (1)
  ) i_tx_id_rr (
    .clk_i  (clk_i       ),
    .rst_ni (rst_ni      ),
    .flush_i('0          ),
    .rr_i   ('0          ),
    .req_i  (~tx_vld_o   ),
    .gnt_o  (            ),
    .data_i ('0          ),
    .gnt_i  (dirty_rd_en ),
    .req_o  (            ),
    .data_o (            ),
    .idx_o  (tx_id       )
  );
  assign rd_tag_d   = rd_paddr>>DCACHE_INDEX_WIDTH;
  
  assign rd_tag_only_o = 1'b1;
  assign rd_paddr   = wbuffer_check_mux.wtag<<3;
  assign rd_req_o   = |tocheck;
  assign rd_tag_o   = rd_tag_q;
  assign rd_idx_o   = rd_paddr[DCACHE_INDEX_WIDTH-1:DCACHE_OFFSET_WIDTH];
  assign rd_off_o   = rd_paddr[DCACHE_OFFSET_WIDTH-1:0];
  assign check_en_d = rd_req_o & rd_ack_i;
  
  assign rtrn_ptr     = tx_stat_q[rtrn_id].ptr;
  
  
  assign wr_data_be_o = tx_stat_q[rtrn_id].be & (~wbuffer_q[rtrn_ptr].dirty);
  assign wr_paddr     = wbuffer_q[rtrn_ptr].wtag<<3;
  assign wr_idx_o     = wr_paddr[DCACHE_INDEX_WIDTH-1:DCACHE_OFFSET_WIDTH];
  assign wr_off_o     = wr_paddr[DCACHE_OFFSET_WIDTH-1:0];
  assign wr_data_o    = wbuffer_q[rtrn_ptr].data;
  logic [DCACHE_WBUF_DEPTH-1:0][DCACHE_CL_IDX_WIDTH-1:0] wtag_comp;
  assign wr_cl_vld_d = wr_cl_vld_i;
  assign wr_cl_idx_d = wr_cl_idx_i;
  for (genvar k=0; k<DCACHE_WBUF_DEPTH; k++) begin : gen_flags
    
    assign debug_paddr[k] = wbuffer_q[k].wtag << 3;
    
    
    
    assign bdirty[k] = (|wbuffer_q[k].txblock) ? '0 : wbuffer_q[k].dirty & wbuffer_q[k].valid;
    assign dirty[k]          = |bdirty[k];
    assign valid[k]          = |wbuffer_q[k].valid;
    assign wbuffer_hit_oh[k] = valid[k] & (wbuffer_q[k].wtag == {req_port_i.address_tag, req_port_i.address_index[DCACHE_INDEX_WIDTH-1:3]});
    
    
    
    assign wtag_comp[k] = wbuffer_q[k].wtag[DCACHE_INDEX_WIDTH-4:DCACHE_OFFSET_WIDTH-3];
    assign inval_hit[k]  = (wr_cl_vld_d & valid[k] & (wtag_comp[k] == wr_cl_idx_d)) |
                           (wr_cl_vld_q & valid[k] & (wtag_comp[k] == wr_cl_idx_q));
    
    assign tocheck[k]       = (~wbuffer_q[k].checked) & valid[k];
  end
  assign wr_ptr     = (|wbuffer_hit_oh) ? hit_ptr : next_ptr;
  assign rdy        = (|wbuffer_hit_oh) | (~full);
  
  lzc #(
    .WIDTH ( DCACHE_WBUF_DEPTH )
  ) i_vld_lzc (
    .in_i    ( ~valid        ),
    .cnt_o   ( next_ptr      ),
    .empty_o ( full          )
  );
  
  lzc #(
    .WIDTH ( DCACHE_WBUF_DEPTH )
  ) i_hit_lzc (
    .in_i    ( wbuffer_hit_oh ),
    .cnt_o   ( hit_ptr        ),
    .empty_o (                )
  );
  
  rr_arb_tree #(
    .NumIn     ( DCACHE_WBUF_DEPTH ),
    .LockIn    ( 1'b1              ),
    .DataType  ( wbuffer_t         )
  ) i_dirty_rr (
    .clk_i  ( clk_i             ),
    .rst_ni ( rst_ni            ),
    .flush_i( '0                ),
    .rr_i   ( '0                ),
    .req_i  ( dirty             ),
    .gnt_o  (                   ),
    .data_i ( wbuffer_q         ),
    .gnt_i  ( dirty_rd_en       ),
    .req_o  (                   ),
    .data_o ( wbuffer_dirty_mux ),
    .idx_o  ( dirty_ptr         )
  );
  
  rr_arb_tree #(
    .NumIn     ( DCACHE_WBUF_DEPTH ),
    .DataType  ( wbuffer_t         )
  ) i_clean_rr (
    .clk_i  ( clk_i             ),
    .rst_ni ( rst_ni            ),
    .flush_i( '0                ),
    .rr_i   ( '0                ),
    .req_i  ( tocheck           ),
    .gnt_o  (                   ),
    .data_i ( wbuffer_q         ),
    .gnt_i  ( check_en_d        ),
    .req_o  (                   ),
    .data_o ( wbuffer_check_mux ),
    .idx_o  ( check_ptr_d       )
  );
  assign req_port_o.data_rvalid = '0;
  assign req_port_o.data_rdata  = '0;
  assign rd_hit_oh_d = rd_hit_oh_i;
 
  logic ni_inside,ni_conflict; 
  assign ni_inside = |ni_pending_q;
  assign ni_conflict = is_ni && ni_inside;
  assign not_ni_o = !ni_inside;
  assign empty_o    = !(|valid);
  
  always_comb begin : p_buffer
    wbuffer_d           = wbuffer_q;
    ni_pending_d        = ni_pending_q;
    dirty_rd_en         = 1'b0;
    req_port_o.data_gnt = 1'b0;
    wbuffer_wren        = 1'b0;
    
    if (check_en_q1) begin
      if (wbuffer_q[check_ptr_q1].valid) begin
        wbuffer_d[check_ptr_q1].checked = 1'b1;
        wbuffer_d[check_ptr_q1].hit_oh = rd_hit_oh_q;
      end
    end
    
    
    for (int k=0; k<DCACHE_WBUF_DEPTH; k++) begin
      if (inval_hit[k]) begin
        wbuffer_d[k].checked = 1'b0;
      end
    end
    
    
    if (evict) begin
      for (int k=0; k<8; k++) begin
        if (tx_stat_q[rtrn_id].be[k]) begin
          wbuffer_d[rtrn_ptr].txblock[k] = 1'b0;
          if (!wbuffer_q[rtrn_ptr].dirty[k]) begin
            wbuffer_d[rtrn_ptr].valid[k] = 1'b0;
            
            
            
          end
        end
      end
      
      if (wbuffer_d[rtrn_ptr].valid == 0) begin
        wbuffer_d[rtrn_ptr].checked = 1'b0;
        ni_pending_d[rtrn_ptr] = 1'b0;
      end
    end
    
    if (miss_req_o && miss_ack_i) begin
      dirty_rd_en = 1'b1;
      for (int k=0; k<8; k++) begin
        if (tx_be[k]) begin
          wbuffer_d[dirty_ptr].dirty[k]   = 1'b0;
          wbuffer_d[dirty_ptr].txblock[k] = 1'b1;
        end
      end
    end
    
    if (req_port_i.data_req && rdy) begin
      
      
      if (!ni_conflict) begin 
        wbuffer_wren              = 1'b1;
        req_port_o.data_gnt       = 1'b1;
        ni_pending_d[wr_ptr]      = is_ni;
        wbuffer_d[wr_ptr].checked = 1'b0;
        wbuffer_d[wr_ptr].wtag    = {req_port_i.address_tag, req_port_i.address_index[DCACHE_INDEX_WIDTH-1:3]};
        
        for (int k=0; k<8; k++) begin
          if (req_port_i.data_be[k]) begin
            wbuffer_d[wr_ptr].valid[k]       = 1'b1;
            wbuffer_d[wr_ptr].dirty[k]       = 1'b1;
            wbuffer_d[wr_ptr].data[k*8 +: 8] = req_port_i.data_wdata[k*8 +: 8];
          end
        end
      end
    end
  end
  always_ff @(posedge clk_i or negedge rst_ni) begin : p_regs
    if (!rst_ni) begin
      wbuffer_q     <= '{default: '0};
      tx_stat_q     <= '{default: '0};
      ni_pending_q  <= '0;
      check_ptr_q   <= '0;
      check_ptr_q1  <= '0;
      check_en_q    <= '0;
      check_en_q1   <= '0;
      rd_tag_q      <= '0;
      rd_hit_oh_q   <= '0;
      wr_cl_vld_q   <= '0;
      wr_cl_idx_q   <= '0;
    end else begin
      wbuffer_q     <= wbuffer_d;
      tx_stat_q     <= tx_stat_d;
      ni_pending_q  <= ni_pending_d;
      check_ptr_q   <= check_ptr_d;
      check_ptr_q1  <= check_ptr_q;
      check_en_q    <= check_en_d;
      check_en_q1   <= check_en_q;
      rd_tag_q      <= rd_tag_d;
      rd_hit_oh_q   <= rd_hit_oh_d;
      wr_cl_vld_q   <= wr_cl_vld_d;
      wr_cl_idx_q   <= wr_cl_idx_d;
    end
  end
endmodule 
module wt_dcache import ariane_pkg::*; import wt_cache_pkg::*; #(
  
  
  parameter logic [CACHE_ID_WIDTH-1:0]   RdAmoTxId          = 1,
  
  parameter ariane_pkg::ariane_cfg_t     ArianeCfg          = ariane_pkg::ArianeDefaultConfig
) (
  input  logic                           clk_i,       
  input  logic                           rst_ni,      
  
  input  logic                           enable_i,    
  input  logic                           flush_i,     
  output logic                           flush_ack_o, 
  output logic                           miss_o,      
  output logic                           wbuffer_empty_o,
  output logic                           wbuffer_not_ni_o,
  
  input  amo_req_t                       amo_req_i,
  output amo_resp_t                      amo_resp_o,
  
  input  dcache_req_i_t [2:0]            req_ports_i,
  output dcache_req_o_t [2:0]            req_ports_o,
  input  logic                           mem_rtrn_vld_i,
  input  dcache_rtrn_t                   mem_rtrn_i,
  output logic                           mem_data_req_o,
  input  logic                           mem_data_ack_i,
  output dcache_req_t                    mem_data_o
);
  
  localparam NumPorts = 3;
  
  logic cache_en;
  
  logic                           wr_cl_vld;
  logic                           wr_cl_nc;
  logic [DCACHE_SET_ASSOC-1:0]    wr_cl_we;
  logic [DCACHE_TAG_WIDTH-1:0]    wr_cl_tag;
  logic [DCACHE_CL_IDX_WIDTH-1:0] wr_cl_idx;
  logic [DCACHE_OFFSET_WIDTH-1:0] wr_cl_off;
  logic [DCACHE_LINE_WIDTH-1:0]   wr_cl_data;
  logic [DCACHE_LINE_WIDTH/8-1:0] wr_cl_data_be;
  logic [DCACHE_SET_ASSOC-1:0]    wr_vld_bits;
  logic [DCACHE_SET_ASSOC-1:0]    wr_req;
  logic                           wr_ack;
  logic [DCACHE_CL_IDX_WIDTH-1:0] wr_idx;
  logic [DCACHE_OFFSET_WIDTH-1:0] wr_off;
  logic [63:0]                    wr_data;
  logic [7:0]                     wr_data_be;
  
  logic [NumPorts-1:0]                          miss_req;
  logic [NumPorts-1:0]                          miss_ack;
  logic [NumPorts-1:0]                          miss_nc;
  logic [NumPorts-1:0]                          miss_we;
  logic [NumPorts-1:0][63:0]                    miss_wdata;
  logic [NumPorts-1:0][riscv::PLEN-1:0]         miss_paddr;
  logic [NumPorts-1:0][DCACHE_SET_ASSOC-1:0]    miss_vld_bits;
  logic [NumPorts-1:0][2:0]                     miss_size;
  logic [NumPorts-1:0][CACHE_ID_WIDTH-1:0]      miss_id;
  logic [NumPorts-1:0]                          miss_replay;
  logic [NumPorts-1:0]                          miss_rtrn_vld;
  logic [CACHE_ID_WIDTH-1:0]                    miss_rtrn_id;
  
  logic [NumPorts-1:0]                          rd_prio;
  logic [NumPorts-1:0]                          rd_tag_only;
  logic [NumPorts-1:0]                          rd_req;
  logic [NumPorts-1:0]                          rd_ack;
  logic [NumPorts-1:0][DCACHE_TAG_WIDTH-1:0]    rd_tag;
  logic [NumPorts-1:0][DCACHE_CL_IDX_WIDTH-1:0] rd_idx;
  logic [NumPorts-1:0][DCACHE_OFFSET_WIDTH-1:0] rd_off;
  logic [63:0]                                  rd_data;
  logic [DCACHE_SET_ASSOC-1:0]                  rd_vld_bits;
  logic [DCACHE_SET_ASSOC-1:0]                  rd_hit_oh;
  
  logic [DCACHE_MAX_TX-1:0][riscv::PLEN-1:0]    tx_paddr;
  logic [DCACHE_MAX_TX-1:0]                     tx_vld;
  
  wbuffer_t [DCACHE_WBUF_DEPTH-1:0]             wbuffer_data;
  wt_dcache_missunit #(
    .Axi64BitCompliant ( ArianeCfg.Axi64BitCompliant ),
    .AmoTxId           ( RdAmoTxId                   ),
    .NumPorts          ( NumPorts                    )
  ) i_wt_dcache_missunit (
    .clk_i              ( clk_i              ),
    .rst_ni             ( rst_ni             ),
    .enable_i           ( enable_i           ),
    .flush_i            ( flush_i            ),
    .flush_ack_o        ( flush_ack_o        ),
    .miss_o             ( miss_o             ),
    .wbuffer_empty_i    ( wbuffer_empty_o    ),
    .cache_en_o         ( cache_en           ),
    
    .amo_req_i          ( amo_req_i          ),
    .amo_resp_o         ( amo_resp_o         ),
    
    .miss_req_i         ( miss_req           ),
    .miss_ack_o         ( miss_ack           ),
    .miss_nc_i          ( miss_nc            ),
    .miss_we_i          ( miss_we            ),
    .miss_wdata_i       ( miss_wdata         ),
    .miss_paddr_i       ( miss_paddr         ),
    .miss_vld_bits_i    ( miss_vld_bits      ),
    .miss_size_i        ( miss_size          ),
    .miss_id_i          ( miss_id            ),
    .miss_replay_o      ( miss_replay        ),
    .miss_rtrn_vld_o    ( miss_rtrn_vld      ),
    .miss_rtrn_id_o     ( miss_rtrn_id       ),
    
    .tx_paddr_i         ( tx_paddr           ),
    .tx_vld_i           ( tx_vld             ),
    
    .wr_cl_vld_o        ( wr_cl_vld          ),
    .wr_cl_nc_o         ( wr_cl_nc           ),
    .wr_cl_we_o         ( wr_cl_we           ),
    .wr_cl_tag_o        ( wr_cl_tag          ),
    .wr_cl_idx_o        ( wr_cl_idx          ),
    .wr_cl_off_o        ( wr_cl_off          ),
    .wr_cl_data_o       ( wr_cl_data         ),
    .wr_cl_data_be_o    ( wr_cl_data_be      ),
    .wr_vld_bits_o      ( wr_vld_bits        ),
    
    .mem_rtrn_vld_i     ( mem_rtrn_vld_i     ),
    .mem_rtrn_i         ( mem_rtrn_i         ),
    .mem_data_req_o     ( mem_data_req_o     ),
    .mem_data_ack_i     ( mem_data_ack_i     ),
    .mem_data_o         ( mem_data_o         )
  );
  
  for(genvar k=0; k<NumPorts-1; k++) begin : gen_rd_ports
    
    assign rd_prio[k] = 1'b1;
    wt_dcache_ctrl #(
      .RdTxId        ( RdAmoTxId     ),
      .ArianeCfg     ( ArianeCfg     )
    ) i_wt_dcache_ctrl (
      .clk_i           ( clk_i             ),
      .rst_ni          ( rst_ni            ),
      .cache_en_i      ( cache_en          ),
      
      .req_port_i      ( req_ports_i   [k] ),
      .req_port_o      ( req_ports_o   [k] ),
      
      .miss_req_o      ( miss_req      [k] ),
      .miss_ack_i      ( miss_ack      [k] ),
      .miss_we_o       ( miss_we       [k] ),
      .miss_wdata_o    ( miss_wdata    [k] ),
      .miss_vld_bits_o ( miss_vld_bits [k] ),
      .miss_paddr_o    ( miss_paddr    [k] ),
      .miss_nc_o       ( miss_nc       [k] ),
      .miss_size_o     ( miss_size     [k] ),
      .miss_id_o       ( miss_id       [k] ),
      .miss_replay_i   ( miss_replay   [k] ),
      .miss_rtrn_vld_i ( miss_rtrn_vld [k] ),
      
      .wr_cl_vld_i     ( wr_cl_vld         ),
      
      .rd_tag_o        ( rd_tag        [k] ),
      .rd_idx_o        ( rd_idx        [k] ),
      .rd_off_o        ( rd_off        [k] ),
      .rd_req_o        ( rd_req        [k] ),
      .rd_tag_only_o   ( rd_tag_only   [k] ),
      .rd_ack_i        ( rd_ack        [k] ),
      .rd_data_i       ( rd_data           ),
      .rd_vld_bits_i   ( rd_vld_bits       ),
      .rd_hit_oh_i     ( rd_hit_oh         )
    );
  end
  
  assign rd_prio[2] = 1'b0;
  wt_dcache_wbuffer #(
    .ArianeCfg     ( ArianeCfg     )
  ) i_wt_dcache_wbuffer (
    .clk_i           ( clk_i               ),
    .rst_ni          ( rst_ni              ),
    .empty_o         ( wbuffer_empty_o     ),
    .not_ni_o        ( wbuffer_not_ni_o    ),
    
    .cache_en_i      ( cache_en            ),
    
    
    .req_port_i      ( req_ports_i   [2]   ),
    .req_port_o      ( req_ports_o   [2]   ),
    
    .miss_req_o      ( miss_req      [2]   ),
    .miss_ack_i      ( miss_ack      [2]   ),
    .miss_we_o       ( miss_we       [2]   ),
    .miss_wdata_o    ( miss_wdata    [2]   ),
    .miss_vld_bits_o ( miss_vld_bits [2]   ),
    .miss_paddr_o    ( miss_paddr    [2]   ),
    .miss_nc_o       ( miss_nc       [2]   ),
    .miss_size_o     ( miss_size     [2]   ),
    .miss_id_o       ( miss_id       [2]   ),
    .miss_rtrn_vld_i ( miss_rtrn_vld [2]   ),
    .miss_rtrn_id_i  ( miss_rtrn_id        ),
    
    .rd_tag_o        ( rd_tag        [2]   ),
    .rd_idx_o        ( rd_idx        [2]   ),
    .rd_off_o        ( rd_off        [2]   ),
    .rd_req_o        ( rd_req        [2]   ),
    .rd_tag_only_o   ( rd_tag_only   [2]   ),
    .rd_ack_i        ( rd_ack        [2]   ),
    .rd_data_i       ( rd_data             ),
    .rd_vld_bits_i   ( rd_vld_bits         ),
    .rd_hit_oh_i     ( rd_hit_oh           ),
     
    .wr_cl_vld_i     ( wr_cl_vld           ),
    .wr_cl_idx_i     ( wr_cl_idx           ),
    
    .wr_req_o        ( wr_req              ),
    .wr_ack_i        ( wr_ack              ),
    .wr_idx_o        ( wr_idx              ),
    .wr_off_o        ( wr_off              ),
    .wr_data_o       ( wr_data             ),
    .wr_data_be_o    ( wr_data_be          ),
    
    .wbuffer_data_o  ( wbuffer_data        ),
    .tx_paddr_o      ( tx_paddr            ),
    .tx_vld_o        ( tx_vld              )
  );
  wt_dcache_mem #(
    .Axi64BitCompliant ( ArianeCfg.Axi64BitCompliant ),
    .NumPorts          ( NumPorts                    )
  ) i_wt_dcache_mem (
    .clk_i             ( clk_i              ),
    .rst_ni            ( rst_ni             ),
    
    .rd_prio_i         ( rd_prio            ),
    .rd_tag_i          ( rd_tag             ),
    .rd_idx_i          ( rd_idx             ),
    .rd_off_i          ( rd_off             ),
    .rd_req_i          ( rd_req             ),
    .rd_tag_only_i     ( rd_tag_only        ),
    .rd_ack_o          ( rd_ack             ),
    .rd_vld_bits_o     ( rd_vld_bits        ),
    .rd_hit_oh_o       ( rd_hit_oh          ),
    .rd_data_o         ( rd_data            ),
    
    .wr_cl_vld_i       ( wr_cl_vld          ),
    .wr_cl_nc_i        ( wr_cl_nc           ),
    .wr_cl_we_i        ( wr_cl_we           ),
    .wr_cl_tag_i       ( wr_cl_tag          ),
    .wr_cl_idx_i       ( wr_cl_idx          ),
    .wr_cl_off_i       ( wr_cl_off          ),
    .wr_cl_data_i      ( wr_cl_data         ),
    .wr_cl_data_be_i   ( wr_cl_data_be      ),
    .wr_vld_bits_i     ( wr_vld_bits        ),
    
    .wr_req_i          ( wr_req             ),
    .wr_ack_o          ( wr_ack             ),
    .wr_idx_i          ( wr_idx             ),
    .wr_off_i          ( wr_off             ),
    .wr_data_i         ( wr_data            ),
    .wr_data_be_i      ( wr_data_be         ),
    
    .wbuffer_data_i    ( wbuffer_data       )
  );
endmodule 
module cva6_icache import ariane_pkg::*; import wt_cache_pkg::*; #(
  parameter logic [CACHE_ID_WIDTH-1:0]  RdTxId             = 0,                                  
  parameter ariane_pkg::ariane_cfg_t    ArianeCfg          = ariane_pkg::ArianeDefaultConfig     
) (
  input  logic                      clk_i,
  input  logic                      rst_ni,
  input  logic                      flush_i,              
  input  logic                      en_i,                 
  output logic                      miss_o,               
  
  input  icache_areq_i_t            areq_i,
  output icache_areq_o_t            areq_o,
  
  input  icache_dreq_i_t            dreq_i,
  output icache_dreq_o_t            dreq_o,
  
  input  logic                      mem_rtrn_vld_i,
  input  icache_rtrn_t              mem_rtrn_i,
  output logic                      mem_data_req_o,
  input  logic                      mem_data_ack_i,
  output icache_req_t               mem_data_o
);
  
  logic                                 cache_en_d, cache_en_q;       
  logic [riscv::VLEN-1:0]               vaddr_d, vaddr_q;
  logic                                 paddr_is_nc;                  
  logic [ICACHE_SET_ASSOC-1:0]          cl_hit;                       
  logic                                 cache_rden;                   
  logic                                 cache_wren;                   
  logic                                 cmp_en_d, cmp_en_q;           
  logic                                 flush_d, flush_q;             
  
  logic                                 update_lfsr;                  
  logic [$clog2(ICACHE_SET_ASSOC)-1:0]  inv_way;                      
  logic [$clog2(ICACHE_SET_ASSOC)-1:0]  rnd_way;                      
  logic [$clog2(ICACHE_SET_ASSOC)-1:0]  repl_way;                     
  logic [ICACHE_SET_ASSOC-1:0]          repl_way_oh_d, repl_way_oh_q; 
  logic                                 all_ways_valid;               
  
  logic                                 inv_en;                       
  logic                                 inv_d, inv_q;                 
  logic                                 flush_en, flush_done;         
  logic [ICACHE_CL_IDX_WIDTH-1:0]       flush_cnt_d, flush_cnt_q;     
  
  logic                                 cl_we;                        
  logic [ICACHE_SET_ASSOC-1:0]          cl_req;                       
  logic [ICACHE_CL_IDX_WIDTH-1:0]       cl_index;                     
  logic [ICACHE_OFFSET_WIDTH-1:0]       cl_offset_d, cl_offset_q;     
  logic [ICACHE_TAG_WIDTH-1:0]          cl_tag_d, cl_tag_q;           
  logic [ICACHE_TAG_WIDTH-1:0]          cl_tag_rdata [ICACHE_SET_ASSOC-1:0]; 
  logic [ICACHE_LINE_WIDTH-1:0]         cl_rdata     [ICACHE_SET_ASSOC-1:0]; 
  logic [ICACHE_SET_ASSOC-1:0][FETCH_WIDTH-1:0]cl_sel;                
  logic [ICACHE_SET_ASSOC-1:0]          vld_req;                      
  logic                                 vld_we;                       
  logic [ICACHE_SET_ASSOC-1:0]          vld_wdata;                    
  logic [ICACHE_SET_ASSOC-1:0]          vld_rdata;                    
  logic [ICACHE_CL_IDX_WIDTH-1:0]       vld_addr;                     
  
  typedef enum logic[2:0] {FLUSH, IDLE, READ, MISS, KILL_ATRANS, KILL_MISS} state_e;
  state_e state_d, state_q;
  
  assign cl_tag_d  = (areq_i.fetch_valid) ? areq_i.fetch_paddr[ICACHE_TAG_WIDTH+ICACHE_INDEX_WIDTH-1:ICACHE_INDEX_WIDTH] : cl_tag_q;
  
  assign paddr_is_nc = (~cache_en_q) | (~ariane_pkg::is_inside_cacheable_regions(ArianeCfg, {{{64-riscv::PLEN}{1'b0}}, cl_tag_d, {ICACHE_INDEX_WIDTH{1'b0}}}));
  
  assign dreq_o.ex = areq_i.fetch_exception;
  
  
  assign vaddr_d = (dreq_o.ready & dreq_i.req) ? dreq_i.vaddr : vaddr_q;
  assign areq_o.fetch_vaddr = {vaddr_q>>2, 2'b0};
  
  assign cl_index    = vaddr_d[ICACHE_INDEX_WIDTH-1:ICACHE_OFFSET_WIDTH];
  if (ArianeCfg.Axi64BitCompliant) begin : gen_axi_offset
    
    assign cl_offset_d = ( dreq_o.ready & dreq_i.req)      ? {dreq_i.vaddr>>2, 2'b0} :
                         ( paddr_is_nc  & mem_data_req_o ) ? cl_offset_q[2]<<2 : 
                                                             cl_offset_q;
    
    assign mem_data_o.paddr = (paddr_is_nc) ? {cl_tag_d, vaddr_q[ICACHE_INDEX_WIDTH-1:3], 3'b0} :                                         
                                              {cl_tag_d, vaddr_q[ICACHE_INDEX_WIDTH-1:ICACHE_OFFSET_WIDTH], {ICACHE_OFFSET_WIDTH{1'b0}}}; 
end else begin : gen_piton_offset
    
    
    assign cl_offset_d = ( dreq_o.ready & dreq_i.req)      ? {dreq_i.vaddr>>2, 2'b0} :
                                                             cl_offset_q;
    
    assign mem_data_o.paddr = (paddr_is_nc) ? {cl_tag_d, vaddr_q[ICACHE_INDEX_WIDTH-1:2], 2'b0} :                                         
                                              {cl_tag_d, vaddr_q[ICACHE_INDEX_WIDTH-1:ICACHE_OFFSET_WIDTH], {ICACHE_OFFSET_WIDTH{1'b0}}}; 
  end
  assign mem_data_o.tid   = RdTxId;
  assign mem_data_o.nc    = paddr_is_nc;
  
  assign mem_data_o.way   = repl_way;
  assign dreq_o.vaddr     = vaddr_q;
  
  assign inv_d = inv_en;
  logic addr_ni;
  assign addr_ni = is_inside_nonidempotent_regions(ArianeCfg, areq_i.fetch_paddr);
  always_comb begin : p_fsm
    
    state_d      = state_q;
    cache_en_d   = cache_en_q & en_i;
    flush_en     = 1'b0;
    cmp_en_d     = 1'b0;
    cache_rden   = 1'b0;
    cache_wren   = 1'b0;
    inv_en       = 1'b0;
    flush_d      = flush_q | flush_i; 
    
    dreq_o.ready     = 1'b0;
    areq_o.fetch_req = 1'b0;
    dreq_o.valid     = 1'b0;
    mem_data_req_o   = 1'b0;
    
    miss_o           = 1'b0;
    
    
    
    
    
    if (mem_rtrn_vld_i && mem_rtrn_i.rtype == ICACHE_INV_REQ) begin
      inv_en = 1'b1;
    end
    unique case (state_q)
      
      
      FLUSH: begin
          flush_en = 1'b1;
        if (flush_done) begin
          state_d = IDLE;
          flush_d = 1'b0;
          
          cache_en_d = en_i;
        end
      end
      
      
      IDLE: begin
          
          cmp_en_d = cache_en_q;
          
          if (flush_d || (en_i && !cache_en_q)) begin
            state_d    = FLUSH;
          
          end else begin
            
            if (!mem_rtrn_vld_i) begin
              dreq_o.ready = 1'b1;
              
              if (dreq_i.req) begin
                cache_rden       = 1'b1;
                state_d          = READ;
              end
            end
            if (dreq_i.kill_s1) begin
              state_d = IDLE;
            end
          end
      end
      
      
      
      
      
      
      READ: begin
          areq_o.fetch_req = '1;
          
          cmp_en_d    = cache_en_q;
          
          cache_rden  = cache_en_q;
          if (areq_i.fetch_valid && (!dreq_i.spec || !addr_ni) ) begin
            
            if (flush_d) begin
              state_d  = IDLE;
            
            end else if (((|cl_hit && cache_en_q) || areq_i.fetch_exception.valid) && !inv_q) begin
              dreq_o.valid     = ~dreq_i.kill_s2;
              state_d          = IDLE;
              
              
              
              if (!mem_rtrn_vld_i) begin
                dreq_o.ready     = 1'b1;
                if (dreq_i.req) begin
                  state_d          = READ;
                end
              end
              
              
              if (dreq_i.kill_s1) begin
                state_d = IDLE;
              end
            
            end else if (dreq_i.kill_s2) begin
              state_d = IDLE;
            end else if (!inv_q) begin
              cmp_en_d = 1'b0;
              
              
              
              mem_data_req_o = 1'b1;
              if (mem_data_ack_i) begin
                miss_o         = ~paddr_is_nc;
                state_d        = MISS;
              end
            end
          
          end else if (dreq_i.kill_s2 || flush_d) begin
            state_d  = KILL_ATRANS;
          end
      end
      
      
      
      
      MISS: begin
        
        
        if (mem_rtrn_vld_i && mem_rtrn_i.rtype == ICACHE_IFILL_ACK) begin
          state_d      = IDLE;
          
          if (!(dreq_i.kill_s2 || flush_d)) begin
            dreq_o.valid = 1'b1;
            
            cache_wren   = ~paddr_is_nc;
          end
        
        end else if (dreq_i.kill_s2 || flush_d) begin
          state_d  = KILL_MISS;
        end
      end
      
      
      
      
      KILL_ATRANS: begin
        areq_o.fetch_req = '1;
        if (areq_i.fetch_valid) begin
          state_d      = IDLE;
        end
      end
      
      
      
      
      KILL_MISS: begin
        if (mem_rtrn_vld_i && mem_rtrn_i.rtype == ICACHE_IFILL_ACK) begin
          state_d      = IDLE;
        end
      end
      default: begin
        
        state_d = FLUSH;
      end
    endcase 
  end
  
  
  
  
  assign flush_cnt_d = (flush_done) ? '0               :
                       (flush_en)   ?  flush_cnt_q + 1 :
                                       flush_cnt_q;
  assign flush_done  = (flush_cnt_q==(ICACHE_NUM_WORDS-1));
  
  
  assign vld_addr = (flush_en)       ? flush_cnt_q        :
                    (inv_en)         ? mem_rtrn_i.inv.idx[ICACHE_INDEX_WIDTH-1:ICACHE_OFFSET_WIDTH] :
                                       cl_index;
  assign vld_req  = (flush_en || cache_rden)        ? '1                                    :
                    (mem_rtrn_i.inv.all && inv_en)  ? '1                                    :
                    (mem_rtrn_i.inv.vld && inv_en)  ? icache_way_bin2oh(mem_rtrn_i.inv.way) :
                                                      repl_way_oh_q;
  assign vld_wdata = (cache_wren) ? '1 : '0;
  assign vld_we    = (cache_wren | inv_en | flush_en);
  
  
  assign update_lfsr   = cache_wren & all_ways_valid;
  assign repl_way      = (all_ways_valid) ? rnd_way : inv_way;
  assign repl_way_oh_d = (cmp_en_q) ? icache_way_bin2oh(repl_way) : repl_way_oh_q;
  
  assign cl_req   = (cache_rden) ? '1            :
                    (cache_wren) ? repl_way_oh_q :
                                   '0;
  assign cl_we    = cache_wren;
  
  lzc #(
    .WIDTH ( ICACHE_SET_ASSOC )
  ) i_lzc (
    .in_i    ( ~vld_rdata     ),
    .cnt_o   ( inv_way        ),
    .empty_o ( all_ways_valid )
  );
  
  lfsr #(
    .LfsrWidth  ( ariane_pkg::ICACHE_SET_ASSOC        ),
    .OutWidth   ( $clog2(ariane_pkg::ICACHE_SET_ASSOC))
  ) i_lfsr (
    .clk_i          ( clk_i       ),
    .rst_ni         ( rst_ni      ),
    .en_i           ( update_lfsr ),
    .out_o          ( rnd_way     )
  );
  logic [$clog2(ICACHE_SET_ASSOC)-1:0] hit_idx;
  for (genvar i=0;i<ICACHE_SET_ASSOC;i++) begin : gen_tag_cmpsel
    assign cl_hit[i] = (cl_tag_rdata[i] == cl_tag_d) & vld_rdata[i];
    assign cl_sel[i] = cl_rdata[i][{cl_offset_q,3'b0} +: FETCH_WIDTH];
  end
  lzc #(
    .WIDTH ( ICACHE_SET_ASSOC )
  ) i_lzc_hit (
    .in_i    ( cl_hit  ),
    .cnt_o   ( hit_idx ),
    .empty_o (         )
  );
  assign dreq_o.data = (cmp_en_q) ? cl_sel[hit_idx] :
                                    mem_rtrn_i.data[{cl_offset_q,3'b0} +: FETCH_WIDTH];
  logic [ICACHE_TAG_WIDTH:0] cl_tag_valid_rdata [ICACHE_SET_ASSOC-1:0];
  for (genvar i = 0; i < ICACHE_SET_ASSOC; i++) begin : gen_sram
    
    sram #(
      
      .DATA_WIDTH ( ICACHE_TAG_WIDTH+1 ),
      .NUM_WORDS  ( ICACHE_NUM_WORDS   )
    ) tag_sram (
      .clk_i     ( clk_i                    ),
      .rst_ni    ( rst_ni                   ),
      .req_i     ( vld_req[i]               ),
      .we_i      ( vld_we                   ),
      .addr_i    ( vld_addr                 ),
      
      
      .wdata_i   ( {vld_wdata[i], cl_tag_q} ),
      .be_i      ( '1                       ),
      .rdata_o   ( cl_tag_valid_rdata[i]    )
    );
    assign cl_tag_rdata[i] = cl_tag_valid_rdata[i][ICACHE_TAG_WIDTH-1:0];
    assign vld_rdata[i]    = cl_tag_valid_rdata[i][ICACHE_TAG_WIDTH];
    
    sram #(
      .DATA_WIDTH ( ICACHE_LINE_WIDTH ),
      .NUM_WORDS  ( ICACHE_NUM_WORDS  )
    ) data_sram (
      .clk_i     ( clk_i               ),
      .rst_ni    ( rst_ni              ),
      .req_i     ( cl_req[i]           ),
      .we_i      ( cl_we               ),
      .addr_i    ( cl_index            ),
      .wdata_i   ( mem_rtrn_i.data     ),
      .be_i      ( '1                  ),
      .rdata_o   ( cl_rdata[i]         )
    );
  end
  always_ff @(posedge clk_i or negedge rst_ni) begin : p_regs
    if(!rst_ni) begin
      cl_tag_q      <= '0;
      flush_cnt_q   <= '0;
      vaddr_q       <= '0;
      cmp_en_q      <= '0;
      cache_en_q    <= '0;
      flush_q       <= '0;
      state_q       <= FLUSH;
      cl_offset_q   <= '0;
      repl_way_oh_q <= '0;
      inv_q         <= '0;
    end else begin
      cl_tag_q      <= cl_tag_d;
      flush_cnt_q   <= flush_cnt_d;
      vaddr_q       <= vaddr_d;
      cmp_en_q      <= cmp_en_d;
      cache_en_q    <= cache_en_d;
      flush_q       <= flush_d;
      state_q       <= state_d;
      cl_offset_q   <= cl_offset_d;
      repl_way_oh_q <= repl_way_oh_d;
      inv_q         <= inv_d;
    end
  end
endmodule 
module wt_l15_adapter import ariane_pkg::*; import wt_cache_pkg::*; #(
  parameter bit          SwapEndianess = 1
) (
  input logic                  clk_i,
  input logic                  rst_ni,
  
  input  logic                 icache_data_req_i,
  output logic                 icache_data_ack_o,
  input  icache_req_t          icache_data_i,
  
  output logic                 icache_rtrn_vld_o,
  output icache_rtrn_t         icache_rtrn_o,
  
  input  logic                 dcache_data_req_i,
  output logic                 dcache_data_ack_o,
  input  dcache_req_t          dcache_data_i,
  
  output logic                 dcache_rtrn_vld_o,
  output dcache_rtrn_t         dcache_rtrn_o,
  
  output l15_req_t             l15_req_o,
  input  l15_rtrn_t            l15_rtrn_i
);
icache_req_t icache_data;
logic icache_data_full, icache_data_empty;
dcache_req_t dcache_data;
logic dcache_data_full, dcache_data_empty;
logic [1:0] arb_req, arb_ack;
logic       arb_idx;
logic rtrn_fifo_empty, rtrn_fifo_full, rtrn_fifo_pop;
l15_rtrn_t rtrn_fifo_data;
  
  
  
  
  
  
  
  
  
  
  
  assign icache_data_ack_o  = icache_data_req_i & ~icache_data_full;
  assign dcache_data_ack_o  = dcache_data_req_i & ~dcache_data_full;
  
  assign l15_req_o.l15_nc                   = (arb_idx)        ? dcache_data.nc    : icache_data.nc;
  
  assign l15_req_o.l15_size                 = (arb_idx)        ? dcache_data.size  :
                                              (icache_data.nc) ? 3'b010            : 3'b111;
  assign l15_req_o.l15_threadid             = (arb_idx)        ? dcache_data.tid   : icache_data.tid;
  assign l15_req_o.l15_prefetch             = '0; 
  assign l15_req_o.l15_invalidate_cacheline = '0; 
  assign l15_req_o.l15_blockstore           = '0; 
  assign l15_req_o.l15_blockinitstore       = '0; 
  assign l15_req_o.l15_l1rplway             = (arb_idx) ? dcache_data.way   : icache_data.way;
  assign l15_req_o.l15_address              = (arb_idx) ? dcache_data.paddr :
                                                          icache_data.paddr;
  assign l15_req_o.l15_data_next_entry      = '0; 
  assign l15_req_o.l15_csm_data             = '0; 
  assign l15_req_o.l15_amo_op               = dcache_data.amo_op;
  
  if (SwapEndianess) assign l15_req_o.l15_data = swendian64(dcache_data.data);
  else               assign l15_req_o.l15_data = dcache_data.data;
  
  rrarbiter #(
    .NUM_REQ(2),
    .LOCK_IN(1)
  ) i_rrarbiter (
    .clk_i  ( clk_i                ),
    .rst_ni ( rst_ni               ),
    .flush_i( '0                   ),
    .en_i   ( l15_rtrn_i.l15_ack   ),
    .req_i  ( arb_req              ),
    .ack_o  ( arb_ack              ),
    .vld_o  (                      ),
    .idx_o  ( arb_idx              )
  );
  assign arb_req           = {~dcache_data_empty, ~icache_data_empty};
  assign l15_req_o.l15_val = (|arb_req);
  
  always_comb begin : p_req
    l15_req_o.l15_rqtype = L15_LOAD_RQ;
    unique case (arb_idx)
      0: begin
        l15_req_o.l15_rqtype = L15_IMISS_RQ;
      end
      1: begin
        unique case (dcache_data.rtype)
          DCACHE_STORE_REQ: begin
            l15_req_o.l15_rqtype = L15_STORE_RQ;
          end
          DCACHE_LOAD_REQ: begin
            l15_req_o.l15_rqtype = L15_LOAD_RQ;
          end
          DCACHE_ATOMIC_REQ: begin
            l15_req_o.l15_rqtype = L15_ATOMIC_RQ;
          end
          
          
          
          default: begin
            ;
          end
        endcase 
      end
      default: begin
        ;
      end
    endcase
  end 
  fifo_v2 #(
    .dtype       (  icache_req_t            ),
    .DEPTH       (  ADAPTER_REQ_FIFO_DEPTH  )
    ) i_icache_data_fifo (
    .clk_i       (  clk_i                   ),
    .rst_ni      (  rst_ni                  ),
    .flush_i     (  1'b0                    ),
    .testmode_i  (  1'b0                    ),
    .full_o      (  icache_data_full        ),
    .empty_o     (  icache_data_empty       ),
    .alm_full_o  (                          ),
    .alm_empty_o (                          ),
    .data_i      (  icache_data_i           ),
    .push_i      (  icache_data_ack_o       ),
    .data_o      (  icache_data             ),
    .pop_i       (  arb_ack[0]              )
  );
  fifo_v2 #(
    .dtype       (  dcache_req_t            ),
    .DEPTH       (  ADAPTER_REQ_FIFO_DEPTH  )
    ) i_dcache_data_fifo (
    .clk_i       (  clk_i                   ),
    .rst_ni      (  rst_ni                  ),
    .flush_i     (  1'b0                    ),
    .testmode_i  (  1'b0                    ),
    .full_o      (  dcache_data_full        ),
    .empty_o     (  dcache_data_empty       ),
    .alm_full_o  (                          ),
    .alm_empty_o (                          ),
    .data_i      (  dcache_data_i           ),
    .push_i      (  dcache_data_ack_o       ),
    .data_o      (  dcache_data             ),
    .pop_i       (  arb_ack[1]              )
  );
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  assign l15_req_o.l15_req_ack = l15_rtrn_i.l15_val & ~rtrn_fifo_full;
  
  assign rtrn_fifo_pop = ~rtrn_fifo_empty;
  
  always_comb begin : p_rtrn_logic
    icache_rtrn_o.rtype = ICACHE_IFILL_ACK;
    dcache_rtrn_o.rtype = DCACHE_LOAD_ACK;
    icache_rtrn_vld_o   = 1'b0;
    dcache_rtrn_vld_o   = 1'b0;
    if(!rtrn_fifo_empty) begin
      unique case (rtrn_fifo_data.l15_returntype)
        L15_LOAD_RET:  begin
          dcache_rtrn_o.rtype = DCACHE_LOAD_ACK;
          dcache_rtrn_vld_o   = 1'b1;
        end
        L15_ST_ACK:    begin
          dcache_rtrn_o.rtype = DCACHE_STORE_ACK;
          dcache_rtrn_vld_o   = 1'b1;
        end
        L15_IFILL_RET: begin
          icache_rtrn_o.rtype = ICACHE_IFILL_ACK;
          icache_rtrn_vld_o   = 1'b1;
        end
        L15_EVICT_REQ: begin
          icache_rtrn_o.rtype = ICACHE_INV_REQ;
          dcache_rtrn_o.rtype = DCACHE_INV_REQ;
          icache_rtrn_vld_o   = icache_rtrn_o.inv.vld | icache_rtrn_o.inv.all;
          dcache_rtrn_vld_o   = dcache_rtrn_o.inv.vld | dcache_rtrn_o.inv.all;
        end
        L15_CPX_RESTYPE_ATOMIC_RES: begin
          dcache_rtrn_o.rtype = DCACHE_ATOMIC_ACK;
          dcache_rtrn_vld_o   = 1'b1;
        end
        
        
        
        
        default: begin
        ;
        end
      endcase 
    end
  end
  
  if (SwapEndianess) begin : gen_swap
    assign dcache_rtrn_o.data = { swendian64(rtrn_fifo_data.l15_data_1),
                                  swendian64(rtrn_fifo_data.l15_data_0) };
    assign icache_rtrn_o.data = { swendian64(rtrn_fifo_data.l15_data_3),
                                  swendian64(rtrn_fifo_data.l15_data_2),
                                  swendian64(rtrn_fifo_data.l15_data_1),
                                  swendian64(rtrn_fifo_data.l15_data_0) };
  end else begin : gen_no_swap
    assign dcache_rtrn_o.data = { rtrn_fifo_data.l15_data_1,
                                  rtrn_fifo_data.l15_data_0 };
    assign icache_rtrn_o.data = { rtrn_fifo_data.l15_data_3,
                                  rtrn_fifo_data.l15_data_2,
                                  rtrn_fifo_data.l15_data_1,
                                  rtrn_fifo_data.l15_data_0 };
  end
  
  assign icache_rtrn_o.tid      = rtrn_fifo_data.l15_threadid;
  assign dcache_rtrn_o.tid      = rtrn_fifo_data.l15_threadid;
  
  assign icache_rtrn_o.inv.idx  = {rtrn_fifo_data.l15_inval_address_15_4, 4'b0000};
  assign icache_rtrn_o.inv.way  = rtrn_fifo_data.l15_inval_way;
  assign icache_rtrn_o.inv.vld  = rtrn_fifo_data.l15_inval_icache_inval;
  assign icache_rtrn_o.inv.all  = rtrn_fifo_data.l15_inval_icache_all_way;
  assign dcache_rtrn_o.inv.idx  = {rtrn_fifo_data.l15_inval_address_15_4, 4'b0000};
  assign dcache_rtrn_o.inv.way  = rtrn_fifo_data.l15_inval_way;
  assign dcache_rtrn_o.inv.vld  = rtrn_fifo_data.l15_inval_dcache_inval;
  assign dcache_rtrn_o.inv.all  = rtrn_fifo_data.l15_inval_dcache_all_way;
  fifo_v2 #(
    .dtype       (  l15_rtrn_t               ),
    .DEPTH       (  ADAPTER_RTRN_FIFO_DEPTH  )
  ) i_rtrn_fifo (
    .clk_i       (  clk_i                    ),
    .rst_ni      (  rst_ni                   ),
    .flush_i     (  1'b0                     ),
    .testmode_i  (  1'b0                     ),
    .full_o      (  rtrn_fifo_full           ),
    .empty_o     (  rtrn_fifo_empty          ),
    .alm_full_o  (                           ),
    .alm_empty_o (                           ),
    .data_i      (  l15_rtrn_i               ),
    .push_i      (  l15_req_o.l15_req_ack    ),
    .data_o      (  rtrn_fifo_data           ),
    .pop_i       (  rtrn_fifo_pop            )
  );
endmodule 
module wt_cache_subsystem import ariane_pkg::*; import wt_cache_pkg::*; #(
  parameter ariane_pkg::ariane_cfg_t ArianeCfg       = ariane_pkg::ArianeDefaultConfig  
) (
  input logic                            clk_i,
  input logic                            rst_ni,
  
  input  logic                           icache_en_i,            
  input  logic                           icache_flush_i,         
  output logic                           icache_miss_o,          
  
  input  icache_areq_i_t                 icache_areq_i,          
  output icache_areq_o_t                 icache_areq_o,
  
  input  icache_dreq_i_t                 icache_dreq_i,          
  output icache_dreq_o_t                 icache_dreq_o,
  
  
  input  logic                           dcache_enable_i,        
  input  logic                           dcache_flush_i,         
  output logic                           dcache_flush_ack_o,     
  output logic                           dcache_miss_o,          
  
  input amo_req_t                        dcache_amo_req_i,
  output amo_resp_t                      dcache_amo_resp_o,
  
  input  dcache_req_i_t   [2:0]          dcache_req_ports_i,     
  output dcache_req_o_t   [2:0]          dcache_req_ports_o,     
  
  output logic                           wbuffer_empty_o,
  output logic                           wbuffer_not_ni_o,
  
  output l15_req_t                       l15_req_o,
  input  l15_rtrn_t                      l15_rtrn_i
  
);
  logic icache_adapter_data_req, adapter_icache_data_ack, adapter_icache_rtrn_vld;
  wt_cache_pkg::icache_req_t  icache_adapter;
  wt_cache_pkg::icache_rtrn_t adapter_icache;
  logic dcache_adapter_data_req, adapter_dcache_data_ack, adapter_dcache_rtrn_vld;
  wt_cache_pkg::dcache_req_t  dcache_adapter;
  wt_cache_pkg::dcache_rtrn_t adapter_dcache;
  cva6_icache #(
    
    .RdTxId             ( 0             ),
    .ArianeCfg          ( ArianeCfg     )
  ) i_cva6_icache (
    .clk_i              ( clk_i                   ),
    .rst_ni             ( rst_ni                  ),
    .flush_i            ( icache_flush_i          ),
    .en_i               ( icache_en_i             ),
    .miss_o             ( icache_miss_o           ),
    .areq_i             ( icache_areq_i           ),
    .areq_o             ( icache_areq_o           ),
    .dreq_i             ( icache_dreq_i           ),
    .dreq_o             ( icache_dreq_o           ),
    .mem_rtrn_vld_i     ( adapter_icache_rtrn_vld ),
    .mem_rtrn_i         ( adapter_icache          ),
    .mem_data_req_o     ( icache_adapter_data_req ),
    .mem_data_ack_i     ( adapter_icache_data_ack ),
    .mem_data_o         ( icache_adapter          )
  );
  
  
  
  
  wt_dcache #(
    
    
    .RdAmoTxId       ( 1             ),
    .ArianeCfg       ( ArianeCfg     )
  ) i_wt_dcache (
    .clk_i           ( clk_i                   ),
    .rst_ni          ( rst_ni                  ),
    .enable_i        ( dcache_enable_i         ),
    .flush_i         ( dcache_flush_i          ),
    .flush_ack_o     ( dcache_flush_ack_o      ),
    .miss_o          ( dcache_miss_o           ),
    .wbuffer_empty_o ( wbuffer_empty_o         ),
    .wbuffer_not_ni_o ( wbuffer_not_ni_o       ),
    .amo_req_i       ( dcache_amo_req_i        ),
    .amo_resp_o      ( dcache_amo_resp_o       ),
    .req_ports_i     ( dcache_req_ports_i      ),
    .req_ports_o     ( dcache_req_ports_o      ),
    .mem_rtrn_vld_i  ( adapter_dcache_rtrn_vld ),
    .mem_rtrn_i      ( adapter_dcache          ),
    .mem_data_req_o  ( dcache_adapter_data_req ),
    .mem_data_ack_i  ( adapter_dcache_data_ack ),
    .mem_data_o      ( dcache_adapter          )
  );
  wt_l15_adapter #(
    .SwapEndianess   ( ArianeCfg.SwapEndianess )
  ) i_adapter (
    .clk_i              ( clk_i                   ),
    .rst_ni             ( rst_ni                  ),
    .icache_data_req_i  ( icache_adapter_data_req ),
    .icache_data_ack_o  ( adapter_icache_data_ack ),
    .icache_data_i      ( icache_adapter          ),
    .icache_rtrn_vld_o  ( adapter_icache_rtrn_vld ),
    .icache_rtrn_o      ( adapter_icache          ),
    .dcache_data_req_i  ( dcache_adapter_data_req ),
    .dcache_data_ack_o  ( adapter_dcache_data_ack ),
    .dcache_data_i      ( dcache_adapter          ),
    .dcache_rtrn_vld_o  ( adapter_dcache_rtrn_vld ),
    .dcache_rtrn_o      ( adapter_dcache          ),
    .l15_req_o          ( l15_req_o               ),
    .l15_rtrn_i         ( l15_rtrn_i              )
  );
endmodule 
module clint #(
    parameter int unsigned AXI_ADDR_WIDTH = 64,
    parameter int unsigned AXI_DATA_WIDTH = 64,
    parameter int unsigned AXI_ID_WIDTH   = 10,
    parameter int unsigned NR_CORES       = 1 
) (
    input  logic                clk_i,       
    input  logic                rst_ni,      
    input  logic                testmode_i,
    input  ariane_axi::req_t    axi_req_i,
    output ariane_axi::resp_t   axi_resp_o,
    input  logic                rtc_i,       
    output logic [NR_CORES-1:0] timer_irq_o, 
    output logic [NR_CORES-1:0] ipi_o        
);
    
    localparam logic [15:0] MSIP_BASE     = 16'h0;
    localparam logic [15:0] MTIMECMP_BASE = 16'h4000;
    localparam logic [15:0] MTIME_BASE    = 16'hbff8;
    localparam AddrSelWidth = (NR_CORES == 1) ? 1 : $clog2(NR_CORES);
    
    logic [AXI_ADDR_WIDTH-1:0] address;
    logic                      en;
    logic                      we;
    logic [63:0] wdata;
    logic [63:0] rdata;
    
    logic [15:0] register_address;
    assign register_address = address[15:0];
    
    logic [63:0]               mtime_n, mtime_q;
    logic [NR_CORES-1:0][63:0] mtimecmp_n, mtimecmp_q;
    logic [NR_CORES-1:0]       msip_n, msip_q;
    
    logic increase_timer;
    
    
    
    axi_lite_interface #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH ),
        .AXI_DATA_WIDTH ( AXI_DATA_WIDTH ),
        .AXI_ID_WIDTH   ( AXI_ID_WIDTH    )
    ) axi_lite_interface_i (
        .clk_i      ( clk_i      ),
        .rst_ni     ( rst_ni     ),
        .axi_req_i  ( axi_req_i  ),
        .axi_resp_o ( axi_resp_o ),
        .address_o  ( address    ),
        .en_o       ( en         ),
        .we_o       ( we         ),
        .data_i     ( rdata      ),
        .data_o     ( wdata      )
    );
    
    
    
    
    always_comb begin
        mtime_n    = mtime_q;
        mtimecmp_n = mtimecmp_q;
        msip_n     = msip_q;
        
        if (increase_timer)
            mtime_n = mtime_q + 1;
        
        if (en && we) begin
            case (register_address) inside
                [MSIP_BASE:MSIP_BASE+4*NR_CORES]: begin
                    msip_n[$unsigned(address[AddrSelWidth-1+2:2])] = wdata[32*address[2]];
                end
                [MTIMECMP_BASE:MTIMECMP_BASE+8*NR_CORES]: begin
                    mtimecmp_n[$unsigned(address[AddrSelWidth-1+3:3])] = wdata;
                end
                MTIME_BASE: begin
                    mtime_n = wdata;
                end
                default:;
            endcase
        end
    end
    
    always_comb begin
        rdata = 'b0;
        if (en && !we) begin
            case (register_address) inside
                [MSIP_BASE:MSIP_BASE+4*NR_CORES]: begin
                    rdata = msip_q[$unsigned(address[AddrSelWidth-1+2:2])];
                end
                [MTIMECMP_BASE:MTIMECMP_BASE+8*NR_CORES]: begin
                    rdata = mtimecmp_q[$unsigned(address[AddrSelWidth-1+3:3])];
                end
                MTIME_BASE: begin
                    rdata = mtime_q;
                end
                default:;
            endcase
        end
    end
    
    
    
    
    
    
    
    
    always_comb begin : irq_gen
        
        for (int unsigned i = 0; i < NR_CORES; i++) begin
            if (mtime_q >= mtimecmp_q[i]) begin
                timer_irq_o[i] = 1'b1;
            end else begin
                timer_irq_o[i] = 1'b0;
            end
        end
    end
    
    
    
    
    
    clint_sync_wedge i_sync_edge (
        .clk_i,
        .rst_ni,
        .serial_i  ( rtc_i          ),
        .r_edge_o  ( increase_timer ),
        .f_edge_o  (                ), 
        .serial_o  (                )  
    );
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (~rst_ni) begin
            mtime_q    <= 64'b0;
            mtimecmp_q <= 'b0;
            msip_q     <= '0;
        end else begin
            mtime_q    <= mtime_n;
            mtimecmp_q <= mtimecmp_n;
            msip_q     <= msip_n;
        end
    end
    assign ipi_o = msip_q;
    
    
    
    
    
    
    
endmodule
module clint_sync_wedge #(
    parameter int unsigned STAGES = 2
) (
    input  logic clk_i,
    input  logic rst_ni,
    input  logic serial_i,
    output logic r_edge_o,
    output logic f_edge_o,
    output logic serial_o
);
    logic serial, serial_q;
    assign serial_o =  serial_q;
    assign f_edge_o = (~serial) & serial_q;
    assign r_edge_o =  serial & (~serial_q);
    clint_sync #(
        .STAGES (STAGES)
    ) i_sync (
        .clk_i,
        .rst_ni,
        .serial_i,
        .serial_o ( serial )
    );
    always_ff @(posedge clk_i, negedge rst_ni) begin
        if (!rst_ni) begin
            serial_q <= 1'b0;
        end else begin
            serial_q <= serial;
        end
    end
endmodule
module clint_sync #(
    parameter int unsigned STAGES = 2
) (
    input  logic clk_i,
    input  logic rst_ni,
    input  logic serial_i,
    output logic serial_o
);
   logic [STAGES-1:0] reg_q;
    always_ff @(posedge clk_i, negedge rst_ni) begin
        if (!rst_ni) begin
            reg_q <= 'h0;
        end else begin
            reg_q <= {reg_q[STAGES-2:0], serial_i};
        end
    end
    assign serial_o = reg_q[STAGES-1];
endmodule
module axi_lite_interface #(
    parameter int unsigned AXI_ADDR_WIDTH = 64,
    parameter int unsigned AXI_DATA_WIDTH = 64,
    parameter int unsigned AXI_ID_WIDTH   = 10
) (
    input logic                       clk_i,    
    input logic                       rst_ni,  
    input  ariane_axi::req_t          axi_req_i,
    output ariane_axi::resp_t         axi_resp_o,
    output logic [AXI_ADDR_WIDTH-1:0] address_o,
    output logic                      en_o,        
    output logic                      we_o,        
    input  logic [AXI_DATA_WIDTH-1:0] data_i,      
    output logic [AXI_DATA_WIDTH-1:0] data_o
);
    
    enum logic [1:0] { IDLE, READ, WRITE, WRITE_B } state_q, state_d;
    
    logic [AXI_ID_WIDTH-1:0]   trans_id_n, trans_id_q;
    
    logic [AXI_ADDR_WIDTH-1:0] address_n,  address_q;
    
    assign axi_resp_o.r.data = data_i;
    
    assign axi_resp_o.r.id = trans_id_q;
    assign axi_resp_o.b.id = trans_id_q;
    
    assign axi_resp_o.r.last = 1'b1;
    
    assign axi_resp_o.b.resp = 2'b0;
    assign axi_resp_o.r.resp = 2'b0;
    
    assign data_o = axi_req_i.w.data;
    
    
    
    always_comb begin
        
        state_d    = state_q;
        address_n  = address_q;
        trans_id_n = trans_id_q;
        
        axi_resp_o.aw_ready = 1'b0;
        axi_resp_o.w_ready  = 1'b0;
        axi_resp_o.b_valid  = 1'b0;
        axi_resp_o.ar_ready = 1'b0;
        axi_resp_o.r_valid  = 1'b0;
        address_o      = '0;
        we_o           = 1'b0;
        en_o           = 1'b0;
        case (state_q)
            
            IDLE: begin
                
                if (axi_req_i.aw_valid) begin
                    axi_resp_o.aw_ready = 1'b1;
                    
                    
                    state_d = WRITE;
                    
                    address_n = axi_req_i.aw.addr;
                    
                    trans_id_n = axi_req_i.aw.id;
                
                end else if (axi_req_i.ar_valid) begin
                    axi_resp_o.ar_ready = 1'b1;
                    state_d = READ;
                    
                    address_n = axi_req_i.ar.addr;
                    
                    trans_id_n = axi_req_i.ar.id;
                end
            end
            
            
            READ: begin
                
                en_o       = 1'b1;
                
                address_o = address_q;
                
                axi_resp_o.r_valid = 1'b1;
                
                if (axi_req_i.r_ready)
                    state_d = IDLE;
            end
            
            
            WRITE: begin
                if (axi_req_i.w_valid) begin
                    axi_resp_o.w_ready = 1'b1;
                    
                    address_o = address_q;
                    en_o = 1'b1;
                    we_o = 1'b1;
                    
                    state_d = WRITE_B;
                end
            end
            WRITE_B: begin
                axi_resp_o.b_valid  = 1'b1;
                
                if (axi_req_i.b_ready)
                    state_d = IDLE;
            end
            default:;
        endcase
    end
    
    
    
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (!rst_ni) begin
            state_q    <= IDLE;
            address_q  <= '0;
            trans_id_q <= '0;
        end else begin
            state_q    <= state_d;
            address_q  <= address_n;
            trans_id_q <= trans_id_n;
        end
    end
    
    
    
    
    
    
    
    
endmodule
module dm_csrs #(
    parameter int                 NrHarts          = 1,
    parameter int                 BusWidth         = 32,
    parameter logic [NrHarts-1:0] SelectableHarts  = 1
) (
    input  logic                              clk_i,           
    input  logic                              rst_ni,          
    input  logic                              testmode_i,
    input  logic                              dmi_rst_ni,      
    input  logic                              dmi_req_valid_i,
    output logic                              dmi_req_ready_o,
    input  dm::dmi_req_t                      dmi_req_i,
    
    output logic                              dmi_resp_valid_o,
    input  logic                              dmi_resp_ready_i,
    output dm::dmi_resp_t                     dmi_resp_o,
    
    output logic                              ndmreset_o,      
    output logic                              dmactive_o,      
                                                               
    
    input  dm::hartinfo_t [NrHarts-1:0]       hartinfo_i,      
    input  logic [NrHarts-1:0]                halted_i,        
    input  logic [NrHarts-1:0]                unavailable_i,   
    input  logic [NrHarts-1:0]                resumeack_i,     
    
    output logic [19:0]                       hartsel_o,       
    output logic [NrHarts-1:0]                haltreq_o,       
    output logic [NrHarts-1:0]                resumereq_o,     
    output logic                              clear_resumeack_o,
    output logic                              cmd_valid_o,       
    output dm::command_t                      cmd_o,             
    input  logic                              cmderror_valid_i,  
    input  dm::cmderr_e                       cmderror_i,        
    input  logic                              cmdbusy_i,         
    output logic [dm::ProgBufSize-1:0][31:0]  progbuf_o, 
    output logic [dm::DataCount-1:0][31:0]    data_o,
    input  logic [dm::DataCount-1:0][31:0]    data_i,
    input  logic                              data_valid_i,
    
    output logic [BusWidth-1:0]               sbaddress_o,
    input  logic [BusWidth-1:0]               sbaddress_i,
    output logic                              sbaddress_write_valid_o,
    
    output logic                              sbreadonaddr_o,
    output logic                              sbautoincrement_o,
    output logic [2:0]                        sbaccess_o,
    
    output logic                              sbreadondata_o,
    output logic [BusWidth-1:0]               sbdata_o,
    output logic                              sbdata_read_valid_o,
    output logic                              sbdata_write_valid_o,
    
    input  logic [BusWidth-1:0]               sbdata_i,
    input  logic                              sbdata_valid_i,
    
    input  logic                              sbbusy_i,
    input  logic                              sberror_valid_i, 
    input  logic [2:0]                        sberror_i 
);
    
    localparam HartSelLen = (NrHarts == 1) ? 1 : $clog2(NrHarts);
    dm::dtm_op_e dtm_op;
    assign dtm_op = dm::dtm_op_e'(dmi_req_i.op);
    logic        resp_queue_full;
    logic        resp_queue_empty;
    logic        resp_queue_push;
    logic        resp_queue_pop;
    logic [31:0] resp_queue_data;
    localparam dm::dm_csr_e DataEnd = dm::dm_csr_e'((dm::Data0 + {4'b0, dm::DataCount}));
    localparam dm::dm_csr_e ProgBufEnd = dm::dm_csr_e'((dm::ProgBuf0 + {4'b0, dm::ProgBufSize}));
    logic [31:0] haltsum0, haltsum1, haltsum2, haltsum3;
    logic [NrHarts/2**5 :0][31:0] halted_reshaped0;
    logic [NrHarts/2**10:0][31:0] halted_reshaped1;
    logic [NrHarts/2**15:0][31:0] halted_reshaped2;
    logic [(NrHarts/2**10+1)*32-1:0] halted_flat1;
    logic [(NrHarts/2**15+1)*32-1:0] halted_flat2;
    logic [32-1:0] halted_flat3;
    
    assign halted_reshaped0 = halted_i;
    assign haltsum0         = halted_reshaped0[hartsel_o[19:5]];
    
    always_comb begin : p_reduction1
        halted_flat1 = '0;
        for (int k=0; k<NrHarts/2**5+1; k++) begin
            halted_flat1[k] = |halted_reshaped0[k];
        end
        halted_reshaped1 = halted_flat1;
        haltsum1         = halted_reshaped1[hartsel_o[19:10]];
    end
    
    always_comb begin : p_reduction2
        halted_flat2 = '0;
        for (int k=0; k<NrHarts/2**10+1; k++) begin
            halted_flat2[k] = |halted_reshaped1[k];
        end
        halted_reshaped2 = halted_flat2;
        haltsum2         = halted_reshaped2[hartsel_o[19:15]];
    end
    
    always_comb begin : p_reduction3
        halted_flat3 = '0;
        for (int k=0; k<NrHarts/2**15+1; k++) begin
            halted_flat3[k] = |halted_reshaped2[k];
        end
        haltsum3 = halted_flat3;
    end
    dm::dmstatus_t      dmstatus;
    dm::dmcontrol_t     dmcontrol_d, dmcontrol_q;
    dm::abstractcs_t    abstractcs;
    dm::cmderr_e        cmderr_d, cmderr_q;
    dm::command_t       command_d, command_q;
    logic               cmd_valid_d, cmd_valid_q;
    dm::abstractauto_t  abstractauto_d, abstractauto_q;
    dm::sbcs_t          sbcs_d, sbcs_q;
    logic [63:0]        sbaddr_d, sbaddr_q;
    logic [63:0]        sbdata_d, sbdata_q;
    logic [NrHarts-1:0] havereset_d, havereset_q;
    
    logic [dm::ProgBufSize-1:0][31:0] progbuf_d, progbuf_q;
    
    logic [({3'b0, dm::DataCount} + dm::Data0 - 1):(dm::Data0)][31:0] data_d, data_q;
    logic [HartSelLen-1:0] selected_hart;
    
    assign dmi_resp_o.resp = dm::DTM_SUCCESS;
    assign dmi_resp_valid_o     = ~resp_queue_empty;
    assign dmi_req_ready_o      = ~resp_queue_full;
    assign resp_queue_push      = dmi_req_valid_i & dmi_req_ready_o;
    
    assign sbautoincrement_o = sbcs_q.sbautoincrement;
    assign sbreadonaddr_o    = sbcs_q.sbreadonaddr;
    assign sbreadondata_o    = sbcs_q.sbreadondata;
    assign sbaccess_o        = sbcs_q.sbaccess;
    assign sbdata_o          = sbdata_q[BusWidth-1:0];
    assign sbaddress_o       = sbaddr_q[BusWidth-1:0];
    assign hartsel_o         = {dmcontrol_q.hartselhi, dmcontrol_q.hartsello};
    always_comb begin : csr_read_write
        
        
        
        
        dmstatus    = '0;
        dmstatus.version = dm::DbgVersion013;
        
        dmstatus.authenticated = 1'b1;
        
        dmstatus.hasresethaltreq = 1'b0;
        
        dmstatus.allhavereset = havereset_q[selected_hart];
        dmstatus.anyhavereset = havereset_q[selected_hart];
        dmstatus.allresumeack = resumeack_i[selected_hart];
        dmstatus.anyresumeack = resumeack_i[selected_hart];
        dmstatus.allunavail   = unavailable_i[selected_hart];
        dmstatus.anyunavail   = unavailable_i[selected_hart];
        
        
        dmstatus.allnonexistent = (hartsel_o > (NrHarts[19:0] - 1)) ? 1'b1 : 1'b0;
        dmstatus.anynonexistent = (hartsel_o > (NrHarts[19:0] - 1)) ? 1'b1 : 1'b0;
        
        
        dmstatus.allhalted    = halted_i[selected_hart] & ~unavailable_i[selected_hart];
        dmstatus.anyhalted    = halted_i[selected_hart] & ~unavailable_i[selected_hart];
        dmstatus.allrunning   = ~halted_i[selected_hart] & ~unavailable_i[selected_hart];
        dmstatus.anyrunning   = ~halted_i[selected_hart] & ~unavailable_i[selected_hart];
        
        abstractcs = '0;
        abstractcs.datacount = dm::DataCount;
        abstractcs.progbufsize = dm::ProgBufSize;
        abstractcs.busy = cmdbusy_i;
        abstractcs.cmderr = cmderr_q;
        
        abstractauto_d = abstractauto_q;
        abstractauto_d.zero0 = '0;
        
        havereset_d = havereset_q;
        dmcontrol_d = dmcontrol_q;
        cmderr_d    = cmderr_q;
        command_d   = command_q;
        progbuf_d   = progbuf_q;
        data_d      = data_q;
        sbcs_d      = sbcs_q;
        sbaddr_d    = sbaddress_i;
        sbdata_d    = sbdata_q;
        resp_queue_data         = 32'b0;
        cmd_valid_d             = 1'b0;
        sbaddress_write_valid_o = 1'b0;
        sbdata_read_valid_o     = 1'b0;
        sbdata_write_valid_o    = 1'b0;
        clear_resumeack_o       = 1'b0;
        
        if (dmi_req_ready_o && dmi_req_valid_i && dtm_op == dm::DTM_READ) begin
            unique case ({1'b0, dmi_req_i.addr}) inside
                [(dm::Data0):DataEnd]: begin
                    if (dm::DataCount > 0) begin
                        resp_queue_data = data_q[dmi_req_i.addr[4:0]];
                    end
                    if (!cmdbusy_i) begin
                        
                        cmd_valid_d = abstractauto_q.autoexecdata[dmi_req_i.addr[3:0] -
                                      int'(dm::Data0)];
                    end
                end
                dm::DMControl:    resp_queue_data = dmcontrol_q;
                dm::DMStatus:     resp_queue_data = dmstatus;
                dm::Hartinfo:     resp_queue_data = hartinfo_i[selected_hart];
                dm::AbstractCS:   resp_queue_data = abstractcs;
                dm::AbstractAuto: resp_queue_data = abstractauto_q;
                
                dm::Command:    resp_queue_data = '0;
                [(dm::ProgBuf0):ProgBufEnd]: begin
                    resp_queue_data = progbuf_q[dmi_req_i.addr[4:0]];
                    if (!cmdbusy_i) begin
                        
                        
                        cmd_valid_d = abstractauto_q.autoexecprogbuf[dmi_req_i.addr[3:0]+16];
                    end
                end
                dm::HaltSum0: resp_queue_data = haltsum0;
                dm::HaltSum1: resp_queue_data = haltsum1;
                dm::HaltSum2: resp_queue_data = haltsum2;
                dm::HaltSum3: resp_queue_data = haltsum3;
                dm::SBCS: begin
                    resp_queue_data = sbcs_q;
                end
                dm::SBAddress0: begin
                    
                    if (sbbusy_i) begin
                       sbcs_d.sbbusyerror = 1'b1;
                    end else begin
                        resp_queue_data = sbaddr_q[31:0];
                    end
                end
                dm::SBAddress1: begin
                    
                    if (sbbusy_i) begin
                       sbcs_d.sbbusyerror = 1'b1;
                    end else begin
                        resp_queue_data = sbaddr_q[63:32];
                    end
                end
                dm::SBData0: begin
                    
                    if (sbbusy_i) begin
                       sbcs_d.sbbusyerror = 1'b1;
                    end else begin
                        sbdata_read_valid_o = (sbcs_q.sberror == '0);
                        resp_queue_data = sbdata_q[31:0];
                    end
                end
                dm::SBData1: begin
                    
                    if (sbbusy_i) begin
                       sbcs_d.sbbusyerror = 1'b1;
                    end else begin
                        resp_queue_data = sbdata_q[63:32];
                    end
                end
                default:;
            endcase
        end
        
        if (dmi_req_ready_o && dmi_req_valid_i && dtm_op == dm::DTM_WRITE) begin
            unique case (dm::dm_csr_e'({1'b0, dmi_req_i.addr})) inside
                [(dm::Data0):DataEnd]: begin
                    
                    if (!cmdbusy_i && dm::DataCount > 0) begin
                        data_d[dmi_req_i.addr[4:0]] = dmi_req_i.data;
                        
                        cmd_valid_d = abstractauto_q.autoexecdata[dmi_req_i.addr[3:0] -
                                      int'(dm::Data0)];
                    end
                end
                dm::DMControl: begin
                    automatic dm::dmcontrol_t dmcontrol;
                    dmcontrol = dm::dmcontrol_t'(dmi_req_i.data);
                    
                    if (dmcontrol.ackhavereset) begin
                        havereset_d[selected_hart] = 1'b0;
                    end
                    dmcontrol_d = dmi_req_i.data;
                end
                dm::DMStatus:; 
                dm::Hartinfo:; 
                
                dm::AbstractCS: begin 
                    
                    
                    
                    
                    automatic dm::abstractcs_t a_abstractcs;
                    a_abstractcs = dm::abstractcs_t'(dmi_req_i.data);
                    
                    if (!cmdbusy_i) begin
                        cmderr_d = dm::cmderr_e'(~a_abstractcs.cmderr & cmderr_q);
                    end else if (cmderr_q == dm::CmdErrNone) begin
                        cmderr_d = dm::CmdErrBusy;
                    end
                end
                dm::Command: begin
                    
                    if (!cmdbusy_i) begin
                        cmd_valid_d = 1'b1;
                        command_d = dm::command_t'(dmi_req_i.data);
                    
                    
                    end else if (cmderr_q == dm::CmdErrNone) begin
                        cmderr_d = dm::CmdErrBusy;
                    end
                end
                dm::AbstractAuto: begin
                    
                    if (!cmdbusy_i) begin
                        abstractauto_d                 = 32'b0;
                        abstractauto_d.autoexecdata    = dmi_req_i.data[dm::DataCount-1:0];
                        abstractauto_d.autoexecprogbuf = dmi_req_i.data[dm::ProgBufSize-1+16:16];
                    end else if (cmderr_q == dm::CmdErrNone) begin
                        cmderr_d = dm::CmdErrBusy;
                    end
                end
                [(dm::ProgBuf0):ProgBufEnd]: begin
                    
                    if (!cmdbusy_i) begin
                        progbuf_d[dmi_req_i.addr[4:0]] = dmi_req_i.data;
                        
                        
                        
                        
                        
                        cmd_valid_d = abstractauto_q.autoexecprogbuf[dmi_req_i.addr[3:0]+16];
                    end
                end
                dm::SBCS: begin
                    
                    if (sbbusy_i) begin
                        sbcs_d.sbbusyerror = 1'b1;
                    end else begin
                        automatic dm::sbcs_t sbcs = dm::sbcs_t'(dmi_req_i.data);
                        sbcs_d = sbcs;
                        
                        sbcs_d.sbbusyerror = sbcs_q.sbbusyerror & (~sbcs.sbbusyerror);
                        sbcs_d.sberror     = sbcs_q.sberror     & (~sbcs.sberror);
                    end
                end
                dm::SBAddress0: begin
                    
                    if (sbbusy_i) begin
                       sbcs_d.sbbusyerror = 1'b1;
                    end else begin
                        sbaddr_d[31:0] = dmi_req_i.data;
                        sbaddress_write_valid_o = (sbcs_q.sberror == '0);
                    end
                end
                dm::SBAddress1: begin
                    
                    if (sbbusy_i) begin
                       sbcs_d.sbbusyerror = 1'b1;
                    end else begin
                        sbaddr_d[63:32] = dmi_req_i.data;
                    end
                end
                dm::SBData0: begin
                    
                    if (sbbusy_i) begin
                       sbcs_d.sbbusyerror = 1'b1;
                    end else begin
                        sbdata_d[31:0] = dmi_req_i.data;
                        sbdata_write_valid_o = (sbcs_q.sberror == '0);
                    end
                end
                dm::SBData1: begin
                    
                    if (sbbusy_i) begin
                       sbcs_d.sbbusyerror = 1'b1;
                    end else begin
                        sbdata_d[63:32] = dmi_req_i.data;
                    end
                end
                default:;
            endcase
        end
        
        if (cmderror_valid_i) begin
            cmderr_d = cmderror_i;
        end
        
        if (data_valid_i)
            data_d = data_i;
        
        if (ndmreset_o) begin
            havereset_d = '1;
        end
        
        
        
        
        if (sberror_valid_i) begin
            sbcs_d.sberror = sberror_i;
        end
        
        if (sbdata_valid_i) begin
            sbdata_d = sbdata_i;
        end
        
        
        dmcontrol_d.hasel           = 1'b0;
        
        dmcontrol_d.hartreset       = 1'b0;
        dmcontrol_d.setresethaltreq = 1'b0;
        dmcontrol_d.clrresethaltreq = 1'b0;
        dmcontrol_d.zero1           = '0;
        dmcontrol_d.zero0           = '0;
        
        dmcontrol_d.ackhavereset    = 1'b0;
        if (!dmcontrol_q.resumereq && dmcontrol_d.resumereq) begin
            clear_resumeack_o = 1'b1;
        end
        if (dmcontrol_q.resumereq && resumeack_i) begin
            dmcontrol_d.resumereq = 1'b0;
        end
        
        sbcs_d.sbversion            = 3'b1;
        sbcs_d.sbbusy               = sbbusy_i;
        sbcs_d.sbasize              = BusWidth;
        sbcs_d.sbaccess128          = 1'b0;
        sbcs_d.sbaccess64           = BusWidth == 64;
        sbcs_d.sbaccess32           = BusWidth == 32;
        sbcs_d.sbaccess16           = 1'b0;
        sbcs_d.sbaccess8            = 1'b0;
        sbcs_d.sbaccess             = BusWidth == 64 ? 2'd3 : 2'd2;
    end
    
    always_comb begin
        selected_hart = hartsel_o[HartSelLen-1:0];
        
        haltreq_o = '0;
        resumereq_o = '0;
        haltreq_o[selected_hart] = dmcontrol_q.haltreq;
        resumereq_o[selected_hart] = dmcontrol_q.resumereq;
    end
    assign dmactive_o  = dmcontrol_q.dmactive;
    assign cmd_o       = command_q;
    assign cmd_valid_o = cmd_valid_q;
    assign progbuf_o   = progbuf_q;
    assign data_o      = data_q;
    assign resp_queue_pop = dmi_resp_ready_i & ~resp_queue_empty;
    assign ndmreset_o = dmcontrol_q.ndmreset;
    
    fifo_v2 #(
        .dtype            ( logic [31:0]         ),
        .DEPTH            ( 2                    )
    ) i_fifo (
        .clk_i            ( clk_i                ),
        .rst_ni           ( dmi_rst_ni           ), 
        .flush_i          ( 1'b0                 ), 
        .testmode_i       ( testmode_i           ),
        .full_o           ( resp_queue_full      ),
        .empty_o          ( resp_queue_empty     ),
        .alm_full_o       (                      ),
        .alm_empty_o      (                      ),
        .data_i           ( resp_queue_data      ),
        .push_i           ( resp_queue_push      ),
        .data_o           ( dmi_resp_o.data      ),
        .pop_i            ( resp_queue_pop       )
    );
    always_ff @(posedge clk_i or negedge rst_ni) begin
        
        if (!rst_ni) begin
            dmcontrol_q    <= '0;
            
            cmderr_q       <= dm::CmdErrNone;
            command_q      <= '0;
            abstractauto_q <= '0;
            progbuf_q      <= '0;
            data_q         <= '0;
            sbcs_q         <= '0;
            sbaddr_q       <= '0;
            sbdata_q       <= '0;
        end else begin
            
            if (!dmcontrol_q.dmactive) begin
                dmcontrol_q.haltreq          <= '0;
                dmcontrol_q.resumereq        <= '0;
                dmcontrol_q.hartreset        <= '0;
                dmcontrol_q.zero1            <= '0;
                dmcontrol_q.hasel            <= '0;
                dmcontrol_q.hartsello        <= '0;
                dmcontrol_q.hartselhi        <= '0;
                dmcontrol_q.zero0            <= '0;
                dmcontrol_q.setresethaltreq  <= '0;
                dmcontrol_q.clrresethaltreq  <= '0;
                dmcontrol_q.ndmreset         <= '0;
                
                dmcontrol_q.dmactive         <= dmcontrol_d.dmactive;
                cmderr_q                     <= dm::CmdErrNone;
                command_q                    <= '0;
                cmd_valid_q                  <= '0;
                abstractauto_q               <= '0;
                progbuf_q                    <= '0;
                data_q                       <= '0;
                sbcs_q                       <= '0;
                sbaddr_q                     <= '0;
                sbdata_q                     <= '0;
            end else begin
                dmcontrol_q                  <= dmcontrol_d;
                cmderr_q                     <= cmderr_d;
                command_q                    <= command_d;
                cmd_valid_q                  <= cmd_valid_d;
                abstractauto_q               <= abstractauto_d;
                progbuf_q                    <= progbuf_d;
                data_q                       <= data_d;
                sbcs_q                       <= sbcs_d;
                sbaddr_q                     <= sbaddr_d;
                sbdata_q                     <= sbdata_d;
            end
        end
    end
    for (genvar k = 0; k < NrHarts; k++) begin : gen_havereset
        always_ff @(posedge clk_i or negedge rst_ni) begin
            if (!rst_ni) begin
                havereset_q[k] <= 1'b1;
            end else begin
                havereset_q[k] <= SelectableHarts[k] ? havereset_d[k] : 1'b0;
            end
        end
    end
endmodule
module dm_mem #(
    parameter int                 NrHarts          = -1,
    parameter int                 BusWidth         = -1,
    parameter logic [NrHarts-1:0] SelectableHarts  = -1
)(
    input  logic                             clk_i,       
    input  logic                             rst_ni,      
    output logic [NrHarts-1:0]               debug_req_o,
    input  logic [19:0]                      hartsel_i,
    
    input  logic [NrHarts-1:0]               haltreq_i,
    input  logic [NrHarts-1:0]               resumereq_i,
    input  logic                             clear_resumeack_i,
    
    output logic [NrHarts-1:0]               halted_o,    
    output logic [NrHarts-1:0]               resuming_o,  
    input  logic [dm::ProgBufSize-1:0][31:0] progbuf_i,    
    input  logic [dm::DataCount-1:0][31:0]   data_i,       
    output logic [dm::DataCount-1:0][31:0]   data_o,       
    output logic                             data_valid_o, 
    
    input  logic                             cmd_valid_i,
    input  dm::command_t                     cmd_i,
    output logic                             cmderror_valid_o,
    output dm::cmderr_e                      cmderror_o,
    output logic                             cmdbusy_o,
    
    
    input  logic                             req_i,
    input  logic                             we_i,
    input  logic [BusWidth-1:0]              addr_i,
    input  logic [BusWidth-1:0]              wdata_i,
    input  logic [BusWidth/8-1:0]            be_i,
    output logic [BusWidth-1:0]              rdata_o
);
    localparam int HartSelLen = (NrHarts == 1) ? 1 : $clog2(NrHarts);
    localparam int MaxAar = (BusWidth == 64) ? 4 : 3;
    localparam DbgAddressBits = 12;
    localparam logic [DbgAddressBits-1:0] DataBase = (dm::DataAddr);
    localparam logic [DbgAddressBits-1:0] DataEnd = (dm::DataAddr + 4*dm::DataCount);
    localparam logic [DbgAddressBits-1:0] ProgBufBase = (dm::DataAddr - 4*dm::ProgBufSize);
    localparam logic [DbgAddressBits-1:0] ProgBufEnd = (dm::DataAddr - 1);
    localparam logic [DbgAddressBits-1:0] AbstractCmdBase = (ProgBufBase - 4*10);
    localparam logic [DbgAddressBits-1:0] AbstractCmdEnd = (ProgBufBase - 1);
    localparam logic [DbgAddressBits-1:0] WhereTo   = 'h300;
    localparam logic [DbgAddressBits-1:0] FlagsBase = 'h400;
    localparam logic [DbgAddressBits-1:0] FlagsEnd  = 'h7FF;
    localparam logic [DbgAddressBits-1:0] Halted    = 'h100;
    localparam logic [DbgAddressBits-1:0] Going     = 'h104;
    localparam logic [DbgAddressBits-1:0] Resuming  = 'h108;
    localparam logic [DbgAddressBits-1:0] Exception = 'h10C;
    logic [dm::ProgBufSize/2-1:0][63:0]   progbuf;
    logic [4:0][63:0]   abstract_cmd;
    logic [NrHarts-1:0] halted_d, halted_q;
    logic [NrHarts-1:0] resuming_d, resuming_q;
    logic               resume, go, going;
    logic [NrHarts-1:0] halted;
    logic [HartSelLen-1:0] hart_sel;
    logic exception;
    logic unsupported_command;
    logic [63:0] rom_rdata;
    logic [63:0] rdata_d, rdata_q;
    logic        word_enable32_q;
    
    
    logic fwd_rom_d, fwd_rom_q;
    dm::ac_ar_cmd_t ac_ar;
    
    assign ac_ar       = dm::ac_ar_cmd_t'(cmd_i.control);
    assign hart_sel    = wdata_i[HartSelLen-1:0];
    assign debug_req_o = haltreq_i;
    assign halted_o    = halted_q;
    assign resuming_o  = resuming_q;
    
    assign progbuf = progbuf_i;
    typedef enum logic [1:0] { Idle, Go, Resume, CmdExecuting } state_e;
    state_e state_d, state_q;
    
    always_comb begin
        cmderror_valid_o = 1'b0;
        cmderror_o       = dm::CmdErrNone;
        state_d          = state_q;
        go               = 1'b0;
        resume           = 1'b0;
        cmdbusy_o        = 1'b1;
        case (state_q)
            Idle: begin
                cmdbusy_o = 1'b0;
                if (cmd_valid_i && halted_q[hartsel_i]) begin
                    
                    state_d = Go;
                end else if (cmd_valid_i) begin
                    
                    cmderror_valid_o = 1'b1;
                    cmderror_o = dm::CmdErrorHaltResume;
                end
                
                
                if (resumereq_i[hartsel_i] && !resuming_q[hartsel_i] &&
                     !haltreq_i[hartsel_i] &&    halted_q[hartsel_i]) begin
                    state_d = Resume;
                end
            end
            Go: begin
                
                cmdbusy_o = 1'b1;
                go        = 1'b1;
                
                if (going)
                    state_d = CmdExecuting;
            end
            Resume: begin
                cmdbusy_o = 1'b1;
                resume = 1'b1;
                if (resuming_o[hartsel_i])
                    state_d = Idle;
            end
            CmdExecuting: begin
                cmdbusy_o = 1'b1;
                go        = 1'b0;
                
                if (halted[hartsel_i]) begin
                    state_d = Idle;
                end
            end
        endcase
        
        
        if (unsupported_command && cmd_valid_i) begin
            cmderror_valid_o = 1'b1;
            cmderror_o = dm::CmdErrNotSupported;
        end
        if (exception) begin
            cmderror_valid_o = 1'b1;
            cmderror_o = dm::CmdErrorException;
        end
    end
    
    always_comb begin
        automatic logic [63:0] data_bits;
        halted_d     = halted_q;
        resuming_d   = resuming_q;
        rdata_o      = (BusWidth == 64) ?
                          (fwd_rom_q ? rom_rdata : rdata_q) :
                          (word_enable32_q ?
                              (fwd_rom_q ? rom_rdata[63:32] : rdata_q[63:32]) :
                              (fwd_rom_q ? rom_rdata[31: 0] : rdata_q[31: 0]));
        rdata_d      = rdata_q;
        
        data_bits    = data_i;
        
        data_valid_o = 1'b0;
        exception    = 1'b0;
        halted       = '0;
        going        = 1'b0;
        
        if (clear_resumeack_i) begin
            resuming_d[hartsel_i] = 1'b0;
        end
        
        if (req_i) begin
            
            if (we_i) begin
                unique case (addr_i[DbgAddressBits-1:0]) inside
                    Halted: begin
                        halted[hart_sel] = 1'b1;
                        halted_d[hart_sel] = 1'b1;
                    end
                    Going: begin
                        going = 1'b1;
                    end
                    Resuming: begin
                        
                        halted_d[hart_sel] = 1'b0;
                        
                        resuming_d[hart_sel] = 1'b1;
                    end
                    
                    Exception: exception = 1'b1;
                    
                    [(dm::DataAddr):DataEnd]: begin
                        data_valid_o = 1'b1;
                        for (int i = 0; i < $bits(be_i); i++) begin
                            if (be_i[i]) begin
                                data_bits[i*8+:8] = wdata_i[i*8+:8];
                            end
                        end
                    end
                    default ;
                endcase
            
            end else begin
                unique case (addr_i[DbgAddressBits-1:0]) inside
                    
                    WhereTo: begin
                        
                        if (resumereq_i[hart_sel]) begin
                            rdata_d = {32'b0, dm::jal('0, dm::ResumeAddress[11:0]-WhereTo)};
                        end
                        
                        if (cmdbusy_o) begin
                            
                            
                            if (cmd_i.cmdtype == dm::AccessRegister &&
                                !ac_ar.transfer && ac_ar.postexec) begin
                                rdata_d = {32'b0, dm::jal('0, ProgBufBase-WhereTo)};
                            
                            end else begin
                                rdata_d = {32'b0, dm::jal('0, AbstractCmdBase-WhereTo)};
                            end
                        end
                    end
                    [DataBase:DataEnd]: begin
                        rdata_d = {
                                  data_i[(addr_i[DbgAddressBits-1:3] - DataBase[DbgAddressBits-1:3] + 1)],
                                  data_i[(addr_i[DbgAddressBits-1:3] - DataBase[DbgAddressBits-1:3])]
                                  };
                    end
                    [ProgBufBase:ProgBufEnd]: begin
                        rdata_d = progbuf[(addr_i[DbgAddressBits-1:3] -
                                      ProgBufBase[DbgAddressBits-1:3])];
                    end
                    
                    [AbstractCmdBase:AbstractCmdEnd]: begin
                        
                        rdata_d = abstract_cmd[(addr_i[DbgAddressBits-1:3] -
                                       AbstractCmdBase[DbgAddressBits-1:3])];
                    end
                    
                    [FlagsBase:FlagsEnd]: begin
                        automatic logic [7:0][7:0] rdata;
                        rdata = '0;
                        
                        if (({addr_i[DbgAddressBits-1:3], 3'b0} - FlagsBase[DbgAddressBits-1:0]) ==
                          {hartsel_i[DbgAddressBits-1:3], 3'b0}) begin
                            rdata[hartsel_i[2:0]] = {6'b0, resume, go};
                        end
                        rdata_d = rdata;
                    end
                    default: ;
                endcase
            end
        end
        data_o = data_bits;
    end
    always_comb begin : abstract_cmd_rom
        
        unsupported_command = 1'b0;
        
        
        abstract_cmd[0][31:0]  = dm::illegal();
        
        abstract_cmd[0][63:32] = dm::auipc(5'd10, '0);
        abstract_cmd[1][31:0]  = dm::srli(5'd10, 5'd10, 6'd12); 
        abstract_cmd[1][63:32] = dm::slli(5'd10, 5'd10, 6'd12);
        abstract_cmd[2][31:0]  = dm::nop();
        abstract_cmd[2][63:32] = dm::nop();
        abstract_cmd[3][31:0]  = dm::nop();
        abstract_cmd[3][63:32] = dm::nop();
        abstract_cmd[4][31:0]  = dm::csrr(dm::CSR_DSCRATCH1, 5'd10);
        abstract_cmd[4][63:32] = dm::ebreak();
        
        unique case (cmd_i.cmdtype)
            
            
            
            dm::AccessRegister: begin
                if (ac_ar.aarsize < MaxAar && ac_ar.transfer && ac_ar.write) begin
                    
                    abstract_cmd[0][31:0] = dm::csrw(dm::CSR_DSCRATCH1, 5'd10);
                    
                    if (ac_ar.regno[15:14] != '0) begin
                        abstract_cmd[0][31:0] = dm::ebreak(); 
                        unsupported_command = 1'b1;
                    
                    
                    end else if (ac_ar.regno[12] && (!ac_ar.regno[5]) &&
                                (ac_ar.regno[4:0] == 5'd10)) begin
                        
                        abstract_cmd[2][31:0]  = dm::csrw(dm::CSR_DSCRATCH0, 5'd8);
                        
                        abstract_cmd[2][63:32] = dm::load(ac_ar.aarsize, 5'd8, 5'd10, dm::DataAddr);
                        
                        abstract_cmd[3][31:0]  = dm::csrw(dm::CSR_DSCRATCH1, 5'd8);
                        
                        abstract_cmd[3][63:32] = dm::csrr(dm::CSR_DSCRATCH0, 5'd8);
                    
                    end else if (ac_ar.regno[12]) begin
                        
                        if (ac_ar.regno[5]) begin
                            abstract_cmd[2][31:0] =
                                dm::float_load(ac_ar.aarsize, ac_ar.regno[4:0], 5'd10, dm::DataAddr);
                        end else begin
                            abstract_cmd[2][31:0] =
                                dm::load(ac_ar.aarsize, ac_ar.regno[4:0], 5'd10, dm::DataAddr);
                        end
                    
                    end else begin
                        
                        
                        abstract_cmd[2][31:0]  = dm::csrw(dm::CSR_DSCRATCH0, 5'd8);
                        
                        abstract_cmd[2][63:32] = dm::load(ac_ar.aarsize, 5'd8, 5'd10, dm::DataAddr);
                        
                        abstract_cmd[3][31:0]  = dm::csrw(dm::csr_reg_t'(ac_ar.regno[11:0]), 5'd8);
                        
                        abstract_cmd[3][63:32] = dm::csrr(dm::CSR_DSCRATCH0, 5'd8);
                    end
                end else if (ac_ar.aarsize < MaxAar && ac_ar.transfer && !ac_ar.write) begin
                    
                    abstract_cmd[0][31:0]  = dm::csrw(dm::CSR_DSCRATCH1, 5'd10);
                    
                    if (ac_ar.regno[15:14] != '0) begin
                        abstract_cmd[0][31:0] = dm::ebreak(); 
                        unsupported_command = 1'b1;
                    
                    
                    end else if (ac_ar.regno[12] && (!ac_ar.regno[5]) &&
                                (ac_ar.regno[4:0] == 5'd10)) begin
                        
                        abstract_cmd[2][31:0]  = dm::csrw(dm::CSR_DSCRATCH0, 5'd8);
                        
                        abstract_cmd[2][63:32] = dm::csrr(dm::CSR_DSCRATCH1, 5'd8);
                        
                        abstract_cmd[3][31:0]  = dm::store(ac_ar.aarsize, 5'd8, 5'd10, dm::DataAddr);
                        
                        abstract_cmd[3][63:32] = dm::csrr(dm::CSR_DSCRATCH0, 5'd8);
                    
                    end else if (ac_ar.regno[12]) begin
                        
                        if (ac_ar.regno[5]) begin
                            abstract_cmd[2][31:0] =
                                dm::float_store(ac_ar.aarsize, ac_ar.regno[4:0], 5'd10, dm::DataAddr);
                        end else begin
                            abstract_cmd[2][31:0] =
                                dm::store(ac_ar.aarsize, ac_ar.regno[4:0], 5'd10, dm::DataAddr);
                        end
                    
                    end else begin
                        
                        
                        abstract_cmd[2][31:0]  = dm::csrw(dm::CSR_DSCRATCH0, 5'd8);
                        
                        abstract_cmd[2][63:32] = dm::csrr(dm::csr_reg_t'(ac_ar.regno[11:0]), 5'd8);
                        
                        abstract_cmd[3][31:0]  = dm::store(ac_ar.aarsize, 5'd8, 5'd10, dm::DataAddr);
                        
                        abstract_cmd[3][63:32] = dm::csrr(dm::CSR_DSCRATCH0, 5'd8);
                    end
                end else if (ac_ar.aarsize >= MaxAar || ac_ar.aarpostincrement == 1'b1) begin
                    
                    
                    
                    abstract_cmd[0][31:0] = dm::ebreak(); 
                    unsupported_command = 1'b1;
                end
                
                
                
                
                if (ac_ar.postexec && !unsupported_command) begin
                    
                    abstract_cmd[4][63:32] = dm::nop();
                end
            end
            
            
            
            default: begin
                abstract_cmd[0][31:0] = dm::ebreak();
                unsupported_command = 1'b1;
            end
        endcase
    end
    logic [63:0] rom_addr;
    assign rom_addr = addr_i;
    debug_rom i_debug_rom (
        .clk_i,
        .req_i,
        .addr_i  ( rom_addr  ),
        .rdata_o ( rom_rdata )
    );
    
    
    assign fwd_rom_d = (addr_i[DbgAddressBits-1:0] >= dm::HaltAddress[DbgAddressBits-1:0]) ?
                           1'b1 : 1'b0;
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (!rst_ni) begin
            fwd_rom_q       <= 1'b0;
            rdata_q         <= '0;
            state_q         <= Idle;
            word_enable32_q <= 1'b0;
        end else begin
            fwd_rom_q       <= fwd_rom_d;
            rdata_q         <= rdata_d;
            state_q         <= state_d;
            word_enable32_q <= addr_i[2];
        end
    end
    for (genvar k = 0; k < NrHarts; k++) begin : gen_halted
        always_ff @(posedge clk_i or negedge rst_ni) begin
            if (!rst_ni) begin
                halted_q[k]   <= 1'b0;
                resuming_q[k] <= 1'b0;
            end else begin
                halted_q[k]   <= SelectableHarts[k] ? halted_d[k]   : 1'b0;
                resuming_q[k] <= SelectableHarts[k] ? resuming_d[k] : 1'b0;
            end
        end
    end
endmodule
module dm_top #(
    parameter int                 NrHarts          = 1,
    parameter int                 BusWidth         = 32,
    parameter logic [NrHarts-1:0] SelectableHarts  = 1  
                                                        
) (
    input  logic                  clk_i,       
    input  logic                  rst_ni,      
    input  logic                  testmode_i,
    output logic                  ndmreset_o,  
    output logic                  dmactive_o,  
    output logic [NrHarts-1:0]    debug_req_o, 
    input  logic [NrHarts-1:0]    unavailable_i, 
    dm::hartinfo_t [NrHarts-1:0]  hartinfo_i,
    input  logic                  slave_req_i,
    input  logic                  slave_we_i,
    input  logic [BusWidth-1:0]   slave_addr_i,
    input  logic [BusWidth/8-1:0] slave_be_i,
    input  logic [BusWidth-1:0]   slave_wdata_i,
    output logic [BusWidth-1:0]   slave_rdata_o,
    output logic                  master_req_o,
    output logic [BusWidth-1:0]   master_add_o,
    output logic                  master_we_o,
    output logic [BusWidth-1:0]   master_wdata_o,
    output logic [BusWidth/8-1:0] master_be_o,
    input  logic                  master_gnt_i,
    input  logic                  master_r_valid_i,
    input  logic [BusWidth-1:0]   master_r_rdata_i,
    
    input  logic                  dmi_rst_ni,
    input  logic                  dmi_req_valid_i,
    output logic                  dmi_req_ready_o,
    input  dm::dmi_req_t          dmi_req_i,
    output logic                  dmi_resp_valid_o,
    input  logic                  dmi_resp_ready_i,
    output dm::dmi_resp_t         dmi_resp_o
);
    
    logic [NrHarts-1:0]               halted;
    
    logic [NrHarts-1:0]               resumeack;
    logic [NrHarts-1:0]               haltreq;
    logic [NrHarts-1:0]               resumereq;
    logic                             clear_resumeack;
    logic                             cmd_valid;
    dm::command_t                     cmd;
    logic                             cmderror_valid;
    dm::cmderr_e                      cmderror;
    logic                             cmdbusy;
    logic [dm::ProgBufSize-1:0][31:0] progbuf;
    logic [dm::DataCount-1:0][31:0]   data_csrs_mem;
    logic [dm::DataCount-1:0][31:0]   data_mem_csrs;
    logic                             data_valid;
    logic [19:0]                      hartsel;
    
    logic [BusWidth-1:0]              sbaddress_csrs_sba;
    logic [BusWidth-1:0]              sbaddress_sba_csrs;
    logic                             sbaddress_write_valid;
    logic                             sbreadonaddr;
    logic                             sbautoincrement;
    logic [2:0]                       sbaccess;
    logic                             sbreadondata;
    logic [BusWidth-1:0]              sbdata_write;
    logic                             sbdata_read_valid;
    logic                             sbdata_write_valid;
    logic [BusWidth-1:0]              sbdata_read;
    logic                             sbdata_valid;
    logic                             sbbusy;
    logic                             sberror_valid;
    logic [2:0]                       sberror;
    dm_csrs #(
        .NrHarts(NrHarts),
        .BusWidth(BusWidth),
        .SelectableHarts(SelectableHarts)
    ) i_dm_csrs (
        .clk_i                   ( clk_i                 ),
        .rst_ni                  ( rst_ni                ),
        .testmode_i              ( testmode_i            ),
        .dmi_rst_ni,
        .dmi_req_valid_i,
        .dmi_req_ready_o,
        .dmi_req_i,
        .dmi_resp_valid_o,
        .dmi_resp_ready_i,
        .dmi_resp_o,
        .ndmreset_o              ( ndmreset_o            ),
        .dmactive_o              ( dmactive_o            ),
        .hartsel_o               ( hartsel               ),
        .hartinfo_i              ( hartinfo_i            ),
        .halted_i                ( halted                ),
        .unavailable_i,
        .resumeack_i             ( resumeack             ),
        .haltreq_o               ( haltreq               ),
        .resumereq_o             ( resumereq             ),
        .clear_resumeack_o       ( clear_resumeack       ),
        .cmd_valid_o             ( cmd_valid             ),
        .cmd_o                   ( cmd                   ),
        .cmderror_valid_i        ( cmderror_valid        ),
        .cmderror_i              ( cmderror              ),
        .cmdbusy_i               ( cmdbusy               ),
        .progbuf_o               ( progbuf               ),
        .data_i                  ( data_mem_csrs         ),
        .data_valid_i            ( data_valid            ),
        .data_o                  ( data_csrs_mem         ),
        .sbaddress_o             ( sbaddress_csrs_sba    ),
        .sbaddress_i             ( sbaddress_sba_csrs    ),
        .sbaddress_write_valid_o ( sbaddress_write_valid ),
        .sbreadonaddr_o          ( sbreadonaddr          ),
        .sbautoincrement_o       ( sbautoincrement       ),
        .sbaccess_o              ( sbaccess              ),
        .sbreadondata_o          ( sbreadondata          ),
        .sbdata_o                ( sbdata_write          ),
        .sbdata_read_valid_o     ( sbdata_read_valid     ),
        .sbdata_write_valid_o    ( sbdata_write_valid    ),
        .sbdata_i                ( sbdata_read           ),
        .sbdata_valid_i          ( sbdata_valid          ),
        .sbbusy_i                ( sbbusy                ),
        .sberror_valid_i         ( sberror_valid         ),
        .sberror_i               ( sberror               )
    );
    dm_sba #(
        .BusWidth(BusWidth)
    ) i_dm_sba (
        .clk_i                   ( clk_i                 ),
        .rst_ni                  ( rst_ni                ),
        .dmactive_i              ( dmactive_o            ),
        .master_req_o            ( master_req_o          ),
        .master_add_o            ( master_add_o          ),
        .master_we_o             ( master_we_o           ),
        .master_wdata_o          ( master_wdata_o        ),
        .master_be_o             ( master_be_o           ),
        .master_gnt_i            ( master_gnt_i          ),
        .master_r_valid_i        ( master_r_valid_i      ),
        .master_r_rdata_i        ( master_r_rdata_i      ),
        .sbaddress_i             ( sbaddress_csrs_sba    ),
        .sbaddress_o             ( sbaddress_sba_csrs    ),
        .sbaddress_write_valid_i ( sbaddress_write_valid ),
        .sbreadonaddr_i          ( sbreadonaddr          ),
        .sbautoincrement_i       ( sbautoincrement       ),
        .sbaccess_i              ( sbaccess              ),
        .sbreadondata_i          ( sbreadondata          ),
        .sbdata_i                ( sbdata_write          ),
        .sbdata_read_valid_i     ( sbdata_read_valid     ),
        .sbdata_write_valid_i    ( sbdata_write_valid    ),
        .sbdata_o                ( sbdata_read           ),
        .sbdata_valid_o          ( sbdata_valid          ),
        .sbbusy_o                ( sbbusy                ),
        .sberror_valid_o         ( sberror_valid         ),
        .sberror_o               ( sberror               )
    );
    dm_mem #(
        .NrHarts(NrHarts),
        .BusWidth(BusWidth),
        .SelectableHarts(SelectableHarts)
    ) i_dm_mem (
        .clk_i                   ( clk_i                 ),
        .rst_ni                  ( rst_ni                ),
        .debug_req_o             ( debug_req_o           ),
        .hartsel_i               ( hartsel               ),
        .haltreq_i               ( haltreq               ),
        .resumereq_i             ( resumereq             ),
        .clear_resumeack_i       ( clear_resumeack       ),
        .halted_o                ( halted                ),
        .resuming_o              ( resumeack             ),
        .cmd_valid_i             ( cmd_valid             ),
        .cmd_i                   ( cmd                   ),
        .cmderror_valid_o        ( cmderror_valid        ),
        .cmderror_o              ( cmderror              ),
        .cmdbusy_o               ( cmdbusy               ),
        .progbuf_i               ( progbuf               ),
        .data_i                  ( data_csrs_mem         ),
        .data_o                  ( data_mem_csrs         ),
        .data_valid_o            ( data_valid            ),
        .req_i                   ( slave_req_i           ),
        .we_i                    ( slave_we_i            ),
        .addr_i                  ( slave_addr_i          ),
        .wdata_i                 ( slave_wdata_i         ),
        .be_i                    ( slave_be_i            ),
        .rdata_o                 ( slave_rdata_o         )
    );
endmodule
module dmi_cdc (
    
    input  logic             tck_i,
    input  logic             trst_ni,
    input  dm::dmi_req_t     jtag_dmi_req_i,
    output logic             jtag_dmi_ready_o,
    input  logic             jtag_dmi_valid_i,
    output dm::dmi_resp_t    jtag_dmi_resp_o,
    output logic             jtag_dmi_valid_o,
    input  logic             jtag_dmi_ready_i,
    
    input  logic             clk_i,
    input  logic             rst_ni,
    output dm::dmi_req_t     core_dmi_req_o,
    output logic             core_dmi_valid_o,
    input  logic             core_dmi_ready_i,
    input dm::dmi_resp_t     core_dmi_resp_i,
    output logic             core_dmi_ready_o,
    input  logic             core_dmi_valid_i
  );
  cdc_2phase #(.T(dm::dmi_req_t)) i_cdc_req (
    .src_rst_ni  ( trst_ni          ),
    .src_clk_i   ( tck_i            ),
    .src_data_i  ( jtag_dmi_req_i   ),
    .src_valid_i ( jtag_dmi_valid_i ),
    .src_ready_o ( jtag_dmi_ready_o ),
    .dst_rst_ni  ( rst_ni           ),
    .dst_clk_i   ( clk_i            ),
    .dst_data_o  ( core_dmi_req_o   ),
    .dst_valid_o ( core_dmi_valid_o ),
    .dst_ready_i ( core_dmi_ready_i )
  );
  cdc_2phase #(.T(dm::dmi_resp_t)) i_cdc_resp (
    .src_rst_ni  ( rst_ni           ),
    .src_clk_i   ( clk_i            ),
    .src_data_i  ( core_dmi_resp_i  ),
    .src_valid_i ( core_dmi_valid_i ),
    .src_ready_o ( core_dmi_ready_o ),
    .dst_rst_ni  ( trst_ni          ),
    .dst_clk_i   ( tck_i            ),
    .dst_data_o  ( jtag_dmi_resp_o  ),
    .dst_valid_o ( jtag_dmi_valid_o ),
    .dst_ready_i ( jtag_dmi_ready_i )
  );
endmodule
module dmi_jtag #(
    parameter logic [31:0] IdcodeValue = 32'h00000001
) (
    input  logic         clk_i,      
    input  logic         rst_ni,     
    input  logic         testmode_i,
    output logic         dmi_rst_no, 
    output dm::dmi_req_t dmi_req_o,
    output logic         dmi_req_valid_o,
    input  logic         dmi_req_ready_i,
    input dm::dmi_resp_t dmi_resp_i,
    output logic         dmi_resp_ready_o,
    input  logic         dmi_resp_valid_i,
    input  logic         tck_i,    
    input  logic         tms_i,    
    input  logic         trst_ni,  
    input  logic         td_i,     
    output logic         td_o,     
    output logic         tdo_oe_o  
);
    assign       dmi_rst_no = rst_ni;
    logic        test_logic_reset;
    logic        shift_dr;
    logic        update_dr;
    logic        capture_dr;
    logic        dmi_access;
    logic        dtmcs_select;
    logic        dmi_reset;
    logic        dmi_tdi;
    logic        dmi_tdo;
    dm::dmi_req_t  dmi_req;
    logic          dmi_req_ready;
    logic          dmi_req_valid;
    dm::dmi_resp_t dmi_resp;
    logic          dmi_resp_valid;
    logic          dmi_resp_ready;
    typedef struct packed {
        logic [6:0]  address;
        logic [31:0] data;
        logic [1:0]  op;
    } dmi_t;
    typedef enum logic [1:0] {
                                DMINoError = 2'h0, DMIReservedError = 2'h1,
                                DMIOPFailed = 2'h2, DMIBusy = 2'h3
                             } dmi_error_e;
    typedef enum logic [2:0] { Idle, Read, WaitReadValid, Write, WaitWriteValid } state_e;
    state_e state_d, state_q;
    logic [$bits(dmi_t)-1:0] dr_d, dr_q;
    logic [6:0] address_d, address_q;
    logic [31:0] data_d, data_q;
    dmi_t  dmi;
    assign dmi          = dmi_t'(dr_q);
    assign dmi_req.addr = address_q;
    assign dmi_req.data = data_q;
    assign dmi_req.op   = (state_q == Write) ? dm::DTM_WRITE : dm::DTM_READ;
    
    assign dmi_resp_ready = 1'b1;
    logic error_dmi_busy;
    dmi_error_e error_d, error_q;
    always_comb begin
        error_dmi_busy = 1'b0;
        
        state_d   = state_q;
        address_d = address_q;
        data_d    = data_q;
        error_d   = error_q;
        dmi_req_valid = 1'b0;
        case (state_q)
            Idle: begin
                
                if (dmi_access && update_dr && (error_q == DMINoError)) begin
                    
                    address_d = dmi.address;
                    data_d = dmi.data;
                    if (dm::dtm_op_e'(dmi.op) == dm::DTM_READ) begin
                        state_d = Read;
                    end else if (dm::dtm_op_e'(dmi.op) == dm::DTM_WRITE) begin
                        state_d = Write;
                    end
                    
                end
            end
            Read: begin
                dmi_req_valid = 1'b1;
                if (dmi_req_ready) begin
                    state_d = WaitReadValid;
                end
            end
            WaitReadValid: begin
                
                if (dmi_resp_valid) begin
                    data_d = dmi_resp.data;
                    state_d = Idle;
                end
            end
            Write: begin
                dmi_req_valid = 1'b1;
                
                if (dmi_req_ready) begin
                    state_d = Idle;
                end
            end
            WaitWriteValid: begin
                
                if (dmi_resp_valid) begin
                    state_d = Idle;
                end
            end
        endcase
        
        
        if (update_dr && state_q != Idle) begin
            error_dmi_busy = 1'b1;
        end
        
        
        
        if (capture_dr && state_q inside {Read, WaitReadValid}) begin
            error_dmi_busy = 1'b1;
        end
        if (error_dmi_busy) begin
            error_d = DMIBusy;
        end
        
        if (dmi_reset && dtmcs_select) begin
            error_d = DMINoError;
        end
    end
    
    assign dmi_tdo = dr_q[0];
    always_comb begin
        dr_d    = dr_q;
        if (capture_dr) begin
            if (dmi_access) begin
                if (error_q == DMINoError && !error_dmi_busy) begin
                    dr_d = {address_q, data_q, DMINoError};
                
                end else if (error_q == DMIBusy || error_dmi_busy) begin
                    dr_d = {address_q, data_q, DMIBusy};
                end
            end
        end
        if (shift_dr) begin
            if (dmi_access) dr_d = {dmi_tdi, dr_q[$bits(dr_q)-1:1]};
        end
        if (test_logic_reset) begin
            dr_d = '0;
        end
    end
    always_ff @(posedge tck_i or negedge trst_ni) begin
        if (!trst_ni) begin
            dr_q      <= '0;
            state_q   <= Idle;
            address_q <= '0;
            data_q    <= '0;
            error_q   <= DMINoError;
        end else begin
            dr_q      <= dr_d;
            state_q   <= state_d;
            address_q <= address_d;
            data_q    <= data_d;
            error_q   <= error_d;
        end
    end
    
    
    
    dmi_jtag_tap #(
        .IrLength (5),
        .IdcodeValue(IdcodeValue)
    ) i_dmi_jtag_tap (
        .tck_i,
        .tms_i,
        .trst_ni,
        .td_i,
        .td_o,
        .tdo_oe_o,
        .testmode_i         ( testmode_i       ),
        .test_logic_reset_o ( test_logic_reset ),
        .shift_dr_o         ( shift_dr         ),
        .update_dr_o        ( update_dr        ),
        .capture_dr_o       ( capture_dr       ),
        .dmi_access_o       ( dmi_access       ),
        .dtmcs_select_o     ( dtmcs_select     ),
        .dmi_reset_o        ( dmi_reset        ),
        .dmi_error_i        ( error_q          ),
        .dmi_tdi_o          ( dmi_tdi          ),
        .dmi_tdo_i          ( dmi_tdo          )
    );
    
    
    
    dmi_cdc i_dmi_cdc (
        
        .tck_i,
        .trst_ni,
        .jtag_dmi_req_i    ( dmi_req          ),
        .jtag_dmi_ready_o  ( dmi_req_ready    ),
        .jtag_dmi_valid_i  ( dmi_req_valid    ),
        .jtag_dmi_resp_o   ( dmi_resp         ),
        .jtag_dmi_valid_o  ( dmi_resp_valid   ),
        .jtag_dmi_ready_i  ( dmi_resp_ready   ),
        
        .clk_i,
        .rst_ni,
        .core_dmi_req_o    ( dmi_req_o        ),
        .core_dmi_valid_o  ( dmi_req_valid_o  ),
        .core_dmi_ready_i  ( dmi_req_ready_i  ),
        .core_dmi_resp_i   ( dmi_resp_i       ),
        .core_dmi_ready_o  ( dmi_resp_ready_o ),
        .core_dmi_valid_i  ( dmi_resp_valid_i )
    );
endmodule
module dm_sba #(
    parameter int BusWidth = -1
) (
    input  logic                   clk_i,       
    input  logic                   rst_ni,
    input  logic                   dmactive_i,  
    output logic                   master_req_o,
    output logic [BusWidth-1:0]    master_add_o,
    output logic                   master_we_o,
    output logic [BusWidth-1:0]    master_wdata_o,
    output logic [BusWidth/8-1:0]  master_be_o,
    input  logic                   master_gnt_i,
    input  logic                   master_r_valid_i,
    input  logic [BusWidth-1:0]    master_r_rdata_i,
    input  logic [BusWidth-1:0]    sbaddress_i,
    input  logic                   sbaddress_write_valid_i,
    
    input  logic                   sbreadonaddr_i,
    output logic [BusWidth-1:0]    sbaddress_o,
    input  logic                   sbautoincrement_i,
    input  logic [2:0]             sbaccess_i,
    
    input  logic                   sbreadondata_i,
    input  logic [BusWidth-1:0]    sbdata_i,
    input  logic                   sbdata_read_valid_i,
    input  logic                   sbdata_write_valid_i,
    
    output logic [BusWidth-1:0]    sbdata_o,
    output logic                   sbdata_valid_o,
    
    output logic                   sbbusy_o,
    output logic                   sberror_valid_o, 
    output logic [2:0]             sberror_o 
);
    typedef enum logic [2:0] { Idle, Read, Write, WaitRead, WaitWrite } state_e;
    state_e state_d, state_q;
    logic [BusWidth-1:0]   address;
    logic                  req;
    logic                  gnt;
    logic                  we;
    logic [BusWidth/8-1:0] be;
    assign sbbusy_o = (state_q != Idle) ? 1'b1 : 1'b0;
    always_comb begin
        req     = 1'b0;
        address = sbaddress_i;
        we      = 1'b0;
        be      = '0;
        sberror_o       = '0;
        sberror_valid_o = 1'b0;
        sbaddress_o     = sbaddress_i;
        state_d = state_q;
        case (state_q)
            Idle: begin
                
                if (sbaddress_write_valid_i && sbreadonaddr_i)  state_d = Read;
                
                if (sbdata_write_valid_i) state_d = Write;
                
                if (sbdata_read_valid_i && sbreadondata_i) state_d = Read;
            end
            Read: begin
                req = 1'b1;
                if (gnt) state_d = WaitRead;
            end
            Write: begin
                req = 1'b1;
                we  = 1'b1;
                
                case (sbaccess_i)
                    3'b000: begin
                        if (BusWidth == 64) be[ sbaddress_i[2:0]] = '1;
                        else                be[ sbaddress_i[1:0]] = '1;
                    end
                    3'b001: begin
                        if (BusWidth == 64) be[{sbaddress_i[2:1], 1'b0} +: 2] = '1;
                        else                be[{sbaddress_i[1:1], 1'b0} +: 2] = '1;
                    end
                    3'b010: begin
                        if (BusWidth == 64) be[{sbaddress_i[2:2], 2'b0} +: 4] = '1;
                        else                be = '1;
                    end
                    3'b011: be = '1;
                    default:;
                endcase
                if (gnt) state_d = WaitWrite;
            end
            WaitRead: begin
                if (sbdata_valid_o) begin
                    state_d = Idle;
                    
                    if (sbautoincrement_i) sbaddress_o = sbaddress_i + (1'b1 << sbaccess_i);
                end
            end
            WaitWrite: begin
                if (sbdata_valid_o) begin
                    state_d = Idle;
                    
                    if (sbautoincrement_i) sbaddress_o = sbaddress_i + (1'b1 << sbaccess_i);
                end
            end
            default:;
        endcase
        
        if (sbaccess_i > 3 && state_q != Idle) begin
            req             = 1'b0;
            state_d         = Idle;
            sberror_valid_o = 1'b1;
            sberror_o       = 3'd3;
        end
        
    end
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (!rst_ni) begin
            state_q <= Idle;
        end else begin
            state_q <= state_d;
        end
    end
    assign master_req_o    = req;
    assign master_add_o    = address[BusWidth-1:0];
    assign master_we_o     = we;
    assign master_wdata_o  = sbdata_i[BusWidth-1:0];
    assign master_be_o     = be[BusWidth/8-1:0];
    assign gnt             = master_gnt_i;
    assign sbdata_valid_o  = master_r_valid_i;
    assign sbdata_o        = master_r_rdata_i[BusWidth-1:0];
    
    
    
    
endmodule
module dmi_jtag_tap #(
    parameter int IrLength = 5,
    
    parameter logic [31:0] IdcodeValue = 32'h00000001
    
    
    
    
)(
    input  logic        tck_i,    
    input  logic        tms_i,    
    input  logic        trst_ni,  
    input  logic        td_i,     
    output logic        td_o,     
    output logic        tdo_oe_o, 
    input  logic        testmode_i,
    output logic        test_logic_reset_o,
    output logic        shift_dr_o,
    output logic        update_dr_o,
    output logic        capture_dr_o,
    
    output logic        dmi_access_o,
    
    output logic        dtmcs_select_o,
    
    output logic        dmi_reset_o,
    input  logic [1:0]  dmi_error_i,
    
    output logic        dmi_tdi_o,
    
    input  logic        dmi_tdo_i
);
    
    assign dmi_tdi_o = td_i;
    typedef enum logic [3:0] { TestLogicReset, RunTestIdle, SelectDrScan,
                     CaptureDr, ShiftDr, Exit1Dr, PauseDr, Exit2Dr,
                     UpdateDr, SelectIrScan, CaptureIr, ShiftIr,
                     Exit1Ir, PauseIr, Exit2Ir, UpdateIr } tap_state_e;
    tap_state_e tap_state_q, tap_state_d;
    typedef enum logic [IrLength-1:0] {
        BYPASS0   = 'h0,
        IDCODE    = 'h1,
        DTMCSR    = 'h10,
        DMIACCESS = 'h11,
        BYPASS1   = 'h1f
    } ir_reg_e;
    typedef struct packed {
        logic [31:18] zero1;
        logic         dmihardreset;
        logic         dmireset;
        logic         zero0;
        logic [14:12] idle;
        logic [11:10] dmistat;
        logic [9:4]   abits;
        logic [3:0]   version;
    } dtmcs_t;
    
    
    
    logic [IrLength-1:0]  jtag_ir_shift_d, jtag_ir_shift_q; 
    ir_reg_e              jtag_ir_d, jtag_ir_q; 
    logic capture_ir, shift_ir, pause_ir, update_ir;
    always_comb begin
        jtag_ir_shift_d = jtag_ir_shift_q;
        jtag_ir_d       = jtag_ir_q;
        
        if (shift_ir) begin
            jtag_ir_shift_d = {td_i, jtag_ir_shift_q[IrLength-1:1]};
        end
        
        if (capture_ir) begin
            jtag_ir_shift_d =  'b0101;
        end
        
        if (update_ir) begin
            jtag_ir_d = ir_reg_e'(jtag_ir_shift_q);
        end
        
        if (test_logic_reset_o) begin
            jtag_ir_shift_d = '0;
            jtag_ir_d       = IDCODE;
        end
    end
    always_ff @(posedge tck_i, negedge trst_ni) begin
        if (!trst_ni) begin
            jtag_ir_shift_q <= '0;
            jtag_ir_q       <= IDCODE;
        end else begin
            jtag_ir_shift_q <= jtag_ir_shift_d;
            jtag_ir_q       <= jtag_ir_d;
        end
    end
    
    
    
    
    
    
    logic [31:0] idcode_d, idcode_q;
    logic        idcode_select;
    logic        bypass_select;
    dtmcs_t      dtmcs_d, dtmcs_q;
    logic        bypass_d, bypass_q;  
    assign dmi_reset_o = dtmcs_q.dmireset;
    always_comb begin
        idcode_d = idcode_q;
        bypass_d = bypass_q;
        dtmcs_d  = dtmcs_q;
        if (capture_dr_o) begin
            if (idcode_select) idcode_d = IdcodeValue;
            if (bypass_select) bypass_d = 1'b0;
            if (dtmcs_select_o) begin
                dtmcs_d  = '{
                                zero1        : '0,
                                dmihardreset : 1'b0,
                                dmireset     : 1'b0,
                                zero0        : '0,
                                idle         : 'd1,         
                                dmistat      : dmi_error_i, 
                                abits        : 'd7, 
                                version      : 'd1  
                            };
            end
        end
        if (shift_dr_o) begin
            if (idcode_select)  idcode_d = {td_i, idcode_q[31:1]};
            if (bypass_select)  bypass_d = td_i;
            if (dtmcs_select_o) dtmcs_d  = {td_i, dtmcs_q[31:1]};
        end
        if (test_logic_reset_o) begin
            idcode_d = IdcodeValue;
            bypass_d = 1'b0;
        end
    end
    
    
    
    always_comb begin
        dmi_access_o   = 1'b0;
        dtmcs_select_o = 1'b0;
        idcode_select  = 1'b0;
        bypass_select  = 1'b0;
        case (jtag_ir_q)
            BYPASS0:   bypass_select  = 1'b1;
            IDCODE:    idcode_select  = 1'b1;
            DTMCSR:    dtmcs_select_o = 1'b1;
            DMIACCESS: dmi_access_o   = 1'b1;
            BYPASS1:   bypass_select  = 1'b1;
            default:   bypass_select  = 1'b1;
        endcase
    end
    
    
    
    logic tdo_mux;
    always_comb begin
        
        if (shift_ir) begin
            tdo_mux = jtag_ir_shift_q[0];
        
        end else begin
          case (jtag_ir_q)    
            IDCODE:         tdo_mux = idcode_q[0];     
            DTMCSR:         tdo_mux = dtmcs_q[0];
            DMIACCESS:      tdo_mux = dmi_tdo_i;       
            default:        tdo_mux = bypass_q;      
          endcase
        end
    end
    
    logic tck_n, tck_ni;
    cluster_clock_inverter i_tck_inv (
        .clk_i ( tck_i  ),
        .clk_o ( tck_ni )
    );
    pulp_clock_mux2 i_dft_tck_mux (
        .clk0_i    ( tck_ni     ),
        .clk1_i    ( tck_i      ), 
        .clk_sel_i ( testmode_i ),
        .clk_o     ( tck_n      )
    );
    
    always_ff @(posedge tck_n, negedge trst_ni) begin
        if (!trst_ni) begin
            td_o     <= 1'b0;
            tdo_oe_o <= 1'b0;
        end else begin
            td_o     <= tdo_mux;
            tdo_oe_o <= (shift_ir | shift_dr_o);
        end
    end
    
    
    
    
    always_comb begin
        test_logic_reset_o = 1'b0;
        capture_dr_o       = 1'b0;
        shift_dr_o         = 1'b0;
        update_dr_o        = 1'b0;
        capture_ir         = 1'b0;
        shift_ir           = 1'b0;
        pause_ir           = 1'b0;
        update_ir          = 1'b0;
        case (tap_state_q)
            TestLogicReset: begin
                tap_state_d = (tms_i) ? TestLogicReset : RunTestIdle;
                test_logic_reset_o = 1'b1;
            end
            RunTestIdle: begin
                tap_state_d = (tms_i) ? SelectDrScan : RunTestIdle;
            end
            
            SelectDrScan: begin
                tap_state_d = (tms_i) ? SelectIrScan : CaptureDr;
            end
            CaptureDr: begin
                capture_dr_o = 1'b1;
                tap_state_d = (tms_i) ? Exit1Dr : ShiftDr;
            end
            ShiftDr: begin
                shift_dr_o = 1'b1;
                tap_state_d = (tms_i) ? Exit1Dr : ShiftDr;
            end
            Exit1Dr: begin
                tap_state_d = (tms_i) ? UpdateDr : PauseDr;
            end
            PauseDr: begin
                tap_state_d = (tms_i) ? Exit2Dr : PauseDr;
            end
            Exit2Dr: begin
                tap_state_d = (tms_i) ? UpdateDr : ShiftDr;
            end
            UpdateDr: begin
                update_dr_o = 1'b1;
                tap_state_d = (tms_i) ? SelectDrScan : RunTestIdle;
            end
            
            SelectIrScan: begin
                tap_state_d = (tms_i) ? TestLogicReset : CaptureIr;
            end
            
            
            
            
            CaptureIr: begin
                capture_ir = 1'b1;
                tap_state_d = (tms_i) ? Exit1Ir : ShiftIr;
            end
            
            
            
            
            ShiftIr: begin
                shift_ir = 1'b1;
                tap_state_d = (tms_i) ? Exit1Ir : ShiftIr;
            end
            Exit1Ir: begin
                tap_state_d = (tms_i) ? UpdateIr : PauseIr;
            end
            PauseIr: begin
                pause_ir = 1'b1;
                tap_state_d = (tms_i) ? Exit2Ir : PauseIr;
            end
            Exit2Ir: begin
                tap_state_d = (tms_i) ? UpdateIr : ShiftIr;
            end
            
            
            
            
            UpdateIr: begin
                update_ir = 1'b1;
                tap_state_d = (tms_i) ? SelectDrScan : RunTestIdle;
            end
            default: tap_state_d = TestLogicReset;  
      endcase
    end
    always_ff @(posedge tck_i or negedge trst_ni) begin
        if (!trst_ni) begin
            tap_state_q <= RunTestIdle;
            idcode_q    <= IdcodeValue;
            bypass_q    <= 1'b0;
            dtmcs_q     <= '0;
        end else begin
            tap_state_q <= tap_state_d;
            idcode_q    <= idcode_d;
            bypass_q    <= bypass_d;
            dtmcs_q     <= dtmcs_d;
        end
    end
endmodule
module debug_rom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 19;
    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_7b200073,
        64'h7b302573_7b202473,
        64'h10852423_f1402473,
        64'ha85ff06f_7b302573,
        64'h7b202473_10052223,
        64'h00100073_7b302573,
        64'h10052623_00c51513,
        64'h00c55513_00000517,
        64'h7b351073_fd5ff06f,
        64'hfa041ce3_00247413,
        64'h40044403_00a40433,
        64'hf1402473_02041c63,
        64'h00147413_40044403,
        64'h00a40433_10852023,
        64'hf1402473_00c51513,
        64'h00c55513_00000517,
        64'h7b351073_7b241073,
        64'h0ff0000f_04c0006f,
        64'h07c0006f_00c0006f
    };
    logic [$clog2(RomSize)-1:0] addr_q;
    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end
    
    
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
module ariane_verilog_wrap
    import ariane_pkg::*;
#(
  parameter int unsigned               RASDepth              = 2,
  parameter int unsigned               BTBEntries            = 32,
  parameter int unsigned               BHTEntries            = 128,
  
  parameter logic [63:0]               DmBaseAddress         = 64'h0,
  
  parameter bit                        SwapEndianess         = 1,
  
  
  parameter int unsigned               NrNonIdempotentRules  =  1,
  parameter logic [NrMaxRules*64-1:0]  NonIdempotentAddrBase = 64'h00C0000000,
  parameter logic [NrMaxRules*64-1:0]  NonIdempotentLength   = 64'hFFFFFFFFFF,
  
  parameter int unsigned               NrExecuteRegionRules  =  0,
  parameter logic [NrMaxRules*64-1:0]  ExecuteRegionAddrBase = '0,
  parameter logic [NrMaxRules*64-1:0]  ExecuteRegionLength   = '0,
  
  parameter int unsigned               NrCachedRegionRules   =  0,
  parameter logic [NrMaxRules*64-1:0]  CachedRegionAddrBase  = '0,
  parameter logic [NrMaxRules*64-1:0]  CachedRegionLength    = '0,
  
  parameter int unsigned               NrPMPEntries          =  8
) (
  input                       clk_i,
  input                       reset_l,      
  output                      spc_grst_l,   
  
  input  [riscv::VLEN-1:0]               boot_addr_i,  
  input  [riscv::XLEN-1:0]               hart_id_i,    
  
  input  [1:0]                irq_i,        
  input                       ipi_i,        
  
  input                       time_irq_i,   
  input                       debug_req_i,  
  
  output [$size(wt_cache_pkg::l15_req_t)-1:0]  l15_req_o,
  input  [$size(wt_cache_pkg::l15_rtrn_t)-1:0] l15_rtrn_i
 );
  
  wt_cache_pkg::l15_req_t  l15_req;
  wt_cache_pkg::l15_rtrn_t l15_rtrn;
  assign l15_req_o = l15_req;
  assign l15_rtrn  = l15_rtrn_i;
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  logic [15:0] wake_up_cnt_d, wake_up_cnt_q;
  logic rst_n;
  assign wake_up_cnt_d = (wake_up_cnt_q[$high(wake_up_cnt_q)]) ? wake_up_cnt_q : wake_up_cnt_q + 1;
  always_ff @(posedge clk_i or negedge reset_l) begin : p_regs
    if(~reset_l) begin
      wake_up_cnt_q <= 0;
    end else begin
      wake_up_cnt_q <= wake_up_cnt_d;
    end
  end
  
  assign rst_n = wake_up_cnt_q[$high(wake_up_cnt_q)] & reset_l;
  
  
  
  logic [1:0] irq;
  logic ipi, time_irq, debug_req;
  
  synchronizer i_sync (
    .clk         ( clk_i      ),
    .presyncdata ( rst_n      ),
    .syncdata    ( spc_grst_l )
  );
  
  for (genvar k=0; k<$size(irq_i); k++) begin
    synchronizer i_irq_sync (
      .clk         ( clk_i      ),
      .presyncdata ( irq_i[k]   ),
      .syncdata    ( irq[k]     )
    );
  end
  synchronizer i_ipi_sync (
    .clk         ( clk_i      ),
    .presyncdata ( ipi_i      ),
    .syncdata    ( ipi        )
  );
  synchronizer i_timer_sync (
    .clk         ( clk_i      ),
    .presyncdata ( time_irq_i ),
    .syncdata    ( time_irq   )
  );
  synchronizer i_debug_sync (
    .clk         ( clk_i       ),
    .presyncdata ( debug_req_i ),
    .syncdata    ( debug_req   )
  );
  
  
  
  localparam ariane_pkg::ariane_cfg_t ArianeOpenPitonCfg = '{
    RASDepth:              RASDepth,
    BTBEntries:            BTBEntries,
    BHTEntries:            BHTEntries,
    
    NrNonIdempotentRules:  NrNonIdempotentRules,
    NonIdempotentAddrBase: NonIdempotentAddrBase,
    NonIdempotentLength:   NonIdempotentLength,
    NrExecuteRegionRules:  NrExecuteRegionRules,
    ExecuteRegionAddrBase: ExecuteRegionAddrBase,
    ExecuteRegionLength:   ExecuteRegionLength,
    
    NrCachedRegionRules:   NrCachedRegionRules,
    CachedRegionAddrBase:  CachedRegionAddrBase,
    CachedRegionLength:    CachedRegionLength,
    
    Axi64BitCompliant:     1'b0,
    SwapEndianess:         SwapEndianess,
    
    DmBaseAddress:         DmBaseAddress,
    NrPMPEntries:          NrPMPEntries
  };
  ariane #(
    .ArianeCfg ( ArianeOpenPitonCfg )
  ) ariane (
    .clk_i       ( clk_i      ),
    .rst_ni      ( spc_grst_l ),
    .boot_addr_i              ,
    .hart_id_i                ,
    .irq_i       ( irq        ),
    .ipi_i       ( ipi        ),
    .time_irq_i  ( time_irq   ),
    .debug_req_i ( debug_req  ),
    .l15_req_o   ( l15_req   ),
    .l15_rtrn_i  ( l15_rtrn  )
  );
endmodule 
module riscv_peripherals #(
    parameter int unsigned DataWidth       = 64,
    parameter int unsigned NumHarts        =  1,
    parameter int unsigned NumSources      =  1,
    parameter int unsigned PlicMaxPriority =  7,
    parameter bit          SwapEndianess   =  0,
    parameter logic [63:0] DmBase          = 64'hfff1000000,
    parameter logic [63:0] RomBase         = 64'hfff1010000,
    parameter logic [63:0] ClintBase       = 64'hfff1020000,
    parameter logic [63:0] PlicBase        = 64'hfff1100000
) (
    input                               clk_i,
    input                               rst_ni,
    input                               testmode_i,
    
    
    input  [DataWidth-1:0]              buf_ariane_debug_noc2_data_i,
    input                               buf_ariane_debug_noc2_valid_i,
    output                              ariane_debug_buf_noc2_ready_o,
    output [DataWidth-1:0]              ariane_debug_buf_noc3_data_o,
    output                              ariane_debug_buf_noc3_valid_o,
    input                               buf_ariane_debug_noc3_ready_i,
    
    input  [DataWidth-1:0]              buf_ariane_bootrom_noc2_data_i,
    input                               buf_ariane_bootrom_noc2_valid_i,
    output                              ariane_bootrom_buf_noc2_ready_o,
    output [DataWidth-1:0]              ariane_bootrom_buf_noc3_data_o,
    output                              ariane_bootrom_buf_noc3_valid_o,
    input                               buf_ariane_bootrom_noc3_ready_i,
    
    input  [DataWidth-1:0]              buf_ariane_clint_noc2_data_i,
    input                               buf_ariane_clint_noc2_valid_i,
    output                              ariane_clint_buf_noc2_ready_o,
    output [DataWidth-1:0]              ariane_clint_buf_noc3_data_o,
    output                              ariane_clint_buf_noc3_valid_o,
    input                               buf_ariane_clint_noc3_ready_i,
    
    input [DataWidth-1:0]               buf_ariane_plic_noc2_data_i,
    input                               buf_ariane_plic_noc2_valid_i,
    output                              ariane_plic_buf_noc2_ready_o,
    output [DataWidth-1:0]              ariane_plic_buf_noc3_data_o,
    output                              ariane_plic_buf_noc3_valid_o,
    input                               buf_ariane_plic_noc3_ready_i,
    
    input                               ariane_boot_sel_i,
    
    output                              ndmreset_o,    
    output                              dmactive_o,    
    output [NumHarts-1:0]               debug_req_o,   
    input  [NumHarts-1:0]               unavailable_i, 
    
    input                               tck_i,
    input                               tms_i,
    input                               trst_ni,
    input                               td_i,
    output                              td_o,
    output                              tdo_oe_o,
    
    input                               rtc_i,        
    output [NumHarts-1:0]               timer_irq_o,  
    output [NumHarts-1:0]               ipi_o,        
    
    input  [NumSources-1:0]             irq_sources_i,
    input  [NumSources-1:0]             irq_le_i,     
    output [NumHarts-1:0][1:0]          irq_o         
);
  localparam int unsigned AxiIdWidth    =  1;
  localparam int unsigned AxiAddrWidth  = 64;
  localparam int unsigned AxiDataWidth  = 64;
  localparam int unsigned AxiUserWidth  =  1;
  
  
  
  logic          debug_req_valid;
  logic          debug_req_ready;
  logic          debug_resp_valid;
  logic          debug_resp_ready;
  dm::dmi_req_t  debug_req;
  dm::dmi_resp_t debug_resp;
 
  logic        tck, tms, trst_n, tdi, tdo, tdo_oe;
  dmi_jtag i_dmi_jtag (
    .clk_i                                ,
    .rst_ni                               ,
    .testmode_i                           ,
    .dmi_req_o        ( debug_req        ),
    .dmi_req_valid_o  ( debug_req_valid  ),
    .dmi_req_ready_i  ( debug_req_ready  ),
    .dmi_resp_i       ( debug_resp       ),
    .dmi_resp_ready_o ( debug_resp_ready ),
    .dmi_resp_valid_i ( debug_resp_valid ),
    .dmi_rst_no       (                  ), 
    .tck_i            ( tck              ),
    .tms_i            ( tms              ),
    .trst_ni          ( trst_n           ),
    .td_i             ( tdi              ),
    .td_o             ( tdo              ),
    .tdo_oe_o         ( tdo_oe           )
  );
 
  assign tck      = tck_i   ;
  assign tms      = tms_i   ;
  assign trst_n   = trst_ni ;
  assign tdi      = td_i    ;
  assign td_o     = tdo     ;
  assign tdo_oe_o = tdo_oe  ;
 
 
  logic                dm_slave_req;
  logic                dm_slave_we;
  logic [64-1:0]       dm_slave_addr;
  logic [64/8-1:0]     dm_slave_be;
  logic [64-1:0]       dm_slave_wdata;
  logic [64-1:0]       dm_slave_rdata;
  logic                dm_master_req;
  logic [64-1:0]       dm_master_add;
  logic                dm_master_we;
  logic [64-1:0]       dm_master_wdata;
  logic [64/8-1:0]     dm_master_be;
  logic                dm_master_gnt;
  logic                dm_master_r_valid;
  logic [64-1:0]       dm_master_r_rdata;
  
  dm_top #(
    .NrHarts              ( NumHarts             ),
    .BusWidth             ( AxiDataWidth         ),
    .SelectableHarts      ( {NumHarts{1'b1}}     )
  ) i_dm_top (
    .clk_i                                        ,
    .rst_ni                                       , 
    .testmode_i                                   ,
    .ndmreset_o                                   ,
    .dmactive_o                                   , 
    .debug_req_o                                  ,
    .unavailable_i                                ,
    .hartinfo_i           ( {NumHarts{ariane_pkg::DebugHartInfo}} ),
    .slave_req_i          ( dm_slave_req         ),
    .slave_we_i           ( dm_slave_we          ),
    .slave_addr_i         ( dm_slave_addr        ),
    .slave_be_i           ( dm_slave_be          ),
    .slave_wdata_i        ( dm_slave_wdata       ),
    .slave_rdata_o        ( dm_slave_rdata       ),
    .master_req_o         ( dm_master_req        ),
    .master_add_o         ( dm_master_add        ),
    .master_we_o          ( dm_master_we         ),
    .master_wdata_o       ( dm_master_wdata      ),
    .master_be_o          ( dm_master_be         ),
    .master_gnt_i         ( dm_master_gnt        ),
    .master_r_valid_i     ( dm_master_r_valid    ),
    .master_r_rdata_i     ( dm_master_r_rdata    ),
    .dmi_rst_ni           ( rst_ni               ),
    .dmi_req_valid_i      ( debug_req_valid      ),
    .dmi_req_ready_o      ( debug_req_ready      ),
    .dmi_req_i            ( debug_req            ),
    .dmi_resp_valid_o     ( debug_resp_valid     ),
    .dmi_resp_ready_i     ( debug_resp_ready     ),
    .dmi_resp_o           ( debug_resp           )
  );
  AXI_BUS #(
      .AXI_ADDR_WIDTH ( AxiAddrWidth     ),
      .AXI_DATA_WIDTH ( AxiDataWidth     ),
      .AXI_ID_WIDTH   ( AxiIdWidth       ),
      .AXI_USER_WIDTH ( AxiUserWidth     )
  ) dm_master();
  axi2mem #(
      .AXI_ID_WIDTH   ( AxiIdWidth   ),
      .AXI_ADDR_WIDTH ( AxiAddrWidth ),
      .AXI_DATA_WIDTH ( AxiDataWidth ),
      .AXI_USER_WIDTH ( AxiUserWidth )
  ) i_dm_axi2mem (
      .clk_i      ( clk_i                     ),
      .rst_ni     ( rst_ni                    ),
      .slave      ( dm_master                 ),
      .req_o      ( dm_slave_req              ),
      .we_o       ( dm_slave_we               ),
      .addr_o     ( dm_slave_addr             ),
      .be_o       ( dm_slave_be               ),
      .data_o     ( dm_slave_wdata            ),
      .data_i     ( dm_slave_rdata            )
  );
  noc_axilite_bridge #(
    .SLAVE_RESP_BYTEWIDTH   ( 8             ),
    .SWAP_ENDIANESS         ( SwapEndianess )
  ) i_debug_axilite_bridge (
    .clk                    ( clk_i                         ),
    .rst                    ( ~rst_ni                       ),
    
    .splitter_bridge_val    ( buf_ariane_debug_noc2_valid_i ),
    .splitter_bridge_data   ( buf_ariane_debug_noc2_data_i  ),
    .bridge_splitter_rdy    ( ariane_debug_buf_noc2_ready_o ),
    .bridge_splitter_val    ( ariane_debug_buf_noc3_valid_o ),
    .bridge_splitter_data   ( ariane_debug_buf_noc3_data_o  ),
    .splitter_bridge_rdy    ( buf_ariane_debug_noc3_ready_i ),
    
    
    .m_axi_awaddr           ( dm_master.aw_addr             ),
    .m_axi_awvalid          ( dm_master.aw_valid            ),
    .m_axi_awready          ( dm_master.aw_ready            ),
    
    .m_axi_wdata            ( dm_master.w_data              ),
    .m_axi_wstrb            ( dm_master.w_strb              ),
    .m_axi_wvalid           ( dm_master.w_valid             ),
    .m_axi_wready           ( dm_master.w_ready             ),
    
    .m_axi_araddr           ( dm_master.ar_addr             ),
    .m_axi_arvalid          ( dm_master.ar_valid            ),
    .m_axi_arready          ( dm_master.ar_ready            ),
    
    .m_axi_rdata            ( dm_master.r_data              ),
    .m_axi_rresp            ( dm_master.r_resp              ),
    .m_axi_rvalid           ( dm_master.r_valid             ),
    .m_axi_rready           ( dm_master.r_ready             ),
    
    .m_axi_bresp            ( dm_master.b_resp              ),
    .m_axi_bvalid           ( dm_master.b_valid             ),
    .m_axi_bready           ( dm_master.b_ready             ),
    
    .w_reqbuf_size          (                               ),
    .r_reqbuf_size          (                               )
  );
  
  
  assign dm_master_gnt      = '0;
  assign dm_master_r_valid  = '0;
  assign dm_master_r_rdata  = '0;
  
  assign dm_master.aw_id     = '0;
  assign dm_master.aw_len    = '0;
  assign dm_master.aw_size   = 3'b11;
  assign dm_master.aw_burst  = '0;
  assign dm_master.aw_lock   = '0;
  assign dm_master.aw_cache  = '0;
  assign dm_master.aw_prot   = '0;
  assign dm_master.aw_qos    = '0;
  assign dm_master.aw_region = '0;
  assign dm_master.aw_atop   = '0;
  assign dm_master.w_last    = 1'b1;
  assign dm_master.ar_id     = '0;
  assign dm_master.ar_len    = '0;
  assign dm_master.ar_size   = 3'b11;
  assign dm_master.ar_burst  = '0;
  assign dm_master.ar_lock   = '0;
  assign dm_master.ar_cache  = '0;
  assign dm_master.ar_prot   = '0;
  assign dm_master.ar_qos    = '0;
  assign dm_master.ar_region = '0;
  
  
  
  logic                    rom_req;
  logic [AxiAddrWidth-1:0] rom_addr;
  logic [AxiDataWidth-1:0] rom_rdata, rom_rdata_bm, rom_rdata_linux;
  AXI_BUS #(
    .AXI_ID_WIDTH   ( AxiIdWidth   ),
    .AXI_ADDR_WIDTH ( AxiAddrWidth ),
    .AXI_DATA_WIDTH ( AxiDataWidth ),
    .AXI_USER_WIDTH ( AxiUserWidth )
  ) br_master();
  axi2mem #(
    .AXI_ID_WIDTH   ( AxiIdWidth    ),
    .AXI_ADDR_WIDTH ( AxiAddrWidth  ),
    .AXI_DATA_WIDTH ( AxiDataWidth  ),
    .AXI_USER_WIDTH ( AxiUserWidth  )
  ) i_axi2rom (
    .clk_i                ,
    .rst_ni               ,
    .slave  ( br_master  ),
    .req_o  ( rom_req    ),
    .we_o   (            ),
    .addr_o ( rom_addr   ),
    .be_o   (            ),
    .data_o (            ),
    .data_i ( rom_rdata  )
  );
  bootrom i_bootrom_bm (
    .clk_i                   ,
    .req_i      ( rom_req   ),
    .addr_i     ( rom_addr  ),
    .rdata_o    ( rom_rdata_bm )
  );
  bootrom_linux i_bootrom_linux (
    .clk_i                   ,
    .req_i      ( rom_req   ),
    .addr_i     ( rom_addr  ),
    .rdata_o    ( rom_rdata_linux )
  );
  
  assign rom_rdata = (ariane_boot_sel_i) ? rom_rdata_bm : rom_rdata_linux;
  noc_axilite_bridge #(
    .SLAVE_RESP_BYTEWIDTH   ( 8             ),
    .SWAP_ENDIANESS         ( SwapEndianess )
  ) i_bootrom_axilite_bridge (
    .clk                    ( clk_i                           ),
    .rst                    ( ~rst_ni                         ),
    
    .splitter_bridge_val    ( buf_ariane_bootrom_noc2_valid_i ),
    .splitter_bridge_data   ( buf_ariane_bootrom_noc2_data_i  ),
    .bridge_splitter_rdy    ( ariane_bootrom_buf_noc2_ready_o ),
    .bridge_splitter_val    ( ariane_bootrom_buf_noc3_valid_o ),
    .bridge_splitter_data   ( ariane_bootrom_buf_noc3_data_o  ),
    .splitter_bridge_rdy    ( buf_ariane_bootrom_noc3_ready_i ),
    
    
    .m_axi_awaddr           ( br_master.aw_addr               ),
    .m_axi_awvalid          ( br_master.aw_valid              ),
    .m_axi_awready          ( br_master.aw_ready              ),
    
    .m_axi_wdata            ( br_master.w_data                ),
    .m_axi_wstrb            ( br_master.w_strb                ),
    .m_axi_wvalid           ( br_master.w_valid               ),
    .m_axi_wready           ( br_master.w_ready               ),
    
    .m_axi_araddr           ( br_master.ar_addr               ),
    .m_axi_arvalid          ( br_master.ar_valid              ),
    .m_axi_arready          ( br_master.ar_ready              ),
    
    .m_axi_rdata            ( br_master.r_data                ),
    .m_axi_rresp            ( br_master.r_resp                ),
    .m_axi_rvalid           ( br_master.r_valid               ),
    .m_axi_rready           ( br_master.r_ready               ),
    
    .m_axi_bresp            ( br_master.b_resp                ),
    .m_axi_bvalid           ( br_master.b_valid               ),
    .m_axi_bready           ( br_master.b_ready               ),
    
    .w_reqbuf_size          (                                 ),
    .r_reqbuf_size          (                                 )
  );
  
  assign br_master.aw_id     = '0;
  assign br_master.aw_len    = '0;
  assign br_master.aw_size   = 3'b11;
  assign br_master.aw_burst  = '0;
  assign br_master.aw_lock   = '0;
  assign br_master.aw_cache  = '0;
  assign br_master.aw_prot   = '0;
  assign br_master.aw_qos    = '0;
  assign br_master.aw_region = '0;
  assign br_master.aw_atop   = '0;
  assign br_master.w_last    = 1'b1;
  assign br_master.ar_id     = '0;
  assign br_master.ar_len    = '0;
  assign br_master.ar_size   = 3'b11;
  assign br_master.ar_burst  = '0;
  assign br_master.ar_lock   = '0;
  assign br_master.ar_cache  = '0;
  assign br_master.ar_prot   = '0;
  assign br_master.ar_qos    = '0;
  assign br_master.ar_region = '0;
  
  
  
  ariane_axi::req_t    clint_axi_req;
  ariane_axi::resp_t   clint_axi_resp;
  clint #(
    .AXI_ADDR_WIDTH ( AxiAddrWidth ),
    .AXI_DATA_WIDTH ( AxiDataWidth ),
    .AXI_ID_WIDTH   ( AxiIdWidth   ),
    .NR_CORES       ( NumHarts     )
  ) i_clint (
    .clk_i                         ,
    .rst_ni                        ,
    .testmode_i                    ,
    .axi_req_i   ( clint_axi_req  ),
    .axi_resp_o  ( clint_axi_resp ),
    .rtc_i                         ,
    .timer_irq_o                   ,
    .ipi_o
  );
  noc_axilite_bridge #(
    .SLAVE_RESP_BYTEWIDTH   ( 8             ),
    .SWAP_ENDIANESS         ( SwapEndianess )
  ) i_clint_axilite_bridge (
    .clk                    ( clk_i                         ),
    .rst                    ( ~rst_ni                       ),
    
    .splitter_bridge_val    ( buf_ariane_clint_noc2_valid_i ),
    .splitter_bridge_data   ( buf_ariane_clint_noc2_data_i  ),
    .bridge_splitter_rdy    ( ariane_clint_buf_noc2_ready_o ),
    .bridge_splitter_val    ( ariane_clint_buf_noc3_valid_o ),
    .bridge_splitter_data   ( ariane_clint_buf_noc3_data_o  ),
    .splitter_bridge_rdy    ( buf_ariane_clint_noc3_ready_i ),
    
    
    .m_axi_awaddr           ( clint_axi_req.aw.addr         ),
    .m_axi_awvalid          ( clint_axi_req.aw_valid        ),
    .m_axi_awready          ( clint_axi_resp.aw_ready       ),
    
    .m_axi_wdata            ( clint_axi_req.w.data          ),
    .m_axi_wstrb            ( clint_axi_req.w.strb          ),
    .m_axi_wvalid           ( clint_axi_req.w_valid         ),
    .m_axi_wready           ( clint_axi_resp.w_ready        ),
    
    .m_axi_araddr           ( clint_axi_req.ar.addr         ),
    .m_axi_arvalid          ( clint_axi_req.ar_valid        ),
    .m_axi_arready          ( clint_axi_resp.ar_ready       ),
    
    .m_axi_rdata            ( clint_axi_resp.r.data         ),
    .m_axi_rresp            ( clint_axi_resp.r.resp         ),
    .m_axi_rvalid           ( clint_axi_resp.r_valid        ),
    .m_axi_rready           ( clint_axi_req.r_ready         ),
    
    .m_axi_bresp            ( clint_axi_resp.b.resp         ),
    .m_axi_bvalid           ( clint_axi_resp.b_valid        ),
    .m_axi_bready           ( clint_axi_req.b_ready         ),
    
    .w_reqbuf_size          (                               ),
    .r_reqbuf_size          (                               )
  );
  
  assign clint_axi_req.aw.id     = '0;
  assign clint_axi_req.aw.len    = '0;
  assign clint_axi_req.aw.size   = 3'b11;
  assign clint_axi_req.aw.burst  = '0;
  assign clint_axi_req.aw.lock   = '0;
  assign clint_axi_req.aw.cache  = '0;
  assign clint_axi_req.aw.prot   = '0;
  assign clint_axi_req.aw.qos    = '0;
  assign clint_axi_req.aw.region = '0;
  assign clint_axi_req.aw.atop   = '0;
  assign clint_axi_req.w.last    = 1'b1;
  assign clint_axi_req.ar.id     = '0;
  assign clint_axi_req.ar.len    = '0;
  assign clint_axi_req.ar.size   = 3'b11;
  assign clint_axi_req.ar.burst  = '0;
  assign clint_axi_req.ar.lock   = '0;
  assign clint_axi_req.ar.cache  = '0;
  assign clint_axi_req.ar.prot   = '0;
  assign clint_axi_req.ar.qos    = '0;
  assign clint_axi_req.ar.region = '0;
  
  
  
  AXI_BUS #(
    .AXI_ID_WIDTH   ( AxiIdWidth   ),
    .AXI_ADDR_WIDTH ( AxiAddrWidth ),
    .AXI_DATA_WIDTH ( AxiDataWidth ),
    .AXI_USER_WIDTH ( AxiUserWidth )
  ) plic_master();
  noc_axilite_bridge #(
    
    
    
    .SLAVE_RESP_BYTEWIDTH   ( 0             ),
    .SWAP_ENDIANESS         ( SwapEndianess ),
    
    .ALIGN_RDATA            ( 0             )
  ) i_plic_axilite_bridge (
    .clk                    ( clk_i                        ),
    .rst                    ( ~rst_ni                      ),
    
    .splitter_bridge_val    ( buf_ariane_plic_noc2_valid_i ),
    .splitter_bridge_data   ( buf_ariane_plic_noc2_data_i  ),
    .bridge_splitter_rdy    ( ariane_plic_buf_noc2_ready_o ),
    .bridge_splitter_val    ( ariane_plic_buf_noc3_valid_o ),
    .bridge_splitter_data   ( ariane_plic_buf_noc3_data_o  ),
    .splitter_bridge_rdy    ( buf_ariane_plic_noc3_ready_i ),
    
    
    .m_axi_awaddr           ( plic_master.aw_addr               ),
    .m_axi_awvalid          ( plic_master.aw_valid              ),
    .m_axi_awready          ( plic_master.aw_ready              ),
    
    .m_axi_wdata            ( plic_master.w_data                ),
    .m_axi_wstrb            ( plic_master.w_strb                ),
    .m_axi_wvalid           ( plic_master.w_valid               ),
    .m_axi_wready           ( plic_master.w_ready               ),
    
    .m_axi_araddr           ( plic_master.ar_addr               ),
    .m_axi_arvalid          ( plic_master.ar_valid              ),
    .m_axi_arready          ( plic_master.ar_ready              ),
    
    .m_axi_rdata            ( plic_master.r_data                ),
    .m_axi_rresp            ( plic_master.r_resp                ),
    .m_axi_rvalid           ( plic_master.r_valid               ),
    .m_axi_rready           ( plic_master.r_ready               ),
    
    .m_axi_bresp            ( plic_master.b_resp                ),
    .m_axi_bvalid           ( plic_master.b_valid               ),
    .m_axi_bready           ( plic_master.b_ready               ),
    
    .w_reqbuf_size          ( plic_master.aw_size               ),
    .r_reqbuf_size          ( plic_master.ar_size               )
  );
  
  assign plic_master.aw_id     = '0;
  assign plic_master.aw_len    = '0;
  assign plic_master.aw_burst  = '0;
  assign plic_master.aw_lock   = '0;
  assign plic_master.aw_cache  = '0;
  assign plic_master.aw_prot   = '0;
  assign plic_master.aw_qos    = '0;
  assign plic_master.aw_region = '0;
  assign plic_master.aw_atop   = '0;
  assign plic_master.w_last    = 1'b1;
  assign plic_master.ar_id     = '0;
  assign plic_master.ar_len    = '0;
  assign plic_master.ar_burst  = '0;
  assign plic_master.ar_lock   = '0;
  assign plic_master.ar_cache  = '0;
  assign plic_master.ar_prot   = '0;
  assign plic_master.ar_qos    = '0;
  assign plic_master.ar_region = '0;
  reg_intf::reg_intf_resp_d32 plic_resp;
  reg_intf::reg_intf_req_a32_d32 plic_req;
  enum logic [2:0] {Idle, WriteSecond, ReadSecond, WriteResp, ReadResp} state_d, state_q;
  logic [31:0] rword_d, rword_q;
  
  assign rword_d = (plic_req.valid && !plic_req.write) ? plic_resp.rdata : rword_q;
  assign plic_master.r_data = {plic_resp.rdata, rword_q};
  always_ff @(posedge clk_i or negedge rst_ni) begin : p_plic_regs
    if (!rst_ni) begin
      state_q <= Idle;
      rword_q <= '0;
    end else begin
      state_q <= state_d;
      rword_q <= rword_d;
    end
  end
  
  
  always_comb begin : p_plic_if
    automatic logic [31:0] waddr, raddr;
    
    waddr = plic_master.aw_addr[31:0] - 32'(PlicBase) + 32'hc000000;
    raddr = plic_master.ar_addr[31:0] - 32'(PlicBase) + 32'hc000000;
    
    plic_master.aw_ready = plic_resp.ready;
    plic_master.w_ready  = plic_resp.ready;
    plic_master.ar_ready = plic_resp.ready;
    plic_master.r_valid  = 1'b0;
    plic_master.r_resp   = '0;
    plic_master.b_valid  = 1'b0;
    plic_master.b_resp   = '0;
    
    plic_req.valid       = 1'b0;
    plic_req.wstrb       = '0;
    plic_req.write       = 1'b0;
    plic_req.wdata       = plic_master.w_data[31:0];
    plic_req.addr        = waddr;
    
    state_d              = state_q;
    unique case (state_q)
      Idle: begin
        if (plic_master.w_valid && plic_master.aw_valid && plic_resp.ready) begin
          plic_req.valid = 1'b1;
          plic_req.write = plic_master.w_strb[3:0];
          plic_req.wstrb = '1;
          
          if (plic_master.aw_size == 3'b11) begin
            state_d = WriteSecond;
          end else begin
            state_d = WriteResp;
          end
        end else if (plic_master.ar_valid && plic_resp.ready) begin
          plic_req.valid = 1'b1;
          plic_req.addr  = raddr;
          
          if (plic_master.ar_size == 3'b11) begin
            state_d = ReadSecond;
          end else begin
            state_d = ReadResp;
          end
        end
      end
      
      WriteSecond: begin
        plic_master.aw_ready = 1'b0;
        plic_master.w_ready  = 1'b0;
        plic_master.ar_ready = 1'b0;
        plic_req.addr        = waddr + 32'h4;
        plic_req.wdata       = plic_master.w_data[63:32];
        if (plic_resp.ready && plic_master.b_ready) begin
          plic_req.valid       = 1'b1;
          plic_req.write       = 1'b1;
          plic_req.wstrb       = '1;
          plic_master.b_valid  = 1'b1;
          state_d              = Idle;
        end
      end
      
      ReadSecond: begin
        plic_master.aw_ready = 1'b0;
        plic_master.w_ready  = 1'b0;
        plic_master.ar_ready = 1'b0;
        plic_req.addr        = raddr + 32'h4;
        if (plic_resp.ready && plic_master.r_ready) begin
          plic_req.valid      = 1'b1;
          plic_master.r_valid = 1'b1;
          state_d             = Idle;
        end
      end
      WriteResp: begin
        plic_master.aw_ready = 1'b0;
        plic_master.w_ready  = 1'b0;
        plic_master.ar_ready = 1'b0;
        if (plic_master.b_ready) begin
          plic_master.b_valid  = 1'b1;
          state_d              = Idle;
        end
      end
      ReadResp: begin
        plic_master.aw_ready = 1'b0;
        plic_master.w_ready  = 1'b0;
        plic_master.ar_ready = 1'b0;
        if (plic_master.r_ready) begin
          plic_master.r_valid = 1'b1;
          state_d             = Idle;
        end
      end
      default: state_d = Idle;
    endcase
  end
  plic_top #(
    .N_SOURCE    ( NumSources      ),
    .N_TARGET    ( 2*NumHarts      ),
    .MAX_PRIO    ( PlicMaxPriority )
  ) i_plic (
    .clk_i,
    .rst_ni,
    .req_i         ( plic_req    ),
    .resp_o        ( plic_resp   ),
    .le_i          ( irq_le_i    ), 
    .irq_sources_i,                 
    .eip_targets_o ( irq_o       )
  );
endmodule 
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 215;
    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00766564,
        64'h6e2c7663_73697200,
        64'h79746972_6f697270,
        64'h2d78616d_2c766373,
        64'h69720073_656d616e,
        64'h2d676572_00646564,
        64'h6e657478_652d7374,
        64'h70757272_65746e69,
        64'h00746669_68732d67,
        64'h65720073_74707572,
        64'h7265746e_6900746e,
        64'h65726170_2d747075,
        64'h72726574_6e690064,
        64'h65657073_2d746e65,
        64'h72727563_00736567,
        64'h6e617200_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h006c6564_6f6d0065,
        64'h6c626974_61706d6f,
        64'h6300736c_6c65632d,
        64'h657a6973_2300736c,
        64'h6c65632d_73736572,
        64'h64646123_09000000,
        64'h02000000_02000000,
        64'h02000000_01000000,
        64'ha9000000_04000000,
        64'h03000000_01000000,
        64'h1d010000_04000000,
        64'h03000000_07000000,
        64'h0a010000_04000000,
        64'h03000000_00000004,
        64'h00000000_000010f1,
        64'hff000000_5b000000,
        64'h10000000_03000000,
        64'h09000000_02000000,
        64'h0b000000_02000000,
        64'hec000000_10000000,
        64'h03000000_94000000,
        64'h00000000_03000000,
        64'h00306369_6c702c76,
        64'h63736972_1b000000,
        64'h0c000000_03000000,
        64'h01000000_83000000,
        64'h04000000_03000000,
        64'h00000000_00000000,
        64'h04000000_03000000,
        64'h00303030_30303131,
        64'h66666640_63696c70,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'h00010000_08000000,
        64'h03000000_00000c00,
        64'h00000000_000002f1,
        64'hff000000_5b000000,
        64'h10000000_03000000,
        64'h07000000_02000000,
        64'h03000000_02000000,
        64'hec000000_10000000,
        64'h03000000_00000000,
        64'h30746e69_6c632c76,
        64'h63736972_1b000000,
        64'h0d000000_03000000,
        64'h00000000_30303030,
        64'h32303166_66664074,
        64'h6e696c63_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_00010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h000000f1_ff000000,
        64'h5b000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_ec000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00303030,
        64'h30303031_66666640,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h00000000_e2000000,
        64'h04000000_03000000,
        64'h01000000_d7000000,
        64'h04000000_03000000,
        64'h01000000_c6000000,
        64'h04000000_03000000,
        64'h00c20100_b8000000,
        64'h04000000_03000000,
        64'h80f0fa02_3f000000,
        64'h04000000_03000000,
        64'h00400d00_00000000,
        64'h00c0c2f0_ff000000,
        64'h5b000000_10000000,
        64'h03000000_00303535,
        64'h3631736e_1b000000,
        64'h08000000_03000000,
        64'h00303030_63326330,
        64'h66666640_74726175,
        64'h01000000_b1000000,
        64'h00000000_03000000,
        64'h00007375_622d656c,
        64'h706d6973_00636f73,
        64'h2d657261_622d656e,
        64'h61697261_2c687465,
        64'h1b000000_1f000000,
        64'h03000000_02000000,
        64'h0f000000_04000000,
        64'h03000000_02000000,
        64'h00000000_04000000,
        64'h03000000_00636f73,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h5b000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_4f000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_a9000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_94000000,
        64'h00000000_03000000,
        64'h01000000_83000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_79000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_70000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_66000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h5f000000_05000000,
        64'h03000000_00000000,
        64'h5b000000_04000000,
        64'h03000000_00757063,
        64'h4f000000_04000000,
        64'h03000000_80f0fa02,
        64'h3f000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'he1f50500_2c000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hd4040000_28010000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h0c050000_38000000,
        64'h34060000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_0000bff5,
        64'h10500073_03c58593,
        64'h00000597_f1402573,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_84020765,
        64'h85930000_0597f140,
        64'h2573047e_0010041b
    };
    logic [$clog2(RomSize)-1:0] addr_q;
    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end
    
    
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
module bootrom_linux (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 732;
    const logic [RomSize-1:0][63:0] mem = {
        64'h000000ff_f0c2c004,
        64'h000000ff_f0c2c003,
        64'h000000ff_f0c2c001,
        64'h000000ff_f0c2c005,
        64'h00000000_00000000,
        64'h0a0d2165_6e6f6420,
        64'h00000000_00206567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f63,
        64'h00000000_00000009,
        64'h3a656d61_6e090a0d,
        64'h00093a73_65747562,
        64'h69727474_61090a0d,
        64'h00000009_3a61626c,
        64'h20747361_6c090a0d,
        64'h0000093a_61626c20,
        64'h74737269_66090a0d,
        64'h00000000_00000000,
        64'h09202020_20203a64,
        64'h69756720_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_00000000,
        64'h093a6469_75672065,
        64'h70797420_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20747067,
        64'h00000009_20203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20657a69_73090a0d,
        64'h00000009_3a736569,
        64'h72746e65_206e6f69,
        64'h74697472_61702072,
        64'h65626d75_6e090a0d,
        64'h00000009_2020203a,
        64'h61626c20_73656972,
        64'h746e6520_6e6f6974,
        64'h69747261_70090a0d,
        64'h00093a61_646c2070,
        64'h756b6361_62090a0d,
        64'h00000000_00000000,
        64'h093a6162_6c20746e,
        64'h65727275_63090a0d,
        64'h00000009_3a646576,
        64'h72657365_72090a0d,
        64'h00093a72_65646165,
        64'h685f6372_63090a0d,
        64'h00000000_00000909,
        64'h3a657a69_73090a0d,
        64'h00000009_3a6e6f69,
        64'h73697665_72090a0d,
        64'h0000093a_65727574,
        64'h616e6769_73090a0d,
        64'h00000000_003a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20747067,
        64'h0000203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_63206473,
        64'h00000000_0000000a,
        64'h0d216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_0a0d676e,
        64'h69746978_65202e2e,
        64'h2e647320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f63,
        64'h00000000_00292520,
        64'h00000000_00000028,
        64'h20736b63_6f6c6220,
        64'h00000000_20666f20,
        64'h0000206b_636f6c62,
        64'h20676e69_79706f63,
        64'h00000000_00000008,
        64'h0000000a_0d202e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e69,
        64'h00000000_203f3f79,
        64'h74706d65_20746f6e,
        64'h206f6669_66207872,
        64'h00000000_00000a0d,
        64'h2164657a_696c6169,
        64'h74696e69_20495053,
        64'h00000000_00007830,
        64'h203a7375_74617473,
        64'h00000000_00000a0d,
        64'h49505320_74696e69,
        64'h00000000_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_00766564,
        64'h6e2c7663_73697200,
        64'h79746972_6f697270,
        64'h2d78616d_2c766373,
        64'h69720073_656d616e,
        64'h2d676572_00646564,
        64'h6e657478_652d7374,
        64'h70757272_65746e69,
        64'h00746669_68732d67,
        64'h65720073_74707572,
        64'h7265746e_6900746e,
        64'h65726170_2d747075,
        64'h72726574_6e690064,
        64'h65657073_2d746e65,
        64'h72727563_00736567,
        64'h6e617200_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h006c6564_6f6d0065,
        64'h6c626974_61706d6f,
        64'h6300736c_6c65632d,
        64'h657a6973_2300736c,
        64'h6c65632d_73736572,
        64'h64646123_09000000,
        64'h02000000_02000000,
        64'h02000000_01000000,
        64'ha9000000_04000000,
        64'h03000000_01000000,
        64'h1d010000_04000000,
        64'h03000000_07000000,
        64'h0a010000_04000000,
        64'h03000000_00000004,
        64'h00000000_000010f1,
        64'hff000000_5b000000,
        64'h10000000_03000000,
        64'h09000000_02000000,
        64'h0b000000_02000000,
        64'hec000000_10000000,
        64'h03000000_94000000,
        64'h00000000_03000000,
        64'h00306369_6c702c76,
        64'h63736972_1b000000,
        64'h0c000000_03000000,
        64'h01000000_83000000,
        64'h04000000_03000000,
        64'h00000000_00000000,
        64'h04000000_03000000,
        64'h00303030_30303131,
        64'h66666640_63696c70,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'h00010000_08000000,
        64'h03000000_00000c00,
        64'h00000000_000002f1,
        64'hff000000_5b000000,
        64'h10000000_03000000,
        64'h07000000_02000000,
        64'h03000000_02000000,
        64'hec000000_10000000,
        64'h03000000_00000000,
        64'h30746e69_6c632c76,
        64'h63736972_1b000000,
        64'h0d000000_03000000,
        64'h00000000_30303030,
        64'h32303166_66664074,
        64'h6e696c63_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_00010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h000000f1_ff000000,
        64'h5b000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_ec000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00303030,
        64'h30303031_66666640,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h00000000_e2000000,
        64'h04000000_03000000,
        64'h01000000_d7000000,
        64'h04000000_03000000,
        64'h01000000_c6000000,
        64'h04000000_03000000,
        64'h00c20100_b8000000,
        64'h04000000_03000000,
        64'h80f0fa02_3f000000,
        64'h04000000_03000000,
        64'h00400d00_00000000,
        64'h00c0c2f0_ff000000,
        64'h5b000000_10000000,
        64'h03000000_00303535,
        64'h3631736e_1b000000,
        64'h08000000_03000000,
        64'h00303030_63326330,
        64'h66666640_74726175,
        64'h01000000_b1000000,
        64'h00000000_03000000,
        64'h00007375_622d656c,
        64'h706d6973_00636f73,
        64'h2d657261_622d656e,
        64'h61697261_2c687465,
        64'h1b000000_1f000000,
        64'h03000000_02000000,
        64'h0f000000_04000000,
        64'h03000000_02000000,
        64'h00000000_04000000,
        64'h03000000_00636f73,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h5b000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_4f000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_a9000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_94000000,
        64'h00000000_03000000,
        64'h01000000_83000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_79000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_70000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_66000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h5f000000_05000000,
        64'h03000000_00000000,
        64'h5b000000_04000000,
        64'h03000000_00757063,
        64'h4f000000_04000000,
        64'h03000000_80f0fa02,
        64'h3f000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'he1f50500_2c000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hd4040000_28010000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h0c050000_38000000,
        64'h34060000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000a0d,
        64'h0a0d0a0d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_0a0d2020,
        64'h20202020_20202020,
        64'h34202f20_426b2034,
        64'h36202020_3a636f73,
        64'h7341202f_20657a69,
        64'h53202032_4c0a0d20,
        64'h20202020_20202020,
        64'h2034202f_20426b20,
        64'h38202020_203a636f,
        64'h73734120_2f20657a,
        64'h69532035_314c0a0d,
        64'h20202020_20202020,
        64'h20203420_2f20426b,
        64'h20382020_20203a63,
        64'h6f737341_202f2065,
        64'h7a695320_44314c0a,
        64'h0d202020_20202020,
        64'h20202034_202f2042,
        64'h6b203631_2020203a,
        64'h636f7373_41202f20,
        64'h657a6953_2049314c,
        64'h0a0d2020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20200a0d_20202020,
        64'h20202020_20202020,
        64'h20202020_424d2034,
        64'h32303120_20202020,
        64'h20202020_3a657a69,
        64'h53204d41_52440a0d,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202068_73656d5f,
        64'h64322020_20202020,
        64'h20202020_203a6b72,
        64'h6f777465_4e0a0d20,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20206e77_6f6e6b6e,
        64'h55202020_20202020,
        64'h20203a71_65724620,
        64'h65726f43_0a0d2020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20312020_20202020,
        64'h20202020_20203a73,
        64'h65726f43_230a0d20,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20203120_20202020,
        64'h20202020_203a7365,
        64'h6c69542d_59230a0d,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202031_20202020,
        64'h20202020_20203a73,
        64'h656c6954_2d58230a,
        64'h0d202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h200a0d20_20202020,
        64'h20202020_20202020,
        64'h20202020_20203833,
        64'h3a35333a_32302031,
        64'h32303220_39312067,
        64'h75412020_20202020,
        64'h20203a65_74614420,
        64'h646c6975_420a0d20,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h2020296e_6f697461,
        64'h6c756d69_53282065,
        64'h6e6f4e20_20202020,
        64'h2020203a_6472616f,
        64'h42204147_50460a0d,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h0a0d2020_20202020,
        64'h20202020_20202020,
        64'h20202020_20273635,
        64'h33666362_62632762,
        64'h20202020_3a6e6f69,
        64'h73726556_20656e61,
        64'h6972410a_0d202020,
        64'h20202020_20202020,
        64'h20202020_20202020,
        64'h27636266_35663666,
        64'h65276220_3a6e6f69,
        64'h73726556_206e6f74,
        64'h69506e65_704f0a0d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h0a0d2d2d_20202020,
        64'h20206d72_6f667461,
        64'h6c502065_6e616972,
        64'h412b6e6f_7469506e,
        64'h65704f20_20202020,
        64'h2d2d0a0d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_2d2d2d2d,
        64'h2d2d2d2d_0a0d0a0d,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_80820141,
        64'h450160a2_cfdff0ef,
        64'h057e65a1_45058e3f,
        64'hf0efb425_05130000,
        64'h15178eff_f0ef1565,
        64'h05130000_05178a1f,
        64'hf0efe406_38050513,
        64'h20058593_114101c9,
        64'hc53765f1_b395913f,
        64'hf0efe2a5_05130000,
        64'h1517bbd9_bc450513,
        64'h00001517_a35ff0ef,
        64'h854a92ff_f0efc865,
        64'h05130000_151793bf,
        64'hf0efc7a5_05130000,
        64'h1517bbfd_bec50513,
        64'h00001517_a5dff0ef,
        64'h8526957f_f0efcae5,
        64'h05130000_1517963f,
        64'hf0efca25_05130000,
        64'h1517c929_84aac97f,
        64'hf0ef8552_8656020b,
        64'h258397ff_f0efc265,
        64'h05130000_151798bf,
        64'hf0efe8a5_05130000,
        64'h1517f579_10e30804,
        64'h849399ff_f0ef2905,
        64'hc4850513_00001517,
        64'hff999be3_b01ff0ef,
        64'h09850009_c5039bbf,
        64'hf0efeaa5_05130000,
        64'h1517ad3f_f0ef6888,
        64'h9cdff0ef_eac50513,
        64'h00001517_ae5ff0ef,
        64'h64889dff_f0efeae5,
        64'h05130000_1517af7f,
        64'hf0ef0604_8c930184,
        64'h89936088_9f9ff0ef,
        64'heb850513_00001517,
        64'hfe999be3_b59ff0ef,
        64'h09850009_c503ff04,
        64'h8993a17f_f0efeb65,
        64'h05130000_1517ff89,
        64'h99e3b77f_f0ef0985,
        64'h0007c503_013c87b3,
        64'h4981a37f_f0effe04,
        64'h8c93eba5_05130000,
        64'h1517b97f_f0ef0ff9,
        64'h7513a4ff_f0efeb65,
        64'h05130000_15174b91,
        64'h4c411005_1e631004,
        64'h892a8b0a_d8dff0ef,
        64'h850a4605_71010489,
        64'h2583a77f_f0efd1e5,
        64'h05130000_1517b4df,
        64'hf0ef4556_a89ff0ef,
        64'hed050513_00001517,
        64'hb5fff0ef_4546a9bf,
        64'hf0efec25_05130000,
        64'h1517bb3f_f0ef6526,
        64'haadff0ef_eb450513,
        64'h00001517_bc5ff0ef,
        64'h7502abff_f0efeb65,
        64'h05130000_1517bd7f,
        64'hf0ef6562_ad1ff0ef,
        64'heb050513_00001517,
        64'hba7ff0ef_4552ae3f,
        64'hf0efeb25_05130000,
        64'h1517bb9f_f0ef4542,
        64'haf5ff0ef_eb450513,
        64'h00001517_bcbff0ef,
        64'h4532b07f_f0efeb65,
        64'h05130000_1517bddf,
        64'hf0ef4522_b19ff0ef,
        64'heb850513_00001517,
        64'hc31ff0ef_6502b2bf,
        64'hf0efeba5_05130000,
        64'h1517b37f_f0efea65,
        64'h05130000_1517bf59,
        64'h54f9b47f_f0efdee5,
        64'h05130000_1517c5ff,
        64'hf0ef8526_b59ff0ef,
        64'heb050513_00001517,
        64'hb65ff0ef_ea450513,
        64'h00001517_c90584aa,
        64'h890ae9bf_f0ef850a,
        64'h45854605_7101b83f,
        64'hf0efde25_05130000,
        64'h15178082_61256ca2,
        64'h6c426be2_7b027aa2,
        64'h7a4279e2_690664a6,
        64'h64468526_60e6fa04,
        64'h011354fd_bb1ff0ef,
        64'hec850513_00001517,
        64'hc905ecbf_f0ef8aae,
        64'h8a2a1080_e466e862,
        64'hec5ef05a_fc4ee0ca,
        64'he4a6ec86_f456f852,
        64'he8a2711d_b7bd2c05,
        64'hbe5ff0ef_ec450513,
        64'h00001517_b7a10b85,
        64'h20048493_ff5799e3,
        64'he29007a1_00e786b3,
        64'h621000f4_86334781,
        64'h974e009b_97139c29,
        64'hc15ff0ef_f2450513,
        64'h00001517_9c29c75f,
        64'hf0ef0325_553b4585,
        64'h036a053b_9c29c33f,
        64'hf0eff325_05130000,
        64'h15179c29_c93ff0ef,
        64'h854a9c29_4585c4bf,
        64'hf0eff425_05130000,
        64'h15179c29_cabff0ef,
        64'h855a0005_041b4585,
        64'hc65ff0ef_f4c50513,
        64'h00001517_09841263,
        64'h060c1363_034b7c3b,
        64'h80826161_45016c02,
        64'h6ba26b42_6ae27a02,
        64'h79a27942_74e26406,
        64'h60a6c97f_f0eff3e5,
        64'h05130000_1517032b,
        64'h6563000b_8b1b2000,
        64'h0a930640_0a134401,
        64'h4b8100f5_84b38932,
        64'h89aae062_e85ae486,
        64'he45eec56_f052f44e,
        64'hf84afc26_e0a21792,
        64'h715d47bd_0177d593,
        64'h02059793_80820141,
        64'h450160a2_ce9ff0ef,
        64'he406fb45_05131141,
        64'h00001517_8082557d,
        64'hb7d900d7_00230785,
        64'h00f60733_06c82683,
        64'hff698b05_5178b77d,
        64'hd6b80785_00074703,
        64'h00f50733_80824501,
        64'hd3b84719_dbb8577d,
        64'h200007b7_02b6e163,
        64'h0007869b_20000837,
        64'h20000537_fff58b85,
        64'h537c2000_0737d3b8,
        64'h200007b7_10600713,
        64'hfff537fd_00010320,
        64'h079304b7_61630007,
        64'h871b4781_200006b7,
        64'hdbb85779_200007b7,
        64'h06b7ee63_10000793,
        64'h80826105_64a2d3b8,
        64'h4719dbb8_64420ff4,
        64'h7513577d_200007b7,
        64'h60e2d97f_f0ef03e5,
        64'h05130000_1517eaff,
        64'hf0ef9101_15024088,
        64'hdadff0ef_05c50513,
        64'h00001517_e3958b85,
        64'h240153fc_57e0ff65,
        64'h8b050647_849353f8,
        64'hd3b81060_07132000,
        64'h07b7fff5_37fd0001,
        64'h06400793_d7a8dbb8,
        64'h5779e426_e822ec06,
        64'h200007b7_1101bbc5,
        64'h610508a5_05130000,
        64'h151764a2_60e26442,
        64'hd03c4799_e09ff0ef,
        64'h0b050513_00001517,
        64'hf21ff0ef_91010204,
        64'h95132481_e21ff0ef,
        64'h0a850513_00001517,
        64'h5064d03c_16600793,
        64'he35ff0ef_0dc50513,
        64'h00001517_f4dff0ef,
        64'h91010204_95132481,
        64'he4dff0ef_0d450513,
        64'h00001517_5064d03c,
        64'h10400793_20000437,
        64'hfff537fd_000147a9,
        64'hc3b84729_200007b7,
        64'he75ff0ef_e426e822,
        64'hec060f45_05131101,
        64'h00001517_80822501,
        64'h41088082_c10c8082,
        64'h61054509_60e2e1ff,
        64'hf0ef0091_4503e27f,
        64'hf0ef0081_4503ed9f,
        64'hf0efec06_002c1101,
        64'h80826145_45416942,
        64'h64e27402_70a2ff24,
        64'h10e3e4bf_f0ef0091,
        64'h4503e53f_f0ef3461,
        64'h00814503_f07ff0ef,
        64'h0ff57513_002c0084,
        64'hd5335961_03800413,
        64'h84aaf406_e84aec26,
        64'hf0227179_80826145,
        64'h45216942_64e27402,
        64'h70a2ff24_10e3e8ff,
        64'hf0ef0091_4503e97f,
        64'hf0ef3461_00814503,
        64'hf4bff0ef_0ff57513,
        64'h002c0084_d53b5961,
        64'h446184aa_f406e84a,
        64'hec26f022_71798082,
        64'h612169e2_854e6b02,
        64'h6aa26a42_790274a2,
        64'h744270e2_fd5913e3,
        64'h397d85d2_eddff0ef,
        64'h0007c503_97ba8bbd,
        64'h02d7d7bb_29856ce7,
        64'h07130000_071702ba,
        64'h706300d7_f4630364,
        64'h543b0009_0a1b0284,
        64'hf4bb0004_069b0004,
        64'h879b5afd_4b294981,
        64'h4925a004_041384aa,
        64'he852fc06_e05ae456,
        64'hec4ef04a_f4263b9a,
        64'hd437f822_71398082,
        64'h00f58023_0007c783,
        64'h00e580a3_97aa8111,
        64'h00074703_973e00f5,
        64'h77137327_87930000,
        64'h0797b7c5_f5dff0ef,
        64'h853e8082_610564a2,
        64'h644260e2_e791fff7,
        64'hc7830084_87b30405,
        64'h0004051b_440184aa,
        64'hec06e426_e8221101,
        64'h808200e7_80230200,
        64'h071354a7_b7830000,
        64'h179700f7_0023478d,
        64'h00a68023_0ff57513,
        64'h00c78023_0085551b,
        64'h0ff57613_07ba30b7,
        64'h879303ff_c7b700f7,
        64'h0023f800_07930006,
        64'h802357a7_b7030000,
        64'h179757a7_b6830000,
        64'h179702b5_553b0045,
        64'h959b8082_00a78023,
        64'h07ba30b7_879303ff,
        64'hc7b7dbe5_0207f793,
        64'h0007c783_59c7b783,
        64'h00001797_80820205,
        64'h75130007_c5035ae7,
        64'hb7830000_17978082,
        64'h0ff57513_00054503,
        64'h808200b5_00238082,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00048067,
        64'h01f49493_0010049b,
        64'hd6058593_00001597,
        64'hf1402573_ff2496e3,
        64'h00100493_0004a903,
        64'h04048493_01a49493,
        64'h0210049b_0924a4af,
        64'h00190913_04048493,
        64'h01a49493_0210049b,
        64'hff2496e3_f14024f3,
        64'h0004a903_04048493,
        64'h01a49493_0210049b,
        64'h081000ef_01a11113,
        64'h0210011b_01249863,
        64'hf1402973_00000493
    };
    logic [$clog2(RomSize)-1:0] addr_q;
    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end
    
    
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
module rv_plic_target #(
  parameter int N_SOURCE = 32,
  parameter int MAX_PRIO = 7,
  parameter     ALGORITHM = "SEQUENTIAL", 
  
  parameter int unsigned SRCW  = $clog2(N_SOURCE+1),
  parameter int unsigned PRIOW = $clog2(MAX_PRIO+1) 
) (
  input clk_i,
  input rst_ni,
  input [N_SOURCE-1:0] ip,
  input [N_SOURCE-1:0] ie,
  input [N_SOURCE-1:0][PRIOW-1:0] prio,
  input [PRIOW-1:0] threshold,
  output logic            irq,
  output logic [SRCW-1:0] irq_id
);
if (ALGORITHM == "SEQUENTIAL") begin : gen_sequential
  
  
  
  logic [PRIOW-1:0] max_prio;
  logic irq_next;
  logic [SRCW-1:0] irq_id_next;
  always_comb begin
    max_prio = threshold + 1'b1; 
    irq_id_next = '0; 
    irq_next = 1'b0;
    for (int i = N_SOURCE-1 ; i >= 0 ; i--) begin
      if ((ip[i] & ie[i]) == 1'b1 && prio[i] >= max_prio) begin
        max_prio = prio[i];
        irq_id_next = SRCW'(i+1);
        irq_next = 1'b1;
      end
    end 
  end
  always_ff @(posedge clk_i, negedge rst_ni) begin
    if (!rst_ni) begin
      irq <= 1'b0;
      irq_id <= '0;
    end else begin
      irq <= irq_next;
      irq_id <= irq_id_next;
    end
  end
end else if (ALGORITHM == "MATRIX") begin : gen_mat
  
  
  
  
  
  
  
  logic [N_SOURCE-1:0] is;
  logic [N_SOURCE-1:0][N_SOURCE-1:0] mat;
  logic [N_SOURCE-1:0] merged_row;
  assign is = ip & ie;
  always_comb begin
    merged_row[N_SOURCE-1] = is[N_SOURCE-1] & (prio[N_SOURCE-1] > threshold);
    for (int i = 0 ; i < N_SOURCE-1 ; i++) begin
      merged_row[i] = 1'b1;
      for (int j = i+1 ; j < N_SOURCE ; j++) begin
        mat[i][j] = (prio[i] <= threshold) ? 1'b0 :         
                    (is[i] & is[j]) ? prio[i] >= prio[j] :
                    (is[i]) ? 1'b 1 : 1'b 0 ;
        merged_row[i] = merged_row[i] & mat[i][j]; 
      end 
    end 
  end 
  
  logic [N_SOURCE-1:0] lod;
  assign lod = merged_row & (~merged_row + 1'b1);
  always_ff @(posedge clk_i, negedge rst_ni) begin
    if (!rst_ni) begin
      irq <= 1'b0;
      irq_id <= '0; 
    end else if (|lod) begin
      
      
      for (int i = N_SOURCE-1 ; i >= 0 ; i--) begin
        if (lod[i] == 1'b1) begin
          irq <= 1'b 1;
          irq_id <= SRCW'(i + 1);
        end
      end 
    end else begin
      
      irq <= 1'b0;
      irq_id <= '0;
    end
  end 
end 
endmodule
module rv_plic_gateway #(
  parameter int N_SOURCE = 32
) (
  input clk_i,
  input rst_ni,
  input [N_SOURCE-1:0] src,
  input [N_SOURCE-1:0] le,      
  input [N_SOURCE-1:0] claim, 
  input [N_SOURCE-1:0] complete, 
  output logic [N_SOURCE-1:0] ip
);
logic [N_SOURCE-1:0] ia;    
logic [N_SOURCE-1:0] set;   
logic [N_SOURCE-1:0] src_d;
always_ff @(posedge clk_i, negedge rst_ni) begin
  if (!rst_ni) src_d <= '0;
  else         src_d <= src;
end
always_comb begin
  for (int i = 0 ; i < N_SOURCE; i++) begin
    set[i] = (le[i]) ? src[i] & ~src_d[i] : src[i] ;
  end
end
always_ff @(posedge clk_i, negedge rst_ni) begin
  if (!rst_ni) begin
    ip <= '0;
  end else begin
    ip <= (ip | (set & ~ia & ~ip)) & (~claim);
  end
end
always_ff @(posedge clk_i, negedge rst_ni) begin
  if (!rst_ni) begin
    ia <= '0;
  end else begin
    ia <= (ia | (set & ~ia)) & (~complete);
  end
end
endmodule
module plic_regs (
  input logic [2:0][2:0] prio_i,
  output logic [2:0][2:0] prio_o,
  output logic [2:0] prio_we_o,
  output logic [2:0] prio_re_o,
  input logic [0:0][2:0] ip_i,
  output logic [0:0] ip_re_o,
  input logic [1:0][2:0] ie_i,
  output logic [1:0][2:0] ie_o,
  output logic [1:0] ie_we_o,
  output logic [1:0] ie_re_o,
  input logic [1:0][2:0] threshold_i,
  output logic [1:0][2:0] threshold_o,
  output logic [1:0] threshold_we_o,
  output logic [1:0] threshold_re_o,
  input logic [1:0][1:0] cc_i,
  output logic [1:0][1:0] cc_o,
  output logic [1:0] cc_we_o,
  output logic [1:0] cc_re_o,
  
  input  reg_intf::reg_intf_req_a32_d32 req_i,
  output reg_intf::reg_intf_resp_d32    resp_o
);
always_comb begin
  resp_o.ready = 1'b1;
  resp_o.rdata = '0;
  resp_o.error = '0;
  prio_o = '0;
  prio_we_o = '0;
  prio_re_o = '0;
  ie_o = '0;
  ie_we_o = '0;
  ie_re_o = '0;
  threshold_o = '0;
  threshold_we_o = '0;
  threshold_re_o = '0;
  cc_o = '0;
  cc_we_o = '0;
  cc_re_o = '0;
  if (req_i.valid) begin
    if (req_i.write) begin
      unique case(req_i.addr)
        32'hc000000: begin
          prio_o[0][2:0] = req_i.wdata[2:0];
          prio_we_o[0] = 1'b1;
        end
        32'hc000004: begin
          prio_o[1][2:0] = req_i.wdata[2:0];
          prio_we_o[1] = 1'b1;
        end
        32'hc000008: begin
          prio_o[2][2:0] = req_i.wdata[2:0];
          prio_we_o[2] = 1'b1;
        end
        32'hc002000: begin
          ie_o[0][2:0] = req_i.wdata[2:0];
          ie_we_o[0] = 1'b1;
        end
        32'hc002080: begin
          ie_o[1][2:0] = req_i.wdata[2:0];
          ie_we_o[1] = 1'b1;
        end
        32'hc200000: begin
          threshold_o[0][2:0] = req_i.wdata[2:0];
          threshold_we_o[0] = 1'b1;
        end
        32'hc201000: begin
          threshold_o[1][2:0] = req_i.wdata[2:0];
          threshold_we_o[1] = 1'b1;
        end
        32'hc200004: begin
          cc_o[0][1:0] = req_i.wdata[1:0];
          cc_we_o[0] = 1'b1;
        end
        32'hc201004: begin
          cc_o[1][1:0] = req_i.wdata[1:0];
          cc_we_o[1] = 1'b1;
        end
        default: resp_o.error = 1'b1;
      endcase
    end else begin
      unique case(req_i.addr)
        32'hc000000: begin
          resp_o.rdata[2:0] = prio_i[0][2:0];
          prio_re_o[0] = 1'b1;
        end
        32'hc000004: begin
          resp_o.rdata[2:0] = prio_i[1][2:0];
          prio_re_o[1] = 1'b1;
        end
        32'hc000008: begin
          resp_o.rdata[2:0] = prio_i[2][2:0];
          prio_re_o[2] = 1'b1;
        end
        32'hc001000: begin
          resp_o.rdata[2:0] = ip_i[0][2:0];
          ip_re_o[0] = 1'b1;
        end
        32'hc002000: begin
          resp_o.rdata[2:0] = ie_i[0][2:0];
          ie_re_o[0] = 1'b1;
        end
        32'hc002080: begin
          resp_o.rdata[2:0] = ie_i[1][2:0];
          ie_re_o[1] = 1'b1;
        end
        32'hc200000: begin
          resp_o.rdata[2:0] = threshold_i[0][2:0];
          threshold_re_o[0] = 1'b1;
        end
        32'hc201000: begin
          resp_o.rdata[2:0] = threshold_i[1][2:0];
          threshold_re_o[1] = 1'b1;
        end
        32'hc200004: begin
          resp_o.rdata[1:0] = cc_i[0][1:0];
          cc_re_o[0] = 1'b1;
        end
        32'hc201004: begin
          resp_o.rdata[1:0] = cc_i[1][1:0];
          cc_re_o[1] = 1'b1;
        end
        default: resp_o.error = 1'b1;
      endcase
    end
  end
end
endmodule
module plic_top #(
  parameter int N_SOURCE    = 30,
  parameter int N_TARGET    = 2,
  parameter int MAX_PRIO    = 7,
  parameter int SRCW        = $clog2(N_SOURCE+1)
) (
  input  logic clk_i,    
  input  logic rst_ni,  
  
  input  reg_intf::reg_intf_req_a32_d32 req_i,
  output reg_intf::reg_intf_resp_d32    resp_o,
  input logic [N_SOURCE-1:0] le_i, 
  
  input  logic [N_SOURCE-1:0] irq_sources_i,
  
  output logic [N_TARGET-1:0] eip_targets_o
);
  localparam PRIOW = $clog2(MAX_PRIO+1);
  logic [N_SOURCE-1:0] ip;
  logic [N_TARGET-1:0][PRIOW-1:0]    threshold_q;
  logic [N_TARGET-1:0]               claim_re; 
  logic [N_TARGET-1:0][SRCW-1:0]     claim_id;
  logic [N_SOURCE-1:0]               claim; 
  logic [N_TARGET-1:0]               complete_we; 
  logic [N_TARGET-1:0][SRCW-1:0]     complete_id;
  logic [N_SOURCE-1:0]               complete; 
  logic [N_SOURCE-1:0][PRIOW-1:0]    prio_q;
  logic [N_TARGET-1:0][N_SOURCE-1:0] ie_q;
  always_comb begin
    claim = '0;
    complete = '0;
    for (int i = 0 ; i < N_TARGET ; i++) begin
      if (claim_re[i] && claim_id[i] != 0) claim[claim_id[i]-1] = 1'b1;
      if (complete_we[i] && complete_id[i] != 0) complete[complete_id[i]-1] = 1'b1;
    end
  end
  
  rv_plic_gateway #(
    .N_SOURCE (N_SOURCE)
  ) i_rv_plic_gateway (
    .clk_i,
    .rst_ni,
    .src(irq_sources_i),
    .le(le_i),
    .claim(claim),
    .complete(complete),
    .ip(ip)
  );
  
  for (genvar i = 0 ; i < N_TARGET; i++) begin : gen_target
    rv_plic_target #(
      .N_SOURCE  ( N_SOURCE ),
      .MAX_PRIO  ( MAX_PRIO ),
      .ALGORITHM ( "SEQUENTIAL" )
    ) i_target (
      .clk_i,
      .rst_ni,
      .ip(ip),
      .ie(ie_q[i]),
      .prio(prio_q),
      .threshold(threshold_q[i]),
      .irq(eip_targets_o[i]),
      .irq_id(claim_id[i])
    );
  end
  logic [N_TARGET-1:0] threshold_we_o;
  logic [N_TARGET-1:0][PRIOW-1:0] threshold_o;
  logic [N_SOURCE:0][PRIOW-1:0] prio_i, prio_o;
  logic [N_SOURCE:0] prio_we_o;
  
  
  logic [N_TARGET-1:0][N_SOURCE:0] ie_i, ie_o;
  logic [N_TARGET-1:0] ie_we_o;
  plic_regs i_plic_regs (
    .prio_i(prio_i),
    .prio_o(prio_o),
    .prio_we_o(prio_we_o),
    .prio_re_o(), 
    
    .ip_i({ip, 1'b0}),
    .ip_re_o(), 
    .ie_i(ie_i),
    .ie_o(ie_o),
    .ie_we_o(ie_we_o),
    .ie_re_o(), 
    .threshold_i(threshold_q),
    .threshold_o(threshold_o),
    .threshold_we_o(threshold_we_o),
    .threshold_re_o(), 
    .cc_i(claim_id),
    .cc_o(complete_id),
    .cc_we_o(complete_we),
    .cc_re_o(claim_re),
    .req_i,
    .resp_o
  );
  assign prio_i[0] = '0;
  for (genvar i = 0; i < N_TARGET; i++) begin
    assign ie_i[i] = {ie_q[i][N_SOURCE-1:0], 1'b0};
  end
  for (genvar i = 1; i < N_SOURCE + 1; i++) begin
    assign prio_i[i] = prio_q[i - 1];
  end
  
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (~rst_ni) begin
      prio_q <= '0;
      ie_q <= '0;
      threshold_q <= '0;
    end else begin
      
      for (int i = 0; i < N_SOURCE; i++) begin
        prio_q[i] <= prio_we_o[i + 1] ? prio_o[i + 1] : prio_q[i];
      end
      for (int i = 0; i < N_TARGET; i++) begin
        threshold_q[i] <= threshold_we_o[i] ? threshold_o[i] : threshold_q[i];
        ie_q[i] <= ie_we_o[i] ? ie_o[i][N_SOURCE:1] : ie_q[i];
      end
    end
  end
endmodule
module axi2apb_wrap #(
    parameter int unsigned AXI_ADDR_WIDTH   = 32,
    parameter int unsigned AXI_DATA_WIDTH   = 32,
    parameter int unsigned AXI_USER_WIDTH   = 6,
    parameter int unsigned AXI_ID_WIDTH     = 6,
    parameter int unsigned APB_ADDR_WIDTH   = 32,
    parameter int unsigned APB_DATA_WIDTH   = 32
)(
    input logic     clk_i,
    input logic     rst_ni,
    input logic     test_en_i,
    AXI_BUS.Slave   axi_slave,
    APB_BUS.Master  apb_master
);
    
    
    
    generate if (AXI_DATA_WIDTH == APB_DATA_WIDTH) begin
        axi2apb #(
            .AXI4_ADDRESS_WIDTH ( AXI_ADDR_WIDTH ),
            .AXI4_RDATA_WIDTH   ( AXI_DATA_WIDTH ),
            .AXI4_WDATA_WIDTH   ( AXI_DATA_WIDTH ),
            .AXI4_ID_WIDTH      ( AXI_ID_WIDTH   ),
            .AXI4_USER_WIDTH    ( AXI_USER_WIDTH ),
            .BUFF_DEPTH_SLAVE   ( 2              ),
            .APB_ADDR_WIDTH     ( APB_ADDR_WIDTH )
        ) axi2apb_i (
            .ACLK       ( clk_i                  ),
            .ARESETn    ( rst_ni                 ),
            .test_en_i  ( test_en_i              ),
            .AWID_i     ( axi_slave.aw_id        ),
            .AWADDR_i   ( axi_slave.aw_addr      ),
            .AWLEN_i    ( axi_slave.aw_len       ),
            .AWSIZE_i   ( axi_slave.aw_size      ),
            .AWBURST_i  ( axi_slave.aw_burst     ),
            .AWLOCK_i   ( axi_slave.aw_lock      ),
            .AWCACHE_i  ( axi_slave.aw_cache     ),
            .AWPROT_i   ( axi_slave.aw_prot      ),
            .AWREGION_i ( axi_slave.aw_region    ),
            .AWUSER_i   ( axi_slave.aw_user      ),
            .AWQOS_i    ( axi_slave.aw_qos       ),
            .AWVALID_i  ( axi_slave.aw_valid     ),
            .AWREADY_o  ( axi_slave.aw_ready     ),
            .WDATA_i    ( axi_slave.w_data       ),
            .WSTRB_i    ( axi_slave.w_strb       ),
            .WLAST_i    ( axi_slave.w_last       ),
            .WUSER_i    ( axi_slave.w_user       ),
            .WVALID_i   ( axi_slave.w_valid      ),
            .WREADY_o   ( axi_slave.w_ready      ),
            .BID_o      ( axi_slave.b_id         ),
            .BRESP_o    ( axi_slave.b_resp       ),
            .BVALID_o   ( axi_slave.b_valid      ),
            .BUSER_o    ( axi_slave.b_user       ),
            .BREADY_i   ( axi_slave.b_ready      ),
            .ARID_i     ( axi_slave.ar_id        ),
            .ARADDR_i   ( axi_slave.ar_addr      ),
            .ARLEN_i    ( axi_slave.ar_len       ),
            .ARSIZE_i   ( axi_slave.ar_size      ),
            .ARBURST_i  ( axi_slave.ar_burst     ),
            .ARLOCK_i   ( axi_slave.ar_lock      ),
            .ARCACHE_i  ( axi_slave.ar_cache     ),
            .ARPROT_i   ( axi_slave.ar_prot      ),
            .ARREGION_i ( axi_slave.ar_region    ),
            .ARUSER_i   ( axi_slave.ar_user      ),
            .ARQOS_i    ( axi_slave.ar_qos       ),
            .ARVALID_i  ( axi_slave.ar_valid     ),
            .ARREADY_o  ( axi_slave.ar_ready     ),
            .RID_o      ( axi_slave.r_id         ),
            .RDATA_o    ( axi_slave.r_data       ),
            .RRESP_o    ( axi_slave.r_resp       ),
            .RLAST_o    ( axi_slave.r_last       ),
            .RUSER_o    ( axi_slave.r_user       ),
            .RVALID_o   ( axi_slave.r_valid      ),
            .RREADY_i   ( axi_slave.r_ready      ),
            .PENABLE    ( apb_master.penable     ),
            .PWRITE     ( apb_master.pwrite      ),
            .PADDR      ( apb_master.paddr       ),
            .PSEL       ( apb_master.psel        ),
            .PWDATA     ( apb_master.pwdata      ),
            .PRDATA     ( apb_master.prdata      ),
            .PREADY     ( apb_master.pready      ),
            .PSLVERR    ( apb_master.pslverr     )
        );
        end else if (AXI_DATA_WIDTH == 64 && APB_DATA_WIDTH == 32) begin
            axi2apb_64_32  #(
                .AXI4_ADDRESS_WIDTH ( AXI_ADDR_WIDTH ),
                .AXI4_RDATA_WIDTH   ( AXI_DATA_WIDTH ),
                .AXI4_WDATA_WIDTH   ( AXI_DATA_WIDTH ),
                .AXI4_ID_WIDTH      ( AXI_ID_WIDTH   ),
                .AXI4_USER_WIDTH    ( AXI_USER_WIDTH ),
                .BUFF_DEPTH_SLAVE   ( 2              ),
                .APB_ADDR_WIDTH     ( APB_ADDR_WIDTH )
            ) axi2apb_i (
                .ACLK       ( clk_i                  ),
                .ARESETn    ( rst_ni                 ),
                .test_en_i  ( test_en_i              ),
                .AWID_i     ( axi_slave.aw_id        ),
                .AWADDR_i   ( axi_slave.aw_addr      ),
                .AWLEN_i    ( axi_slave.aw_len       ),
                .AWSIZE_i   ( axi_slave.aw_size      ),
                .AWBURST_i  ( axi_slave.aw_burst     ),
                .AWLOCK_i   ( axi_slave.aw_lock      ),
                .AWCACHE_i  ( axi_slave.aw_cache     ),
                .AWPROT_i   ( axi_slave.aw_prot      ),
                .AWREGION_i ( axi_slave.aw_region    ),
                .AWUSER_i   ( axi_slave.aw_user      ),
                .AWQOS_i    ( axi_slave.aw_qos       ),
                .AWVALID_i  ( axi_slave.aw_valid     ),
                .AWREADY_o  ( axi_slave.aw_ready     ),
                .WDATA_i    ( axi_slave.w_data       ),
                .WSTRB_i    ( axi_slave.w_strb       ),
                .WLAST_i    ( axi_slave.w_last       ),
                .WUSER_i    ( axi_slave.w_user       ),
                .WVALID_i   ( axi_slave.w_valid      ),
                .WREADY_o   ( axi_slave.w_ready      ),
                .BID_o      ( axi_slave.b_id         ),
                .BRESP_o    ( axi_slave.b_resp       ),
                .BVALID_o   ( axi_slave.b_valid      ),
                .BUSER_o    ( axi_slave.b_user       ),
                .BREADY_i   ( axi_slave.b_ready      ),
                .ARID_i     ( axi_slave.ar_id        ),
                .ARADDR_i   ( axi_slave.ar_addr      ),
                .ARLEN_i    ( axi_slave.ar_len       ),
                .ARSIZE_i   ( axi_slave.ar_size      ),
                .ARBURST_i  ( axi_slave.ar_burst     ),
                .ARLOCK_i   ( axi_slave.ar_lock      ),
                .ARCACHE_i  ( axi_slave.ar_cache     ),
                .ARPROT_i   ( axi_slave.ar_prot      ),
                .ARREGION_i ( axi_slave.ar_region    ),
                .ARUSER_i   ( axi_slave.ar_user      ),
                .ARQOS_i    ( axi_slave.ar_qos       ),
                .ARVALID_i  ( axi_slave.ar_valid     ),
                .ARREADY_o  ( axi_slave.ar_ready     ),
                .RID_o      ( axi_slave.r_id         ),
                .RDATA_o    ( axi_slave.r_data       ),
                .RRESP_o    ( axi_slave.r_resp       ),
                .RLAST_o    ( axi_slave.r_last       ),
                .RUSER_o    ( axi_slave.r_user       ),
                .RVALID_o   ( axi_slave.r_valid      ),
                .RREADY_i   ( axi_slave.r_ready      ),
                .PENABLE    ( apb_master.penable     ),
                .PWRITE     ( apb_master.pwrite      ),
                .PADDR      ( apb_master.paddr       ),
                .PSEL       ( apb_master.psel        ),
                .PWDATA     ( apb_master.pwdata      ),
                .PRDATA     ( apb_master.prdata      ),
                .PREADY     ( apb_master.pready      ),
                .PSLVERR    ( apb_master.pslverr     )
            );
        end
  endgenerate
endmodule
module axi2apb
#(
    parameter AXI4_ADDRESS_WIDTH = 32,
    parameter AXI4_RDATA_WIDTH   = 32,
    parameter AXI4_WDATA_WIDTH   = 32,
    parameter AXI4_ID_WIDTH      = 16,
    parameter AXI4_USER_WIDTH    = 10,
    parameter AXI_NUMBYTES       = AXI4_WDATA_WIDTH/8,
    parameter BUFF_DEPTH_SLAVE   = 4,
    parameter APB_ADDR_WIDTH     = 32
)
(
    input logic                           ACLK,
    input logic                           ARESETn,
    input logic                           test_en_i,
    input  logic [AXI4_ID_WIDTH-1:0]      AWID_i,
    input  logic [AXI4_ADDRESS_WIDTH-1:0] AWADDR_i,
    input  logic [ 7:0]                   AWLEN_i,
    input  logic [ 2:0]                   AWSIZE_i,
    input  logic [ 1:0]                   AWBURST_i,
    input  logic                          AWLOCK_i,
    input  logic [ 3:0]                   AWCACHE_i,
    input  logic [ 2:0]                   AWPROT_i,
    input  logic [ 3:0]                   AWREGION_i,
    input  logic [ AXI4_USER_WIDTH-1:0]   AWUSER_i,
    input  logic [ 3:0]                   AWQOS_i,
    input  logic                          AWVALID_i,
    output logic                          AWREADY_o,
    input  logic [AXI4_WDATA_WIDTH-1:0]   WDATA_i,
    input  logic [AXI_NUMBYTES-1:0]       WSTRB_i,
    input  logic                          WLAST_i,
    input  logic [AXI4_USER_WIDTH-1:0]    WUSER_i,
    input  logic                          WVALID_i,
    output logic                          WREADY_o,
    output logic   [AXI4_ID_WIDTH-1:0]    BID_o,
    output logic   [ 1:0]                 BRESP_o,
    output logic                          BVALID_o,
    output logic   [AXI4_USER_WIDTH-1:0]  BUSER_o,
    input  logic                          BREADY_i,
    input  logic [AXI4_ID_WIDTH-1:0]      ARID_i,
    input  logic [AXI4_ADDRESS_WIDTH-1:0] ARADDR_i,
    input  logic [ 7:0]                   ARLEN_i,
    input  logic [ 2:0]                   ARSIZE_i,
    input  logic [ 1:0]                   ARBURST_i,
    input  logic                          ARLOCK_i,
    input  logic [ 3:0]                   ARCACHE_i,
    input  logic [ 2:0]                   ARPROT_i,
    input  logic [ 3:0]                   ARREGION_i,
    input  logic [ AXI4_USER_WIDTH-1:0]   ARUSER_i,
    input  logic [ 3:0]                   ARQOS_i,
    input  logic                          ARVALID_i,
    output logic                          ARREADY_o,
    output  logic [AXI4_ID_WIDTH-1:0]     RID_o,
    output  logic [AXI4_RDATA_WIDTH-1:0]  RDATA_o,
    output  logic [ 1:0]                  RRESP_o,
    output  logic                         RLAST_o,
    output  logic [AXI4_USER_WIDTH-1:0]   RUSER_o,
    output  logic                         RVALID_o,
    input   logic                         RREADY_i,
    output logic                          PENABLE,
    output logic                          PWRITE,
    output logic [APB_ADDR_WIDTH-1:0]     PADDR,
    output logic                          PSEL,
    output logic [AXI4_WDATA_WIDTH-1:0]   PWDATA,
    input  logic [AXI4_RDATA_WIDTH-1:0]   PRDATA,
    input  logic                          PREADY,
    input  logic                          PSLVERR
);
    
    
    
    logic [AXI4_ID_WIDTH-1:0]       AWID;
    logic [AXI4_ADDRESS_WIDTH-1:0]  AWADDR;
    logic [ 7:0]                    AWLEN;
    logic [ 2:0]                    AWSIZE;
    logic [ 1:0]                    AWBURST;
    logic                           AWLOCK;
    logic [ 3:0]                    AWCACHE;
    logic [ 2:0]                    AWPROT;
    logic [ 3:0]                    AWREGION;
    logic [ AXI4_USER_WIDTH-1:0]    AWUSER;
    logic [ 3:0]                    AWQOS;
    logic                           AWVALID;
    logic                           AWREADY;
    
    
    
    logic [AXI4_WDATA_WIDTH-1:0]    WDATA;  
    logic [AXI_NUMBYTES-1:0]        WSTRB;  
    logic                           WLAST;  
    logic [AXI4_USER_WIDTH-1:0]     WUSER;  
    logic                           WVALID; 
    logic                           WREADY; 
    
    
    
    logic   [AXI4_ID_WIDTH-1:0]     BID;
    logic   [ 1:0]                  BRESP;
    logic                           BVALID;
    logic   [AXI4_USER_WIDTH-1:0]   BUSER;
    logic                           BREADY;
    
    
    
    logic [AXI4_ID_WIDTH-1:0]       ARID;
    logic [AXI4_ADDRESS_WIDTH-1:0]  ARADDR;
    logic [ 7:0]                    ARLEN;
    logic [ 2:0]                    ARSIZE;
    logic [ 1:0]                    ARBURST;
    logic                           ARLOCK;
    logic [ 3:0]                    ARCACHE;
    logic [ 2:0]                    ARPROT;
    logic [ 3:0]                    ARREGION;
    logic [ AXI4_USER_WIDTH-1:0]    ARUSER;
    logic [ 3:0]                    ARQOS;
    logic                           ARVALID;
    logic                           ARREADY;
    
    
    
    logic [AXI4_ID_WIDTH-1:0]       RID;
    logic [AXI4_RDATA_WIDTH-1:0]    RDATA;
    logic [ 1:0]                    RRESP;
    logic                           RLAST;
    logic [AXI4_USER_WIDTH-1:0]     RUSER;
    logic                           RVALID;
    logic                           RREADY;
  enum logic [2:0] { IDLE,
                     DONE_SINGLE_RD,
                     WAIT_W_PREADY,
                     WAIT_R_PREADY,
                     SEND_B_RESP
                    } CS, NS;
  logic [AXI4_ADDRESS_WIDTH-1:0] address;
  logic sample_RDATA;
  logic [AXI4_RDATA_WIDTH-1:0] RDATA_Q;
  logic read_req;
  logic write_req;
  assign PENABLE = write_req | read_req;
  assign PWRITE  = write_req;
  assign PADDR   = address[APB_ADDR_WIDTH-1:0];
  assign PWDATA  = WDATA;
  assign PSEL    = 1'b1;
   
   axi_aw_buffer #(
       .ID_WIDTH     ( AXI4_ID_WIDTH      ),
       .ADDR_WIDTH   ( AXI4_ADDRESS_WIDTH ),
       .USER_WIDTH   ( AXI4_USER_WIDTH    ),
       .BUFFER_DEPTH ( BUFF_DEPTH_SLAVE   )
   ) slave_aw_buffer_i (
      .clk_i           ( ACLK        ),
      .rst_ni          ( ARESETn     ),
      .test_en_i       ( test_en_i   ),
      .slave_valid_i   ( AWVALID_i   ),
      .slave_addr_i    ( AWADDR_i    ),
      .slave_prot_i    ( AWPROT_i    ),
      .slave_region_i  ( AWREGION_i  ),
      .slave_len_i     ( AWLEN_i     ),
      .slave_size_i    ( AWSIZE_i    ),
      .slave_burst_i   ( AWBURST_i   ),
      .slave_lock_i    ( AWLOCK_i    ),
      .slave_cache_i   ( AWCACHE_i   ),
      .slave_qos_i     ( AWQOS_i     ),
      .slave_id_i      ( AWID_i      ),
      .slave_user_i    ( AWUSER_i    ),
      .slave_ready_o   ( AWREADY_o   ),
      .master_valid_o  ( AWVALID     ),
      .master_addr_o   ( AWADDR      ),
      .master_prot_o   ( AWPROT      ),
      .master_region_o ( AWREGION    ),
      .master_len_o    ( AWLEN       ),
      .master_size_o   ( AWSIZE      ),
      .master_burst_o  ( AWBURST     ),
      .master_lock_o   ( AWLOCK      ),
      .master_cache_o  ( AWCACHE     ),
      .master_qos_o    ( AWQOS       ),
      .master_id_o     ( AWID        ),
      .master_user_o   ( AWUSER      ),
      .master_ready_i  ( AWREADY     )
   );
   
   axi_ar_buffer #(
       .ID_WIDTH     ( AXI4_ID_WIDTH      ),
       .ADDR_WIDTH   ( AXI4_ADDRESS_WIDTH ),
       .USER_WIDTH   ( AXI4_USER_WIDTH    ),
       .BUFFER_DEPTH ( BUFF_DEPTH_SLAVE   )
   ) slave_ar_buffer_i (
      .clk_i           ( ACLK       ),
      .rst_ni          ( ARESETn    ),
      .test_en_i       ( test_en_i  ),
      .slave_valid_i   ( ARVALID_i  ),
      .slave_addr_i    ( ARADDR_i   ),
      .slave_prot_i    ( ARPROT_i   ),
      .slave_region_i  ( ARREGION_i ),
      .slave_len_i     ( ARLEN_i    ),
      .slave_size_i    ( ARSIZE_i   ),
      .slave_burst_i   ( ARBURST_i  ),
      .slave_lock_i    ( ARLOCK_i   ),
      .slave_cache_i   ( ARCACHE_i  ),
      .slave_qos_i     ( ARQOS_i    ),
      .slave_id_i      ( ARID_i     ),
      .slave_user_i    ( ARUSER_i   ),
      .slave_ready_o   ( ARREADY_o  ),
      .master_valid_o  ( ARVALID    ),
      .master_addr_o   ( ARADDR     ),
      .master_prot_o   ( ARPROT     ),
      .master_region_o ( ARREGION   ),
      .master_len_o    ( ARLEN      ),
      .master_size_o   ( ARSIZE     ),
      .master_burst_o  ( ARBURST    ),
      .master_lock_o   ( ARLOCK     ),
      .master_cache_o  ( ARCACHE    ),
      .master_qos_o    ( ARQOS      ),
      .master_id_o     ( ARID       ),
      .master_user_o   ( ARUSER     ),
      .master_ready_i  ( ARREADY    )
   );
   axi_w_buffer #(
       .DATA_WIDTH(AXI4_WDATA_WIDTH),
       .USER_WIDTH(AXI4_USER_WIDTH),
       .BUFFER_DEPTH(BUFF_DEPTH_SLAVE)
   ) slave_w_buffer_i (
        .clk_i          ( ACLK      ),
        .rst_ni         ( ARESETn   ),
        .test_en_i      ( test_en_i ),
        .slave_valid_i  ( WVALID_i  ),
        .slave_data_i   ( WDATA_i   ),
        .slave_strb_i   ( WSTRB_i   ),
        .slave_user_i   ( WUSER_i   ),
        .slave_last_i   ( WLAST_i   ),
        .slave_ready_o  ( WREADY_o  ),
        .master_valid_o ( WVALID    ),
        .master_data_o  ( WDATA     ),
        .master_strb_o  ( WSTRB     ),
        .master_user_o  ( WUSER     ),
        .master_last_o  ( WLAST     ),
        .master_ready_i ( WREADY    )
    );
   axi_r_buffer #(
        .ID_WIDTH     ( AXI4_ID_WIDTH    ),
        .DATA_WIDTH   ( AXI4_RDATA_WIDTH ),
        .USER_WIDTH   ( AXI4_USER_WIDTH  ),
        .BUFFER_DEPTH ( BUFF_DEPTH_SLAVE )
   ) slave_r_buffer_i (
        .clk_i          ( ACLK       ),
        .rst_ni         ( ARESETn    ),
        .test_en_i      ( test_en_i  ),
        .slave_valid_i  ( RVALID     ),
        .slave_data_i   ( RDATA      ),
        .slave_resp_i   ( RRESP      ),
        .slave_user_i   ( RUSER      ),
        .slave_id_i     ( RID        ),
        .slave_last_i   ( RLAST      ),
        .slave_ready_o  ( RREADY     ),
        .master_valid_o ( RVALID_o   ),
        .master_data_o  ( RDATA_o    ),
        .master_resp_o  ( RRESP_o    ),
        .master_user_o  ( RUSER_o    ),
        .master_id_o    ( RID_o      ),
        .master_last_o  ( RLAST_o    ),
        .master_ready_i ( RREADY_i   )
   );
   axi_b_buffer #(
        .ID_WIDTH(AXI4_ID_WIDTH),
        .USER_WIDTH(AXI4_USER_WIDTH),
        .BUFFER_DEPTH(BUFF_DEPTH_SLAVE)
   ) slave_b_buffer (
        .clk_i          ( ACLK      ),
        .rst_ni         ( ARESETn   ),
        .test_en_i      ( test_en_i ),
        .slave_valid_i  ( BVALID    ),
        .slave_resp_i   ( BRESP     ),
        .slave_id_i     ( BID       ),
        .slave_user_i   ( BUSER     ),
        .slave_ready_o  ( BREADY    ),
        .master_valid_o ( BVALID_o  ),
        .master_resp_o  ( BRESP_o   ),
        .master_id_o    ( BID_o     ),
        .master_user_o  ( BUSER_o   ),
        .master_ready_i ( BREADY_i  )
    );
    always_comb begin
      read_req     = 1'b0;
      write_req    = 1'b0;
      address      = '0;
      sample_RDATA = 1'b0;
      ARREADY      = 1'b0;
      AWREADY      = 1'b0;
      WREADY       = 1'b0;
      BVALID       = 1'b0;
      BRESP        = 2'b00;
      BID          = AWID;
      BUSER        = AWUSER;
      RVALID       = 1'b0;
      RLAST        = 1'b0;
      RID          = ARID;
      RUSER        = ARUSER;
      RRESP        = 2'b00;
      RDATA        = RDATA_Q;
      case(CS)
        WAIT_R_PREADY: begin
            read_req     = 1'b1;
            address      = ARADDR[APB_ADDR_WIDTH  - 1 : 0];
            sample_RDATA = PREADY;
            if (PREADY == 1'b1) begin 
               NS = DONE_SINGLE_RD;
            end
        end
        WAIT_W_PREADY: begin
            write_req   = 1'b1;
            address     = AWADDR[APB_ADDR_WIDTH - 1:0];
            
            if (PREADY == 1'b1) begin 
                NS = SEND_B_RESP;
            end
        end
        IDLE: begin
            if (ARVALID == 1'b1) begin
                read_req     = 1'b1;
                address      = ARADDR[APB_ADDR_WIDTH - 1:0];;
                sample_RDATA = PREADY;
                if(PREADY == 1'b1) begin 
                    NS   = DONE_SINGLE_RD;
                end else begin 
                    NS = WAIT_R_PREADY;
                end
            end else begin
                if (AWVALID) begin
                    address =  AWADDR[APB_ADDR_WIDTH - 1:0];
                    if (WVALID) begin
                        write_req = 1'b1;
                        
                        if (PREADY == 1'b1) begin
                            NS = SEND_B_RESP;
                        end else begin 
                           NS = WAIT_W_PREADY;
                        end
                    end else begin 
                        write_req       = 1'b0;
                        address         = '0;
                        NS              = IDLE;
                    end
                end
            end
        end
        SEND_B_RESP: begin
            BVALID   = 1'b1;
            address  = '0;
            if (BREADY) begin
                NS      = IDLE;
                AWREADY = 1'b1;
                WREADY  = 1'b1;
            end
        end
        DONE_SINGLE_RD: begin
            RVALID    = 1'b1;
            RLAST     = 1;
            address   = '0;
            if (RREADY) begin 
                NS = IDLE;
                ARREADY = 1'b1;
            end
        end
        default: NS = IDLE;
      endcase
    end
    always_ff @(posedge ACLK, negedge ARESETn) begin
        if (ARESETn == 1'b0) begin
            CS      <= IDLE;
            RDATA_Q <= '0;
        end else begin
            CS      <= NS;
            if (sample_RDATA)
                RDATA_Q <= PRDATA;
        end
    end
endmodule
module axi2apb_64_32 #(
    parameter int unsigned AXI4_ADDRESS_WIDTH = 32,
    parameter int unsigned AXI4_RDATA_WIDTH   = 64,
    parameter int unsigned AXI4_WDATA_WIDTH   = 64,
    parameter int unsigned AXI4_ID_WIDTH      = 16,
    parameter int unsigned AXI4_USER_WIDTH    = 10,
    parameter int unsigned AXI_NUMBYTES       = AXI4_WDATA_WIDTH/8,
    parameter int unsigned BUFF_DEPTH_SLAVE   = 4,
    parameter int unsigned APB_NUM_SLAVES     = 8,
    parameter int unsigned APB_ADDR_WIDTH     = 12
)
(
    input logic                           ACLK,
    input logic                           ARESETn,
    input logic                           test_en_i,
    
    
    
    
    input  logic [AXI4_ID_WIDTH-1:0]       AWID_i     ,
    input  logic [AXI4_ADDRESS_WIDTH-1:0]  AWADDR_i   ,
    input  logic [ 7:0]                    AWLEN_i    ,
    input  logic [ 2:0]                    AWSIZE_i   ,
    input  logic [ 1:0]                    AWBURST_i  ,
    input  logic                           AWLOCK_i   ,
    input  logic [ 3:0]                    AWCACHE_i  ,
    input  logic [ 2:0]                    AWPROT_i   ,
    input  logic [ 3:0]                    AWREGION_i ,
    input  logic [ AXI4_USER_WIDTH-1:0]    AWUSER_i   ,
    input  logic [ 3:0]                    AWQOS_i    ,
    input  logic                           AWVALID_i  ,
    output logic                           AWREADY_o  ,
    
    
    input  logic [AXI_NUMBYTES-1:0][7:0]   WDATA_i    ,
    input  logic [AXI_NUMBYTES-1:0]        WSTRB_i    ,
    input  logic                           WLAST_i    ,
    input  logic [AXI4_USER_WIDTH-1:0]     WUSER_i    ,
    input  logic                           WVALID_i   ,
    output logic                           WREADY_o   ,
    
    
    output logic   [AXI4_ID_WIDTH-1:0]     BID_o      ,
    output logic   [ 1:0]                  BRESP_o    ,
    output logic                           BVALID_o   ,
    output logic   [AXI4_USER_WIDTH-1:0]   BUSER_o    ,
    input  logic                           BREADY_i   ,
    
    
    input  logic [AXI4_ID_WIDTH-1:0]       ARID_i     ,
    input  logic [AXI4_ADDRESS_WIDTH-1:0]  ARADDR_i   ,
    input  logic [ 7:0]                    ARLEN_i    ,
    input  logic [ 2:0]                    ARSIZE_i   ,
    input  logic [ 1:0]                    ARBURST_i  ,
    input  logic                           ARLOCK_i   ,
    input  logic [ 3:0]                    ARCACHE_i  ,
    input  logic [ 2:0]                    ARPROT_i   ,
    input  logic [ 3:0]                    ARREGION_i ,
    input  logic [ AXI4_USER_WIDTH-1:0]    ARUSER_i   ,
    input  logic [ 3:0]                    ARQOS_i    ,
    input  logic                           ARVALID_i  ,
    output logic                           ARREADY_o  ,
    
    
    output  logic [AXI4_ID_WIDTH-1:0]      RID_o      ,
    output  logic [AXI4_RDATA_WIDTH-1:0]   RDATA_o    ,
    output  logic [ 1:0]                   RRESP_o    ,
    output  logic                          RLAST_o    ,
    output  logic [AXI4_USER_WIDTH-1:0]    RUSER_o    ,
    output  logic                          RVALID_o   ,
    input   logic                          RREADY_i   ,
    
    output logic                           PENABLE    ,
    output logic                           PWRITE     ,
    output logic [APB_ADDR_WIDTH-1:0]      PADDR      ,
    output logic                           PSEL       ,
    output logic [31:0]                    PWDATA     ,
    input  logic [31:0]                    PRDATA     ,
    input  logic                           PREADY     ,
    input  logic                           PSLVERR
);
    
    
    
    logic [AXI4_ID_WIDTH-1:0]      AWID;
    logic [AXI4_ADDRESS_WIDTH-1:0] AWADDR;
    logic [ 7:0]                   AWLEN;
    logic [ 2:0]                   AWSIZE;
    logic [ 1:0]                   AWBURST;
    logic                          AWLOCK;
    logic [ 3:0]                   AWCACHE;
    logic [ 2:0]                   AWPROT;
    logic [ 3:0]                   AWREGION;
    logic [ AXI4_USER_WIDTH-1:0]   AWUSER;
    logic [ 3:0]                   AWQOS;
    logic                          AWVALID;
    logic                          AWREADY;
    
    
    
    logic [1:0][31:0]              WDATA;  
    logic [AXI_NUMBYTES-1:0]       WSTRB;  
    logic                          WLAST;  
    logic [AXI4_USER_WIDTH-1:0]    WUSER;  
    logic                          WVALID; 
    logic                          WREADY; 
    
    
    
    logic [AXI4_ID_WIDTH-1:0]      BID;
    logic [ 1:0]                   BRESP;
    logic                          BVALID;
    logic [AXI4_USER_WIDTH-1:0]    BUSER;
    logic                          BREADY;
    
    
    
    logic [AXI4_ID_WIDTH-1:0]      ARID;
    logic [AXI4_ADDRESS_WIDTH-1:0] ARADDR;
    logic [ 7:0]                   ARLEN;
    logic [ 2:0]                   ARSIZE;
    logic [ 1:0]                   ARBURST;
    logic                          ARLOCK;
    logic [ 3:0]                   ARCACHE;
    logic [ 2:0]                   ARPROT;
    logic [ 3:0]                   ARREGION;
    logic [ AXI4_USER_WIDTH-1:0]   ARUSER;
    logic [ 3:0]                   ARQOS;
    logic                          ARVALID;
    logic                          ARREADY;
    
    
    
    logic [AXI4_ID_WIDTH-1:0]    RID;
    logic [1:0][31:0]            RDATA;
    logic [ 1:0]                 RRESP;
    logic                        RLAST;
    logic [AXI4_USER_WIDTH-1:0]  RUSER;
    logic                        RVALID;
    logic                        RREADY;
    enum logic [3:0] { IDLE,
                       SINGLE_RD, SINGLE_RD_64,
                       BURST_RD_1, BURST_RD, BURST_RD_64,
                       BURST_WR, BURST_WR_64,
                       SINGLE_WR,SINGLE_WR_64,
                       WAIT_R_PREADY, WAIT_W_PREADY
                      } CS, NS;
    logic        W_word_sel;
    logic [APB_ADDR_WIDTH-1:0] address;
    logic        read_req;
    logic        write_req;
    logic        sample_AR;
    logic [8:0]  ARLEN_Q;
    logic        decr_ARLEN;
    logic        sample_AW;
    logic [8:0]  AWLEN_Q;
    logic        decr_AWLEN;
    logic [AXI4_ADDRESS_WIDTH-1:0] ARADDR_Q;
    logic                          incr_ARADDR;
    logic [AXI4_ADDRESS_WIDTH-1:0] AWADDR_Q;
    logic                          incr_AWADDR;
    logic        sample_RDATA_0; 
    logic        sample_RDATA_1; 
    logic [31:0] RDATA_Q_0;
    logic [31:0] RDATA_Q_1;
    assign PENABLE = write_req | read_req;
    assign PWRITE  = write_req;
    assign PADDR   = address[APB_ADDR_WIDTH-1:0];
    assign PWDATA  = WDATA[W_word_sel];
    assign PSEL    = 1'b1;
    
    axi_aw_buffer #(
        .ID_WIDTH     ( AXI4_ID_WIDTH      ),
        .ADDR_WIDTH   ( AXI4_ADDRESS_WIDTH ),
        .USER_WIDTH   ( AXI4_USER_WIDTH    ),
        .BUFFER_DEPTH ( BUFF_DEPTH_SLAVE   )
    ) slave_aw_buffer_i (
       .clk_i           ( ACLK        ),
       .rst_ni          ( ARESETn     ),
       .test_en_i       ( test_en_i   ),
       .slave_valid_i   ( AWVALID_i   ),
       .slave_addr_i    ( AWADDR_i    ),
       .slave_prot_i    ( AWPROT_i    ),
       .slave_region_i  ( AWREGION_i  ),
       .slave_len_i     ( AWLEN_i     ),
       .slave_size_i    ( AWSIZE_i    ),
       .slave_burst_i   ( AWBURST_i   ),
       .slave_lock_i    ( AWLOCK_i    ),
       .slave_cache_i   ( AWCACHE_i   ),
       .slave_qos_i     ( AWQOS_i     ),
       .slave_id_i      ( AWID_i      ),
       .slave_user_i    ( AWUSER_i    ),
       .slave_ready_o   ( AWREADY_o   ),
       .master_valid_o  ( AWVALID     ),
       .master_addr_o   ( AWADDR      ),
       .master_prot_o   ( AWPROT      ),
       .master_region_o ( AWREGION    ),
       .master_len_o    ( AWLEN       ),
       .master_size_o   ( AWSIZE      ),
       .master_burst_o  ( AWBURST     ),
       .master_lock_o   ( AWLOCK      ),
       .master_cache_o  ( AWCACHE     ),
       .master_qos_o    ( AWQOS       ),
       .master_id_o     ( AWID        ),
       .master_user_o   ( AWUSER      ),
       .master_ready_i  ( AWREADY     )
    );
    
    axi_ar_buffer #(
        .ID_WIDTH       ( AXI4_ID_WIDTH      ),
        .ADDR_WIDTH     ( AXI4_ADDRESS_WIDTH ),
        .USER_WIDTH     ( AXI4_USER_WIDTH    ),
        .BUFFER_DEPTH   ( BUFF_DEPTH_SLAVE   )
    ) slave_ar_buffer_i (
       .clk_i           ( ACLK       ),
       .rst_ni          ( ARESETn    ),
       .test_en_i       ( test_en_i  ),
       .slave_valid_i   ( ARVALID_i  ),
       .slave_addr_i    ( ARADDR_i   ),
       .slave_prot_i    ( ARPROT_i   ),
       .slave_region_i  ( ARREGION_i ),
       .slave_len_i     ( ARLEN_i    ),
       .slave_size_i    ( ARSIZE_i   ),
       .slave_burst_i   ( ARBURST_i  ),
       .slave_lock_i    ( ARLOCK_i   ),
       .slave_cache_i   ( ARCACHE_i  ),
       .slave_qos_i     ( ARQOS_i    ),
       .slave_id_i      ( ARID_i     ),
       .slave_user_i    ( ARUSER_i   ),
       .slave_ready_o   ( ARREADY_o  ),
       .master_valid_o  ( ARVALID    ),
       .master_addr_o   ( ARADDR     ),
       .master_prot_o   ( ARPROT     ),
       .master_region_o ( ARREGION   ),
       .master_len_o    ( ARLEN      ),
       .master_size_o   ( ARSIZE     ),
       .master_burst_o  ( ARBURST    ),
       .master_lock_o   ( ARLOCK     ),
       .master_cache_o  ( ARCACHE    ),
       .master_qos_o    ( ARQOS      ),
       .master_id_o     ( ARID       ),
       .master_user_o   ( ARUSER     ),
       .master_ready_i  ( ARREADY    )
    );
    axi_w_buffer #(
        .DATA_WIDTH   ( AXI4_WDATA_WIDTH ),
        .USER_WIDTH   ( AXI4_USER_WIDTH  ),
        .BUFFER_DEPTH ( BUFF_DEPTH_SLAVE )
    ) slave_w_buffer_i (
         .clk_i          ( ACLK      ),
         .rst_ni         ( ARESETn   ),
         .test_en_i      ( test_en_i ),
         .slave_valid_i  ( WVALID_i  ),
         .slave_data_i   ( WDATA_i   ),
         .slave_strb_i   ( WSTRB_i   ),
         .slave_user_i   ( WUSER_i   ),
         .slave_last_i   ( WLAST_i   ),
         .slave_ready_o  ( WREADY_o  ),
         .master_valid_o ( WVALID    ),
         .master_data_o  ( WDATA     ),
         .master_strb_o  ( WSTRB     ),
         .master_user_o  ( WUSER     ),
         .master_last_o  ( WLAST     ),
         .master_ready_i ( WREADY    )
    );
    axi_r_buffer #(
         .ID_WIDTH     ( AXI4_ID_WIDTH    ),
         .DATA_WIDTH   ( AXI4_RDATA_WIDTH ),
         .USER_WIDTH   ( AXI4_USER_WIDTH  ),
         .BUFFER_DEPTH ( BUFF_DEPTH_SLAVE )
    ) slave_r_buffer_i (
         .clk_i          ( ACLK       ),
         .rst_ni         ( ARESETn    ),
         .test_en_i      ( test_en_i  ),
         .slave_valid_i  ( RVALID     ),
         .slave_data_i   ( RDATA      ),
         .slave_resp_i   ( RRESP      ),
         .slave_user_i   ( RUSER      ),
         .slave_id_i     ( RID        ),
         .slave_last_i   ( RLAST      ),
         .slave_ready_o  ( RREADY     ),
         .master_valid_o ( RVALID_o   ),
         .master_data_o  ( RDATA_o    ),
         .master_resp_o  ( RRESP_o    ),
         .master_user_o  ( RUSER_o    ),
         .master_id_o    ( RID_o      ),
         .master_last_o  ( RLAST_o    ),
         .master_ready_i ( RREADY_i   )
    );
    axi_b_buffer #(
        .ID_WIDTH       ( AXI4_ID_WIDTH    ),
        .USER_WIDTH     ( AXI4_USER_WIDTH  ),
        .BUFFER_DEPTH   ( BUFF_DEPTH_SLAVE )
    ) slave_b_buffer_i (
        .clk_i          ( ACLK      ),
        .rst_ni         ( ARESETn   ),
        .test_en_i      ( test_en_i ),
        .slave_valid_i  ( BVALID    ),
        .slave_resp_i   ( BRESP     ),
        .slave_id_i     ( BID       ),
        .slave_user_i   ( BUSER     ),
        .slave_ready_o  ( BREADY    ),
        .master_valid_o ( BVALID_o  ),
        .master_resp_o  ( BRESP_o   ),
        .master_id_o    ( BID_o     ),
        .master_user_o  ( BUSER_o   ),
        .master_ready_i ( BREADY_i  )
    );
    always_comb begin
        read_req   = 1'b0;
        write_req  = 1'b0;
        W_word_sel = 1'b0; 
        sample_AW  = 1'b0;
        decr_AWLEN = 1'b0;
        sample_AR  = 1'b0;
        decr_ARLEN = 1'b0;
        incr_AWADDR = 1'b0;
        incr_ARADDR = 1'b0;
        sample_RDATA_0 = 1'b0;
        sample_RDATA_1 = 1'b0;
        ARREADY = 1'b0;
        AWREADY = 1'b0;
        WREADY  = 1'b0;
        RDATA   = '0;
        BVALID = 1'b0;
        BRESP  = 2'b00;
        BID    = AWID;
        BUSER  = AWUSER;
        RVALID = 1'b0;
        RLAST  = 1'b0;
        RID    = ARID;
        RUSER  = ARUSER;
        RRESP  = 2'b00;
        case(CS)
            WAIT_R_PREADY: begin
                sample_AR = 1'b0;
                read_req  = 1'b1;
                address   = ARADDR;
                if (PREADY == 1'b1) begin
                    if (ARLEN == 0) begin
                        case (ARSIZE)
                            3'h3: begin
                                NS = SINGLE_RD_64;
                                if (ARADDR[2:0] == 3'h4)
                                    sample_RDATA_1 = 1'b1;
                                else  sample_RDATA_0 = 1'b1;
                            end
                            default: begin
                                NS = SINGLE_RD;
                                if (ARADDR[2:0] == 3'h4)
                                    sample_RDATA_1 = 1'b1;
                                else
                                    sample_RDATA_0 = 1'b1;
                                end
                            endcase
                    end else begin 
                       NS             = BURST_RD_64;
                       sample_RDATA_0 = 1'b1;
                       decr_ARLEN     = 1'b1;
                       incr_ARADDR    = 1'b1;
                    end
                end else begin 
                    NS = WAIT_R_PREADY;
                end
            end
            WAIT_W_PREADY: begin
                address   = AWADDR;
                write_req = 1'b1;
                if (AWADDR[2:0] == 3'h4)
                    W_word_sel = 1'b1;
                else
                    W_word_sel = 1'b0;
                
                if (PREADY == 1'b1) begin 
                    if (AWLEN == 0) begin 
                        case (AWSIZE)
                            3'h3: NS = SINGLE_WR_64;
                            default: NS = SINGLE_WR;
                        endcase
                    end else begin 
                        sample_AW = 1'b1;
                        NS        = BURST_WR_64;
                    end
                end else begin 
                    NS = WAIT_W_PREADY;
                end
            end
            IDLE: begin
                if (ARVALID == 1'b1)  begin
                    sample_AR = 1'b1;
                    read_req  = 1'b1;
                    address   = ARADDR;
                    if (PREADY == 1'b1) begin 
                        if (ARLEN == 0) begin
                            case (ARSIZE)
                                3'h3: begin
                                    NS = SINGLE_RD_64;
                                    if (ARADDR[2:0] == 4)
                                        sample_RDATA_1 = 1'b1;
                                    else
                                        sample_RDATA_0 = 1'b1;
                                end
                                default: begin
                                    NS = SINGLE_RD;
                                    if (ARADDR[2:0] == 4)
                                        sample_RDATA_1 = 1'b1;
                                    else
                                        sample_RDATA_0 = 1'b1;
                                    end
                            endcase end else begin 
                            NS             = BURST_RD_64;
                            sample_RDATA_0 = 1'b1;
                        end
                    end else begin 
                        NS = WAIT_R_PREADY;
                    end
                end else begin
                    if (AWVALID) begin 
                        if (WVALID) begin 
                            write_req = 1'b1;
                            address   = AWADDR;
                            if (AWADDR[2:0] == 3'h4)
                                W_word_sel = 1'b1;
                            else
                                W_word_sel = 1'b0;
                          
                            if (PREADY == 1'b1) begin
                                  if(AWLEN == 0) begin 
                                        case(AWSIZE)
                                            3'h3: NS = SINGLE_WR_64;
                                            default: NS = SINGLE_WR;
                                        endcase
                                  end else begin 
                                        sample_AW   = 1'b1;
                                        if ((AWADDR[2:0] == 3'h4) && (WSTRB[7:4] == 0))
                                          incr_AWADDR = 1'b0;
                                        else
                                          incr_AWADDR = 1'b1;
                                        NS = BURST_WR_64;
                                  end
                            end else begin
                                NS = WAIT_W_PREADY;
                            end
                        end else begin 
                            write_req = 1'b0;
                            address   = '0;
                            NS        = IDLE;
                        end
                    end else begin
                        NS = IDLE;
                        address =  '0;
                    end
                end
            end
            SINGLE_WR_64: begin
                address    = AWADDR + 4;
                W_word_sel = 1'b1; 
                write_req  = WVALID;
                if (WVALID) begin
                    if (PREADY == 1'b1)
                        NS = SINGLE_WR;
                    else
                        NS = SINGLE_WR_64;
                end else begin
                    NS = SINGLE_WR_64;
                end
            end
            SINGLE_WR:  begin
                BVALID   = 1'b1;
                address  = '0;
                if (BREADY)  begin
                    NS      = IDLE;
                    AWREADY = 1'b1;
                    WREADY  = 1'b1;
                end else begin
                    NS = SINGLE_WR;
                end
            end
            BURST_WR_64: begin
                W_word_sel = 1'b1; 
                write_req  = WVALID & (|WSTRB[7:4]);
                address    = AWADDR_Q; 
                if (WVALID) begin
                    if (&WSTRB[7:4]) begin
                        if(PREADY == 1'b1) begin
                            NS          = BURST_WR;
                            WREADY      = 1'b1; 
                            decr_AWLEN  = 1'b1; 
                            incr_AWADDR = 1'b1; 
                        end else begin
                            NS = BURST_WR_64;
                        end
                    end else begin
                        NS = BURST_WR;
                        WREADY      = 1'b1; 
                        decr_AWLEN  = 1'b1; 
                        incr_AWADDR = 1'b1; 
                    end
                end else begin
                    NS = BURST_WR_64;
                end
            end
            BURST_WR: begin
                address = AWADDR_Q; 
                if (AWLEN_Q == 0) begin 
                    BVALID = 1'b1;
                    if (BREADY) begin
                      NS      = IDLE;
                      AWREADY = 1'b1;
                    end else
                      NS = BURST_WR;
                end else begin 
                    W_word_sel = 1'b0; 
                    write_req  = WVALID & (&WSTRB[3:0]);
                    if (WVALID) begin
                        if (PREADY == 1'b1) begin
                            NS          = BURST_WR_64;
                            incr_AWADDR = 1'b1;
                            decr_AWLEN  = 1'b1; 
                          end else
                            NS = BURST_WR;
                    end else begin
                        NS = BURST_WR_64;
                    end
              end
            end
            BURST_RD_64: begin
               read_req = 1'b1;
               address  = ARADDR_Q;
                if (ARLEN_Q == 0) begin 
                    NS      = IDLE;
                    ARREADY = 1'b1;
                end else begin
                    if (PREADY == 1'b1) begin 
                        decr_ARLEN     = 1'b1;
                        sample_RDATA_1 = 1'b1;
                        NS = BURST_RD;
                        if (ARADDR_Q[2:0] == 3'h4)
                          incr_ARADDR = 1'b1;
                        else
                          incr_ARADDR = 1'b0;
                      end
                    else  begin
                        NS = BURST_RD_64;
                    end
                 end
            end
            BURST_RD: begin
                RVALID   = 1'b1;
                RDATA[0] = RDATA_Q_0;
                RDATA[1] = RDATA_Q_1;
                RLAST    = (ARLEN_Q == 0) ? 1'b1 : 1'b0;
                address  = ARADDR_Q;
                if (RREADY) begin 
                    if (ARLEN_Q == 0) begin 
                        NS      = IDLE;
                        ARREADY = 1'b1;
                    end else begin 
                        read_req = 1'b1;
                        if (PREADY == 1'b1) begin 
                            sample_RDATA_0 = 1'b1;
                            NS             = BURST_RD_64;
                            incr_ARADDR    = 1'b1;
                            decr_ARLEN     = 1'b1;
                        end else begin
                            NS = BURST_RD_1;
                        end
                    end
                end else begin 
                    NS = BURST_RD;
                end
            end
            BURST_RD_1: begin
                read_req = 1'b1;
                address  = ARADDR_Q;
                if (PREADY == 1'b1) begin 
                    sample_RDATA_0 = 1'b1;
                    NS             = BURST_RD_64;
                    incr_ARADDR    = 1'b1;
                    decr_ARLEN     = 1'b1;
                end else begin
                    NS = BURST_RD_1;
                end
            end
            SINGLE_RD: begin
                RVALID   = 1'b1;
                RDATA[0] = RDATA_Q_0;
                RDATA[1] = RDATA_Q_1;
                RLAST    = 1;
                address  = '0;
                if (RREADY) begin 
                    NS      = IDLE;
                    ARREADY = 1'b1;
                end else begin 
                    NS = SINGLE_RD;
                end
            end
            SINGLE_RD_64: begin
                read_req       = 1'b1;
                address        = ARADDR + 4;
                if (PREADY == 1'b1) begin 
                    NS = SINGLE_RD;
                    if(ARADDR[2:0] == 3'h4)
                        sample_RDATA_0 = 1'b1;
                    else
                        sample_RDATA_1 = 1'b1;
                end else begin
                  NS = SINGLE_RD_64;
                end
            end
            default: begin
                NS      = IDLE;
                address = '0;
            end
        endcase
    end
    
    
    
    always_ff @(posedge ACLK, negedge ARESETn) begin
        if (ARESETn == 1'b0) begin
            CS        <= IDLE;
            
            ARLEN_Q   <= '0;
            AWADDR_Q  <= '0;
            
            AWLEN_Q   <= '0;
            RDATA_Q_0 <= '0;
            RDATA_Q_1 <= '0;
            ARADDR_Q  <= '0;
        end else  begin
            CS <= NS;
            if (sample_AR) begin
                ARLEN_Q <= {ARLEN,1'b0} + 2;
            end else if (decr_ARLEN) begin
                ARLEN_Q <= ARLEN_Q - 1;
            end
            if (sample_RDATA_0)
                RDATA_Q_0 <= PRDATA;
            if (sample_RDATA_1)
                RDATA_Q_1 <= PRDATA;
            case ({sample_AW, decr_AWLEN})
                2'b00: AWLEN_Q <= AWLEN_Q;
                2'b01: AWLEN_Q <= AWLEN_Q - 1;
                2'b10: AWLEN_Q <= {AWLEN, 1'b0} + 1;
                2'b11: AWLEN_Q <= {AWLEN, 1'b0};
            endcase
            case ({sample_AW, incr_AWADDR})
                2'b00: AWADDR_Q <= AWADDR_Q;
                2'b01: AWADDR_Q <= AWADDR_Q + 4;
                2'b10: AWADDR_Q <= {AWADDR[AXI4_ADDRESS_WIDTH-1:3], 3'b000};
                2'b11: AWADDR_Q <= {AWADDR[AXI4_ADDRESS_WIDTH-1:3], 3'b000} + 4;
            endcase
            case({sample_AR, incr_ARADDR})
                2'b00: ARADDR_Q <= ARADDR_Q;
                2'b01: ARADDR_Q <= ARADDR_Q + 4;
                2'b10: ARADDR_Q <= {ARADDR[AXI4_ADDRESS_WIDTH-1:3], 3'b000};
                2'b11: ARADDR_Q <= {ARADDR[AXI4_ADDRESS_WIDTH-1:3], 3'b000} + 4;
            endcase
        end
    end
endmodule
module axi_w_buffer #(
    parameter int DATA_WIDTH   = -1,
    parameter int USER_WIDTH   = -1,
    parameter int BUFFER_DEPTH = -1,
    parameter int STRB_WIDTH   = DATA_WIDTH/8   
)(
    input logic                   clk_i,
    input logic                   rst_ni,
    input logic                   test_en_i,
    input logic                   slave_valid_i,
    input logic  [DATA_WIDTH-1:0] slave_data_i,
    input logic  [STRB_WIDTH-1:0] slave_strb_i,
    input logic  [USER_WIDTH-1:0] slave_user_i,
    input logic                   slave_last_i,
    output logic                  slave_ready_o,
    output logic                  master_valid_o,
    output logic [DATA_WIDTH-1:0] master_data_o,
    output logic [STRB_WIDTH-1:0] master_strb_o,
    output logic [USER_WIDTH-1:0] master_user_o,
    output logic                  master_last_o,
    input  logic                  master_ready_i
);
    logic [DATA_WIDTH+STRB_WIDTH+USER_WIDTH:0] s_data_in;
    logic [DATA_WIDTH+STRB_WIDTH+USER_WIDTH:0] s_data_out;
    assign s_data_in = { slave_user_i,  slave_strb_i,  slave_data_i,  slave_last_i  };
    assign             { master_user_o, master_strb_o, master_data_o, master_last_o } = s_data_out;
    axi_single_slice #(.BUFFER_DEPTH(BUFFER_DEPTH), .DATA_WIDTH(1+DATA_WIDTH+STRB_WIDTH+USER_WIDTH)) i_axi_single_slice (
      .clk_i      ( clk_i          ),
      .rst_ni     ( rst_ni         ),
      .testmode_i ( test_en_i      ),
      .valid_i    ( slave_valid_i  ),
      .ready_o    ( slave_ready_o  ),
      .data_i     ( s_data_in      ),
      .ready_i    ( master_ready_i ),
      .valid_o    ( master_valid_o ),
      .data_o     ( s_data_out     )
    );
endmodule
module axi_b_buffer #(
    parameter int ID_WIDTH     = -1,
    parameter int USER_WIDTH   = -1,
    parameter int BUFFER_DEPTH = -1
)(
   input logic                   clk_i,
   input logic                   rst_ni,
   input logic                   test_en_i,
   input logic                   slave_valid_i,
   input logic  [1:0]            slave_resp_i,
   input logic  [ID_WIDTH-1:0]   slave_id_i,
   input logic  [USER_WIDTH-1:0] slave_user_i,
   output logic                  slave_ready_o,
   output logic                  master_valid_o,
   output logic [1:0]            master_resp_o,
   output logic [ID_WIDTH-1:0]   master_id_o,
   output logic [USER_WIDTH-1:0] master_user_o,
   input  logic                  master_ready_i
);
    logic [2+USER_WIDTH+ID_WIDTH-1:0] s_data_in;
    logic [2+USER_WIDTH+ID_WIDTH-1:0] s_data_out;
    assign s_data_in = {slave_id_i,  slave_user_i,  slave_resp_i};
    assign             {master_id_o, master_user_o, master_resp_o} = s_data_out;
    axi_single_slice #(.BUFFER_DEPTH(BUFFER_DEPTH), .DATA_WIDTH(2+USER_WIDTH+ID_WIDTH)) i_axi_single_slice (
      .clk_i      ( clk_i          ),
      .rst_ni     ( rst_ni         ),
      .testmode_i ( test_en_i      ),
      .valid_i    ( slave_valid_i  ),
      .ready_o    ( slave_ready_o  ),
      .data_i     ( s_data_in      ),
      .ready_i    ( master_ready_i ),
      .valid_o    ( master_valid_o ),
      .data_o     ( s_data_out     )
    );
endmodule
module axi_slice_wrap #(
    parameter AXI_ADDR_WIDTH    = 32,
    parameter AXI_DATA_WIDTH    = 64,
    parameter AXI_USER_WIDTH    = 6,
    parameter AXI_ID_WIDTH      = 3,
    parameter SLICE_DEPTH       = 2,
    parameter AXI_STRB_WIDTH    = AXI_DATA_WIDTH/8
)(
    input logic    clk_i,    
    input logic    rst_ni,  
    input logic    test_en_i,
    AXI_BUS.Slave  axi_slave,
    AXI_BUS.Master axi_master
);
    axi_slice #(
        .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH               ),
        .AXI_DATA_WIDTH ( AXI_DATA_WIDTH               ),
        .AXI_USER_WIDTH ( AXI_USER_WIDTH               ),
        .AXI_ID_WIDTH   ( AXI_ID_WIDTH                 ),
        .SLICE_DEPTH    ( SLICE_DEPTH                  ),
        .AXI_STRB_WIDTH ( AXI_STRB_WIDTH               )
    ) i_axi_slice (
        .axi_slave_aw_valid_i   ( axi_slave.aw_valid   ),
        .axi_slave_aw_addr_i    ( axi_slave.aw_addr    ),
        .axi_slave_aw_prot_i    ( axi_slave.aw_prot    ),
        .axi_slave_aw_region_i  ( axi_slave.aw_region  ),
        .axi_slave_aw_len_i     ( axi_slave.aw_len     ),
        .axi_slave_aw_size_i    ( axi_slave.aw_size    ),
        .axi_slave_aw_burst_i   ( axi_slave.aw_burst   ),
        .axi_slave_aw_lock_i    ( axi_slave.aw_lock    ),
        .axi_slave_aw_cache_i   ( axi_slave.aw_cache   ),
        .axi_slave_aw_qos_i     ( axi_slave.aw_qos     ),
        .axi_slave_aw_id_i      ( axi_slave.aw_id      ),
        .axi_slave_aw_user_i    ( axi_slave.aw_user    ),
        .axi_slave_aw_ready_o   ( axi_slave.aw_ready   ),
        .axi_slave_ar_valid_i   ( axi_slave.ar_valid   ),
        .axi_slave_ar_addr_i    ( axi_slave.ar_addr    ),
        .axi_slave_ar_prot_i    ( axi_slave.ar_prot    ),
        .axi_slave_ar_region_i  ( axi_slave.ar_region  ),
        .axi_slave_ar_len_i     ( axi_slave.ar_len     ),
        .axi_slave_ar_size_i    ( axi_slave.ar_size    ),
        .axi_slave_ar_burst_i   ( axi_slave.ar_burst   ),
        .axi_slave_ar_lock_i    ( axi_slave.ar_lock    ),
        .axi_slave_ar_cache_i   ( axi_slave.ar_cache   ),
        .axi_slave_ar_qos_i     ( axi_slave.ar_qos     ),
        .axi_slave_ar_id_i      ( axi_slave.ar_id      ),
        .axi_slave_ar_user_i    ( axi_slave.ar_user    ),
        .axi_slave_ar_ready_o   ( axi_slave.ar_ready   ),
        .axi_slave_w_valid_i    ( axi_slave.w_valid    ),
        .axi_slave_w_data_i     ( axi_slave.w_data     ),
        .axi_slave_w_strb_i     ( axi_slave.w_strb     ),
        .axi_slave_w_user_i     ( axi_slave.w_user     ),
        .axi_slave_w_last_i     ( axi_slave.w_last     ),
        .axi_slave_w_ready_o    ( axi_slave.w_ready    ),
        .axi_slave_r_valid_o    ( axi_slave.r_valid    ),
        .axi_slave_r_data_o     ( axi_slave.r_data     ),
        .axi_slave_r_resp_o     ( axi_slave.r_resp     ),
        .axi_slave_r_last_o     ( axi_slave.r_last     ),
        .axi_slave_r_id_o       ( axi_slave.r_id       ),
        .axi_slave_r_user_o     ( axi_slave.r_user     ),
        .axi_slave_r_ready_i    ( axi_slave.r_ready    ),
        .axi_slave_b_valid_o    ( axi_slave.b_valid    ),
        .axi_slave_b_resp_o     ( axi_slave.b_resp     ),
        .axi_slave_b_id_o       ( axi_slave.b_id       ),
        .axi_slave_b_user_o     ( axi_slave.b_user     ),
        .axi_slave_b_ready_i    ( axi_slave.b_ready    ),
        .axi_master_aw_valid_o  ( axi_master.aw_valid  ),
        .axi_master_aw_addr_o   ( axi_master.aw_addr   ),
        .axi_master_aw_prot_o   ( axi_master.aw_prot   ),
        .axi_master_aw_region_o ( axi_master.aw_region ),
        .axi_master_aw_len_o    ( axi_master.aw_len    ),
        .axi_master_aw_size_o   ( axi_master.aw_size   ),
        .axi_master_aw_burst_o  ( axi_master.aw_burst  ),
        .axi_master_aw_lock_o   ( axi_master.aw_lock   ),
        .axi_master_aw_cache_o  ( axi_master.aw_cache  ),
        .axi_master_aw_qos_o    ( axi_master.aw_qos    ),
        .axi_master_aw_id_o     ( axi_master.aw_id     ),
        .axi_master_aw_user_o   ( axi_master.aw_user   ),
        .axi_master_aw_ready_i  ( axi_master.aw_ready  ),
        .axi_master_ar_valid_o  ( axi_master.ar_valid  ),
        .axi_master_ar_addr_o   ( axi_master.ar_addr   ),
        .axi_master_ar_prot_o   ( axi_master.ar_prot   ),
        .axi_master_ar_region_o ( axi_master.ar_region ),
        .axi_master_ar_len_o    ( axi_master.ar_len    ),
        .axi_master_ar_size_o   ( axi_master.ar_size   ),
        .axi_master_ar_burst_o  ( axi_master.ar_burst  ),
        .axi_master_ar_lock_o   ( axi_master.ar_lock   ),
        .axi_master_ar_cache_o  ( axi_master.ar_cache  ),
        .axi_master_ar_qos_o    ( axi_master.ar_qos    ),
        .axi_master_ar_id_o     ( axi_master.ar_id     ),
        .axi_master_ar_user_o   ( axi_master.ar_user   ),
        .axi_master_ar_ready_i  ( axi_master.ar_ready  ),
        .axi_master_w_valid_o   ( axi_master.w_valid   ),
        .axi_master_w_data_o    ( axi_master.w_data    ),
        .axi_master_w_strb_o    ( axi_master.w_strb    ),
        .axi_master_w_user_o    ( axi_master.w_user    ),
        .axi_master_w_last_o    ( axi_master.w_last    ),
        .axi_master_w_ready_i   ( axi_master.w_ready   ),
        .axi_master_r_valid_i   ( axi_master.r_valid   ),
        .axi_master_r_data_i    ( axi_master.r_data    ),
        .axi_master_r_resp_i    ( axi_master.r_resp    ),
        .axi_master_r_last_i    ( axi_master.r_last    ),
        .axi_master_r_id_i      ( axi_master.r_id      ),
        .axi_master_r_user_i    ( axi_master.r_user    ),
        .axi_master_r_ready_o   ( axi_master.r_ready   ),
        .axi_master_b_valid_i   ( axi_master.b_valid   ),
        .axi_master_b_resp_i    ( axi_master.b_resp    ),
        .axi_master_b_id_i      ( axi_master.b_id      ),
        .axi_master_b_user_i    ( axi_master.b_user    ),
        .axi_master_b_ready_o   ( axi_master.b_ready   ),
        .*
    );
endmodule
module axi_slice
#(
    parameter AXI_ADDR_WIDTH = 32,
    parameter AXI_DATA_WIDTH = 64,
    parameter AXI_USER_WIDTH = 6,
    parameter AXI_ID_WIDTH   = 3,
    parameter SLICE_DEPTH    = 2,
    parameter AXI_STRB_WIDTH = AXI_DATA_WIDTH/8
)
(
    input  logic                      clk_i,
    input  logic                      rst_ni,
    input  logic                      test_en_i,
    
    
    
    input  logic                      axi_slave_aw_valid_i,
    input  logic [AXI_ADDR_WIDTH-1:0] axi_slave_aw_addr_i,
    input  logic [2:0]                axi_slave_aw_prot_i,
    input  logic [3:0]                axi_slave_aw_region_i,
    input  logic [7:0]                axi_slave_aw_len_i,
    input  logic [2:0]                axi_slave_aw_size_i,
    input  logic [1:0]                axi_slave_aw_burst_i,
    input  logic                      axi_slave_aw_lock_i,
    input  logic [3:0]                axi_slave_aw_cache_i,
    input  logic [3:0]                axi_slave_aw_qos_i,
    input  logic [AXI_ID_WIDTH-1:0]   axi_slave_aw_id_i,
    input  logic [AXI_USER_WIDTH-1:0] axi_slave_aw_user_i,
    output logic                      axi_slave_aw_ready_o,
    
    input  logic                      axi_slave_ar_valid_i,
    input  logic [AXI_ADDR_WIDTH-1:0] axi_slave_ar_addr_i,
    input  logic [2:0]                axi_slave_ar_prot_i,
    input  logic [3:0]                axi_slave_ar_region_i,
    input  logic [7:0]                axi_slave_ar_len_i,
    input  logic [2:0]                axi_slave_ar_size_i,
    input  logic [1:0]                axi_slave_ar_burst_i,
    input  logic                      axi_slave_ar_lock_i,
    input  logic [3:0]                axi_slave_ar_cache_i,
    input  logic [3:0]                axi_slave_ar_qos_i,
    input  logic [AXI_ID_WIDTH-1:0]   axi_slave_ar_id_i,
    input  logic [AXI_USER_WIDTH-1:0] axi_slave_ar_user_i,
    output logic                      axi_slave_ar_ready_o,
    
    input  logic                      axi_slave_w_valid_i,
    input  logic [AXI_DATA_WIDTH-1:0] axi_slave_w_data_i,
    input  logic [AXI_STRB_WIDTH-1:0] axi_slave_w_strb_i,
    input  logic [AXI_USER_WIDTH-1:0] axi_slave_w_user_i,
    input  logic                      axi_slave_w_last_i,
    output logic                      axi_slave_w_ready_o,
    
    output logic                      axi_slave_r_valid_o,
    output logic [AXI_DATA_WIDTH-1:0] axi_slave_r_data_o,
    output logic [1:0]                axi_slave_r_resp_o,
    output logic                      axi_slave_r_last_o,
    output logic [AXI_ID_WIDTH-1:0]   axi_slave_r_id_o,
    output logic [AXI_USER_WIDTH-1:0] axi_slave_r_user_o,
    input  logic                      axi_slave_r_ready_i,
    
    output logic                      axi_slave_b_valid_o,
    output logic [1:0]                axi_slave_b_resp_o,
    output logic [AXI_ID_WIDTH-1:0]   axi_slave_b_id_o,
    output logic [AXI_USER_WIDTH-1:0] axi_slave_b_user_o,
    input  logic                      axi_slave_b_ready_i,
        
    
    
    output logic                      axi_master_aw_valid_o,
    output logic [AXI_ADDR_WIDTH-1:0] axi_master_aw_addr_o,
    output logic [2:0]                axi_master_aw_prot_o,
    output logic [3:0]                axi_master_aw_region_o,
    output logic [7:0]                axi_master_aw_len_o,
    output logic [2:0]                axi_master_aw_size_o,
    output logic [1:0]                axi_master_aw_burst_o,
    output logic                      axi_master_aw_lock_o,
    output logic [3:0]                axi_master_aw_cache_o,
    output logic [3:0]                axi_master_aw_qos_o,
    output logic [AXI_ID_WIDTH-1:0]   axi_master_aw_id_o,
    output logic [AXI_USER_WIDTH-1:0] axi_master_aw_user_o,
    input  logic                      axi_master_aw_ready_i,
    
    output logic                      axi_master_ar_valid_o,
    output logic [AXI_ADDR_WIDTH-1:0] axi_master_ar_addr_o,
    output logic [2:0]                axi_master_ar_prot_o,
    output logic [3:0]                axi_master_ar_region_o,
    output logic [7:0]                axi_master_ar_len_o,
    output logic [2:0]                axi_master_ar_size_o,
    output logic [1:0]                axi_master_ar_burst_o,
    output logic                      axi_master_ar_lock_o,
    output logic [3:0]                axi_master_ar_cache_o,
    output logic [3:0]                axi_master_ar_qos_o,
    output logic [AXI_ID_WIDTH-1:0]   axi_master_ar_id_o,
    output logic [AXI_USER_WIDTH-1:0] axi_master_ar_user_o,
    input  logic                      axi_master_ar_ready_i,
    
    output logic                      axi_master_w_valid_o,
    output logic [AXI_DATA_WIDTH-1:0] axi_master_w_data_o,
    output logic [AXI_STRB_WIDTH-1:0] axi_master_w_strb_o,
    output logic [AXI_USER_WIDTH-1:0] axi_master_w_user_o,
    output logic                      axi_master_w_last_o,
    input  logic                      axi_master_w_ready_i,
    
    input  logic                      axi_master_r_valid_i,
    input  logic [AXI_DATA_WIDTH-1:0] axi_master_r_data_i,
    input  logic [1:0]                axi_master_r_resp_i,
    input  logic                      axi_master_r_last_i,
    input  logic [AXI_ID_WIDTH-1:0]   axi_master_r_id_i,
    input  logic [AXI_USER_WIDTH-1:0] axi_master_r_user_i,
    output logic                      axi_master_r_ready_o,
    
    input  logic                      axi_master_b_valid_i,
    input  logic [1:0]                axi_master_b_resp_i,
    input  logic [AXI_ID_WIDTH-1:0]   axi_master_b_id_i,
    input  logic [AXI_USER_WIDTH-1:0] axi_master_b_user_i,
    output logic                      axi_master_b_ready_o
);
   
   axi_aw_buffer
   #(
       .ID_WIDTH     (AXI_ID_WIDTH),
       .ADDR_WIDTH   (AXI_ADDR_WIDTH),
       .USER_WIDTH   (AXI_USER_WIDTH),
       .BUFFER_DEPTH (SLICE_DEPTH)
   )
   aw_buffer_i
   (
      .clk_i            ( clk_i                  ),
      .rst_ni           ( rst_ni                 ),
      .test_en_i        ( test_en_i              ),
      .slave_valid_i    ( axi_slave_aw_valid_i   ),
      .slave_addr_i     ( axi_slave_aw_addr_i    ),
      .slave_prot_i     ( axi_slave_aw_prot_i    ),
      .slave_region_i   ( axi_slave_aw_region_i  ),
      .slave_len_i      ( axi_slave_aw_len_i     ),
      .slave_size_i     ( axi_slave_aw_size_i    ),
      .slave_burst_i    ( axi_slave_aw_burst_i   ),
      .slave_lock_i     ( axi_slave_aw_lock_i    ),
      .slave_cache_i    ( axi_slave_aw_cache_i   ),
      .slave_qos_i      ( axi_slave_aw_qos_i     ),
      .slave_id_i       ( axi_slave_aw_id_i      ),
      .slave_user_i     ( axi_slave_aw_user_i    ),
      .slave_ready_o    ( axi_slave_aw_ready_o   ),
      .master_valid_o   ( axi_master_aw_valid_o  ),
      .master_addr_o    ( axi_master_aw_addr_o   ),
      .master_prot_o    ( axi_master_aw_prot_o   ),
      .master_region_o  ( axi_master_aw_region_o ),
      .master_len_o     ( axi_master_aw_len_o    ),
      .master_size_o    ( axi_master_aw_size_o   ),
      .master_burst_o   ( axi_master_aw_burst_o  ),
      .master_lock_o    ( axi_master_aw_lock_o   ),
      .master_cache_o   ( axi_master_aw_cache_o  ),
      .master_qos_o     ( axi_master_aw_qos_o    ),
      .master_id_o      ( axi_master_aw_id_o     ),
      .master_user_o    ( axi_master_aw_user_o   ),
      .master_ready_i   ( axi_master_aw_ready_i  )
   );
   
   axi_ar_buffer
   #(
       .ID_WIDTH     (AXI_ID_WIDTH),
       .ADDR_WIDTH   (AXI_ADDR_WIDTH),
       .USER_WIDTH   (AXI_USER_WIDTH),
       .BUFFER_DEPTH (SLICE_DEPTH)
   )
   ar_buffer_i
   (
      .clk_i           ( clk_i                   ),
      .rst_ni          ( rst_ni                  ),
      .test_en_i       ( test_en_i               ),
      .slave_valid_i   ( axi_slave_ar_valid_i    ),
      .slave_addr_i    ( axi_slave_ar_addr_i     ),
      .slave_prot_i    ( axi_slave_ar_prot_i     ),
      .slave_region_i  ( axi_slave_ar_region_i   ),
      .slave_len_i     ( axi_slave_ar_len_i      ),
      .slave_size_i    ( axi_slave_ar_size_i     ),
      .slave_burst_i   ( axi_slave_ar_burst_i    ),
      .slave_lock_i    ( axi_slave_ar_lock_i     ),
      .slave_cache_i   ( axi_slave_ar_cache_i    ),
      .slave_qos_i     ( axi_slave_ar_qos_i      ),
      .slave_id_i      ( axi_slave_ar_id_i       ),
      .slave_user_i    ( axi_slave_ar_user_i     ),
      .slave_ready_o   ( axi_slave_ar_ready_o    ),
      .master_valid_o  ( axi_master_ar_valid_o   ),
      .master_addr_o   ( axi_master_ar_addr_o    ),
      .master_prot_o   ( axi_master_ar_prot_o    ),
      .master_region_o ( axi_master_ar_region_o  ),
      .master_len_o    ( axi_master_ar_len_o     ),
      .master_size_o   ( axi_master_ar_size_o    ),
      .master_burst_o  ( axi_master_ar_burst_o   ),
      .master_lock_o   ( axi_master_ar_lock_o    ),
      .master_cache_o  ( axi_master_ar_cache_o   ),
      .master_qos_o    ( axi_master_ar_qos_o     ),
      .master_id_o     ( axi_master_ar_id_o      ),
      .master_user_o   ( axi_master_ar_user_o    ),
      .master_ready_i  ( axi_master_ar_ready_i   )
   );
   
   axi_w_buffer
   #(
       .DATA_WIDTH   (AXI_DATA_WIDTH),
       .USER_WIDTH   (AXI_USER_WIDTH),
       .BUFFER_DEPTH (SLICE_DEPTH)
   )
   w_buffer_i
   (
      .clk_i          ( clk_i                 ),
      .rst_ni         ( rst_ni                ),
      .test_en_i      ( test_en_i             ),
      .slave_valid_i  ( axi_slave_w_valid_i   ),
      .slave_data_i   ( axi_slave_w_data_i    ),
      .slave_strb_i   ( axi_slave_w_strb_i    ),
      .slave_user_i   ( axi_slave_w_user_i    ),
      .slave_last_i   ( axi_slave_w_last_i    ),
      .slave_ready_o  ( axi_slave_w_ready_o   ),
      .master_valid_o ( axi_master_w_valid_o  ),
      .master_data_o  ( axi_master_w_data_o   ),
      .master_strb_o  ( axi_master_w_strb_o   ),
      .master_user_o  ( axi_master_w_user_o   ),
      .master_last_o  ( axi_master_w_last_o   ),
      .master_ready_i ( axi_master_w_ready_i  )
   );
   
   axi_r_buffer
   #(
       .ID_WIDTH     (AXI_ID_WIDTH),
       .DATA_WIDTH   (AXI_DATA_WIDTH),
       .USER_WIDTH   (AXI_USER_WIDTH),
       .BUFFER_DEPTH (SLICE_DEPTH)
   )
   r_buffer_i
   (
      .clk_i           ( clk_i                 ),
      .rst_ni          ( rst_ni                ),
      .test_en_i       ( test_en_i             ),
      .slave_valid_i   ( axi_master_r_valid_i  ),
      .slave_data_i    ( axi_master_r_data_i   ),
      .slave_resp_i    ( axi_master_r_resp_i   ),
      .slave_user_i    ( axi_master_r_user_i   ),
      .slave_id_i      ( axi_master_r_id_i     ),
      .slave_last_i    ( axi_master_r_last_i   ),
      .slave_ready_o   ( axi_master_r_ready_o  ),
      .master_valid_o  ( axi_slave_r_valid_o   ),
      .master_data_o   ( axi_slave_r_data_o    ),
      .master_resp_o   ( axi_slave_r_resp_o    ),
      .master_user_o   ( axi_slave_r_user_o    ),
      .master_id_o     ( axi_slave_r_id_o      ),
      .master_last_o   ( axi_slave_r_last_o    ),
      .master_ready_i  ( axi_slave_r_ready_i   )
   );
   
   axi_b_buffer
   #(
       .ID_WIDTH     (AXI_ID_WIDTH),
       .USER_WIDTH   (AXI_USER_WIDTH),
       .BUFFER_DEPTH (SLICE_DEPTH)
   )
   b_buffer_i
   (
      .clk_i           ( clk_i                 ),
      .rst_ni          ( rst_ni                ),
      .test_en_i       ( test_en_i             ),
      .slave_valid_i   ( axi_master_b_valid_i  ),
      .slave_resp_i    ( axi_master_b_resp_i   ),
      .slave_id_i      ( axi_master_b_id_i     ),
      .slave_user_i    ( axi_master_b_user_i   ),
      .slave_ready_o   ( axi_master_b_ready_o  ),
      .master_valid_o  ( axi_slave_b_valid_o   ),
      .master_resp_o   ( axi_slave_b_resp_o    ),
      .master_id_o     ( axi_slave_b_id_o      ),
      .master_user_o   ( axi_slave_b_user_o    ),
      .master_ready_i  ( axi_slave_b_ready_i   )
   );
endmodule
module axi_single_slice #(
    parameter int BUFFER_DEPTH = -1,
    parameter int DATA_WIDTH   = -1
) (
    input  logic                  clk_i,    
    input  logic                  rst_ni,  
    input  logic                  testmode_i,
    input  logic                  valid_i,
    output logic                  ready_o,
    input  logic [DATA_WIDTH-1:0] data_i,
    input  logic                  ready_i,
    output logic                  valid_o,
    output logic [DATA_WIDTH-1:0] data_o
);
    logic full, empty;
    assign ready_o = ~full;
    assign valid_o = ~empty;
    fifo #(
        .FALL_THROUGH ( 1'b0         ),
        .DATA_WIDTH   ( DATA_WIDTH   ),
        .DEPTH        ( BUFFER_DEPTH )
    ) i_fifo (
        .clk_i      ( clk_i             ),
        .rst_ni     ( rst_ni            ),
        .flush_i    ( 1'b0              ),
        .threshold_o (), 
        .testmode_i ( testmode_i        ),
        .full_o     ( full              ),
        .empty_o    ( empty             ),
        .data_i     ( data_i            ),
        .push_i     ( valid_i & ready_o ),
        .data_o     ( data_o            ),
        .pop_i      ( ready_i & valid_o )
    );
endmodule
module axi_ar_buffer #(
    parameter int ID_WIDTH     = -1,
    parameter int ADDR_WIDTH   = -1,
    parameter int USER_WIDTH   = -1,
    parameter int BUFFER_DEPTH = -1
)(
    input logic                   clk_i,
    input logic                   rst_ni,
    input logic                   test_en_i,
    input  logic                  slave_valid_i,
    input  logic [ADDR_WIDTH-1:0] slave_addr_i,
    input  logic [2:0]            slave_prot_i,
    input  logic [3:0]            slave_region_i,
    input  logic [7:0]            slave_len_i,
    input  logic [2:0]            slave_size_i,
    input  logic [1:0]            slave_burst_i,
    input  logic                  slave_lock_i,
    input  logic [3:0]            slave_cache_i,
    input  logic [3:0]            slave_qos_i,
    input  logic [ID_WIDTH-1:0]   slave_id_i,
    input  logic [USER_WIDTH-1:0] slave_user_i,
    output logic                  slave_ready_o,
    output logic                  master_valid_o,
    output logic [ADDR_WIDTH-1:0] master_addr_o,
    output logic [2:0]            master_prot_o,
    output logic [3:0]            master_region_o,
    output logic [7:0]            master_len_o,
    output logic [2:0]            master_size_o,
    output logic [1:0]            master_burst_o,
    output logic                  master_lock_o,
    output logic [3:0]            master_cache_o,
    output logic [3:0]            master_qos_o,
    output logic [ID_WIDTH-1:0]   master_id_o,
    output logic [USER_WIDTH-1:0] master_user_o,
    input  logic                  master_ready_i
);
   logic [29+ADDR_WIDTH+USER_WIDTH+ID_WIDTH-1:0] s_data_in;
   logic [29+ADDR_WIDTH+USER_WIDTH+ID_WIDTH-1:0] s_data_out;
   assign s_data_in = {slave_cache_i,  slave_prot_i,  slave_lock_i,  slave_burst_i,  slave_size_i,  slave_len_i,  slave_qos_i,  slave_region_i,  slave_addr_i,  slave_user_i,  slave_id_i} ;
   assign             {master_cache_o, master_prot_o, master_lock_o, master_burst_o, master_size_o, master_len_o, master_qos_o, master_region_o, master_addr_o, master_user_o, master_id_o} =  s_data_out;
  axi_single_slice #(.BUFFER_DEPTH(BUFFER_DEPTH), .DATA_WIDTH(29+ADDR_WIDTH+USER_WIDTH+ID_WIDTH)) i_axi_single_slice (
    .clk_i      ( clk_i          ),
    .rst_ni     ( rst_ni         ),
    .testmode_i ( test_en_i      ),
    .valid_i    ( slave_valid_i  ),
    .ready_o    ( slave_ready_o  ),
    .data_i     ( s_data_in      ),
    .ready_i    ( master_ready_i ),
    .valid_o    ( master_valid_o ),
    .data_o     ( s_data_out     )
  );
endmodule
module axi_r_buffer #(
   parameter ID_WIDTH      = 4,
   parameter DATA_WIDTH    = 64,
   parameter USER_WIDTH    = 6,
   parameter BUFFER_DEPTH  = 8,
   parameter STRB_WIDTH    = DATA_WIDTH/8   
)(
   input logic                   clk_i,
   input logic                   rst_ni,
   input logic                   test_en_i,
   input logic                   slave_valid_i,
   input logic  [DATA_WIDTH-1:0] slave_data_i,
   input logic  [1:0]            slave_resp_i,
   input logic  [USER_WIDTH-1:0] slave_user_i,
   input logic  [ID_WIDTH-1:0]   slave_id_i,
   input logic                   slave_last_i,
   output logic                  slave_ready_o,
   output logic                  master_valid_o,
   output logic [DATA_WIDTH-1:0] master_data_o,
   output logic [1:0]            master_resp_o,
   output logic [USER_WIDTH-1:0] master_user_o,
   output logic [ID_WIDTH-1:0]   master_id_o,
   output logic                  master_last_o,
   input  logic                  master_ready_i
);
   logic [2+DATA_WIDTH+USER_WIDTH+ID_WIDTH:0] s_data_in;
   logic [2+DATA_WIDTH+USER_WIDTH+ID_WIDTH:0] s_data_out;
   assign s_data_in =  {slave_id_i,  slave_user_i,  slave_data_i,  slave_resp_i,  slave_last_i};
   assign              {master_id_o, master_user_o, master_data_o, master_resp_o, master_last_o} = s_data_out;
   axi_single_slice #(.BUFFER_DEPTH(BUFFER_DEPTH), .DATA_WIDTH(3+DATA_WIDTH+USER_WIDTH+ID_WIDTH)) i_axi_single_slice (
     .clk_i      ( clk_i          ),
     .rst_ni     ( rst_ni         ),
     .testmode_i ( test_en_i      ),
     .valid_i    ( slave_valid_i  ),
     .ready_o    ( slave_ready_o  ),
     .data_i     ( s_data_in      ),
     .ready_i    ( master_ready_i ),
     .valid_o    ( master_valid_o ),
     .data_o     ( s_data_out     )
   );
endmodule
module axi_aw_buffer #(
    parameter int ID_WIDTH     = -1,
    parameter int ADDR_WIDTH   = -1,
    parameter int USER_WIDTH   = -1,
    parameter int BUFFER_DEPTH = -1
)(
    input logic                   clk_i,
    input logic                   rst_ni,
    input logic                   test_en_i,
    input  logic                  slave_valid_i,
    input  logic [ADDR_WIDTH-1:0] slave_addr_i,
    input  logic [2:0]            slave_prot_i,
    input  logic [3:0]            slave_region_i,
    input  logic [7:0]            slave_len_i,
    input  logic [2:0]            slave_size_i,
    input  logic [1:0]            slave_burst_i,
    input  logic                  slave_lock_i,
    input  logic [3:0]            slave_cache_i,
    input  logic [3:0]            slave_qos_i,
    input  logic [ID_WIDTH-1:0]   slave_id_i,
    input  logic [USER_WIDTH-1:0] slave_user_i,
    output logic                  slave_ready_o,
    output logic                  master_valid_o,
    output logic [ADDR_WIDTH-1:0] master_addr_o,
    output logic [2:0]            master_prot_o,
    output logic [3:0]            master_region_o,
    output logic [7:0]            master_len_o,
    output logic [2:0]            master_size_o,
    output logic [1:0]            master_burst_o,
    output logic                  master_lock_o,
    output logic [3:0]            master_cache_o,
    output logic [3:0]            master_qos_o,
    output logic [ID_WIDTH-1:0]   master_id_o,
    output logic [USER_WIDTH-1:0] master_user_o,
    input  logic                  master_ready_i
);
   logic [29+ADDR_WIDTH+USER_WIDTH+ID_WIDTH-1:0] s_data_in;
   logic [29+ADDR_WIDTH+USER_WIDTH+ID_WIDTH-1:0] s_data_out;
   assign s_data_in = {slave_cache_i,  slave_prot_i,  slave_lock_i,  slave_burst_i,  slave_size_i,  slave_len_i,  slave_qos_i,  slave_region_i,  slave_addr_i,  slave_user_i,  slave_id_i};
   assign             {master_cache_o, master_prot_o, master_lock_o, master_burst_o, master_size_o, master_len_o, master_qos_o, master_region_o, master_addr_o, master_user_o, master_id_o} = s_data_out;
    axi_single_slice #(.BUFFER_DEPTH(BUFFER_DEPTH), .DATA_WIDTH(29+ADDR_WIDTH+USER_WIDTH+ID_WIDTH)) i_axi_single_slice (
      .clk_i      ( clk_i          ),
      .rst_ni     ( rst_ni         ),
      .testmode_i ( test_en_i      ),
      .valid_i    ( slave_valid_i  ),
      .ready_o    ( slave_ready_o  ),
      .data_i     ( s_data_in      ),
      .ready_i    ( master_ready_i ),
      .valid_o    ( master_valid_o ),
      .data_o     ( s_data_out     )
    );
endmodule
module ariane_verilog_wrap
    import ariane_pkg::*;
#(
  parameter int unsigned               RASDepth              = 2,
  parameter int unsigned               BTBEntries            = 32,
  parameter int unsigned               BHTEntries            = 128,
  
  parameter logic [63:0]               DmBaseAddress         = 64'h0,
  
  parameter bit                        SwapEndianess         = 1,
  
  
  parameter int unsigned               NrNonIdempotentRules  =  1,
  parameter logic [NrMaxRules*64-1:0]  NonIdempotentAddrBase = 64'h00C0000000,
  parameter logic [NrMaxRules*64-1:0]  NonIdempotentLength   = 64'hFFFFFFFFFF,
  
  parameter int unsigned               NrExecuteRegionRules  =  0,
  parameter logic [NrMaxRules*64-1:0]  ExecuteRegionAddrBase = '0,
  parameter logic [NrMaxRules*64-1:0]  ExecuteRegionLength   = '0,
  
  parameter int unsigned               NrCachedRegionRules   =  0,
  parameter logic [NrMaxRules*64-1:0]  CachedRegionAddrBase  = '0,
  parameter logic [NrMaxRules*64-1:0]  CachedRegionLength    = '0,
  
  parameter int unsigned               NrPMPEntries          =  8
) (
  input                       clk_i,
  input                       reset_l,      
  output                      spc_grst_l,   
  
  input  [riscv::VLEN-1:0]               boot_addr_i,  
  input  [riscv::XLEN-1:0]               hart_id_i,    
  
  input  [1:0]                irq_i,        
  input                       ipi_i,        
  
  input                       time_irq_i,   
  input                       debug_req_i,  
  
  output [$size(wt_cache_pkg::l15_req_t)-1:0]  l15_req_o,
  input  [$size(wt_cache_pkg::l15_rtrn_t)-1:0] l15_rtrn_i
 );
  
  wt_cache_pkg::l15_req_t  l15_req;
  wt_cache_pkg::l15_rtrn_t l15_rtrn;
  assign l15_req_o = l15_req;
  assign l15_rtrn  = l15_rtrn_i;
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  logic [15:0] wake_up_cnt_d, wake_up_cnt_q;
  logic rst_n;
  assign wake_up_cnt_d = (wake_up_cnt_q[$high(wake_up_cnt_q)]) ? wake_up_cnt_q : wake_up_cnt_q + 1;
  always_ff @(posedge clk_i or negedge reset_l) begin : p_regs
    if(~reset_l) begin
      wake_up_cnt_q <= 0;
    end else begin
      wake_up_cnt_q <= wake_up_cnt_d;
    end
  end
  
  assign rst_n = wake_up_cnt_q[$high(wake_up_cnt_q)] & reset_l;
  
  
  
  logic [1:0] irq;
  logic ipi, time_irq, debug_req;
  
  synchronizer i_sync (
    .clk         ( clk_i      ),
    .presyncdata ( rst_n      ),
    .syncdata    ( spc_grst_l )
  );
  
  for (genvar k=0; k<$size(irq_i); k++) begin
    synchronizer i_irq_sync (
      .clk         ( clk_i      ),
      .presyncdata ( irq_i[k]   ),
      .syncdata    ( irq[k]     )
    );
  end
  synchronizer i_ipi_sync (
    .clk         ( clk_i      ),
    .presyncdata ( ipi_i      ),
    .syncdata    ( ipi        )
  );
  synchronizer i_timer_sync (
    .clk         ( clk_i      ),
    .presyncdata ( time_irq_i ),
    .syncdata    ( time_irq   )
  );
  synchronizer i_debug_sync (
    .clk         ( clk_i       ),
    .presyncdata ( debug_req_i ),
    .syncdata    ( debug_req   )
  );
  
  
  
  localparam ariane_pkg::ariane_cfg_t ArianeOpenPitonCfg = '{
    RASDepth:              RASDepth,
    BTBEntries:            BTBEntries,
    BHTEntries:            BHTEntries,
    
    NrNonIdempotentRules:  NrNonIdempotentRules,
    NonIdempotentAddrBase: NonIdempotentAddrBase,
    NonIdempotentLength:   NonIdempotentLength,
    NrExecuteRegionRules:  NrExecuteRegionRules,
    ExecuteRegionAddrBase: ExecuteRegionAddrBase,
    ExecuteRegionLength:   ExecuteRegionLength,
    
    NrCachedRegionRules:   NrCachedRegionRules,
    CachedRegionAddrBase:  CachedRegionAddrBase,
    CachedRegionLength:    CachedRegionLength,
    
    Axi64BitCompliant:     1'b0,
    SwapEndianess:         SwapEndianess,
    
    DmBaseAddress:         DmBaseAddress,
    NrPMPEntries:          NrPMPEntries
  };
  ariane #(
    .ArianeCfg ( ArianeOpenPitonCfg )
  ) ariane (
    .clk_i       ( clk_i      ),
    .rst_ni      ( spc_grst_l ),
    .boot_addr_i              ,
    .hart_id_i                ,
    .irq_i       ( irq        ),
    .ipi_i       ( ipi        ),
    .time_irq_i  ( time_irq   ),
    .debug_req_i ( debug_req  ),
    .l15_req_o   ( l15_req   ),
    .l15_rtrn_i  ( l15_rtrn  )
  );
endmodule 
module riscv_peripherals #(
    parameter int unsigned DataWidth       = 64,
    parameter int unsigned NumHarts        =  1,
    parameter int unsigned NumSources      =  1,
    parameter int unsigned PlicMaxPriority =  7,
    parameter bit          SwapEndianess   =  0,
    parameter logic [63:0] DmBase          = 64'hfff1000000,
    parameter logic [63:0] RomBase         = 64'hfff1010000,
    parameter logic [63:0] ClintBase       = 64'hfff1020000,
    parameter logic [63:0] PlicBase        = 64'hfff1100000
) (
    input                               clk_i,
    input                               rst_ni,
    input                               testmode_i,
    
    
    input  [DataWidth-1:0]              buf_ariane_debug_noc2_data_i,
    input                               buf_ariane_debug_noc2_valid_i,
    output                              ariane_debug_buf_noc2_ready_o,
    output [DataWidth-1:0]              ariane_debug_buf_noc3_data_o,
    output                              ariane_debug_buf_noc3_valid_o,
    input                               buf_ariane_debug_noc3_ready_i,
    
    input  [DataWidth-1:0]              buf_ariane_bootrom_noc2_data_i,
    input                               buf_ariane_bootrom_noc2_valid_i,
    output                              ariane_bootrom_buf_noc2_ready_o,
    output [DataWidth-1:0]              ariane_bootrom_buf_noc3_data_o,
    output                              ariane_bootrom_buf_noc3_valid_o,
    input                               buf_ariane_bootrom_noc3_ready_i,
    
    input  [DataWidth-1:0]              buf_ariane_clint_noc2_data_i,
    input                               buf_ariane_clint_noc2_valid_i,
    output                              ariane_clint_buf_noc2_ready_o,
    output [DataWidth-1:0]              ariane_clint_buf_noc3_data_o,
    output                              ariane_clint_buf_noc3_valid_o,
    input                               buf_ariane_clint_noc3_ready_i,
    
    input [DataWidth-1:0]               buf_ariane_plic_noc2_data_i,
    input                               buf_ariane_plic_noc2_valid_i,
    output                              ariane_plic_buf_noc2_ready_o,
    output [DataWidth-1:0]              ariane_plic_buf_noc3_data_o,
    output                              ariane_plic_buf_noc3_valid_o,
    input                               buf_ariane_plic_noc3_ready_i,
    
    input                               ariane_boot_sel_i,
    
    output                              ndmreset_o,    
    output                              dmactive_o,    
    output [NumHarts-1:0]               debug_req_o,   
    input  [NumHarts-1:0]               unavailable_i, 
    
    input                               tck_i,
    input                               tms_i,
    input                               trst_ni,
    input                               td_i,
    output                              td_o,
    output                              tdo_oe_o,
    
    input                               rtc_i,        
    output [NumHarts-1:0]               timer_irq_o,  
    output [NumHarts-1:0]               ipi_o,        
    
    input  [NumSources-1:0]             irq_sources_i,
    input  [NumSources-1:0]             irq_le_i,     
    output [NumHarts-1:0][1:0]          irq_o         
);
  localparam int unsigned AxiIdWidth    =  1;
  localparam int unsigned AxiAddrWidth  = 64;
  localparam int unsigned AxiDataWidth  = 64;
  localparam int unsigned AxiUserWidth  =  1;
  
  
  
  logic          debug_req_valid;
  logic          debug_req_ready;
  logic          debug_resp_valid;
  logic          debug_resp_ready;
  dm::dmi_req_t  debug_req;
  dm::dmi_resp_t debug_resp;
 
  logic        tck, tms, trst_n, tdi, tdo, tdo_oe;
  dmi_jtag i_dmi_jtag (
    .clk_i                                ,
    .rst_ni                               ,
    .testmode_i                           ,
    .dmi_req_o        ( debug_req        ),
    .dmi_req_valid_o  ( debug_req_valid  ),
    .dmi_req_ready_i  ( debug_req_ready  ),
    .dmi_resp_i       ( debug_resp       ),
    .dmi_resp_ready_o ( debug_resp_ready ),
    .dmi_resp_valid_i ( debug_resp_valid ),
    .dmi_rst_no       (                  ), 
    .tck_i            ( tck              ),
    .tms_i            ( tms              ),
    .trst_ni          ( trst_n           ),
    .td_i             ( tdi              ),
    .td_o             ( tdo              ),
    .tdo_oe_o         ( tdo_oe           )
  );
 
  assign tck      = tck_i   ;
  assign tms      = tms_i   ;
  assign trst_n   = trst_ni ;
  assign tdi      = td_i    ;
  assign td_o     = tdo     ;
  assign tdo_oe_o = tdo_oe  ;
 
 
  logic                dm_slave_req;
  logic                dm_slave_we;
  logic [64-1:0]       dm_slave_addr;
  logic [64/8-1:0]     dm_slave_be;
  logic [64-1:0]       dm_slave_wdata;
  logic [64-1:0]       dm_slave_rdata;
  logic                dm_master_req;
  logic [64-1:0]       dm_master_add;
  logic                dm_master_we;
  logic [64-1:0]       dm_master_wdata;
  logic [64/8-1:0]     dm_master_be;
  logic                dm_master_gnt;
  logic                dm_master_r_valid;
  logic [64-1:0]       dm_master_r_rdata;
  
  dm_top #(
    .NrHarts              ( NumHarts             ),
    .BusWidth             ( AxiDataWidth         ),
    .SelectableHarts      ( {NumHarts{1'b1}}     )
  ) i_dm_top (
    .clk_i                                        ,
    .rst_ni                                       , 
    .testmode_i                                   ,
    .ndmreset_o                                   ,
    .dmactive_o                                   , 
    .debug_req_o                                  ,
    .unavailable_i                                ,
    .hartinfo_i           ( {NumHarts{ariane_pkg::DebugHartInfo}} ),
    .slave_req_i          ( dm_slave_req         ),
    .slave_we_i           ( dm_slave_we          ),
    .slave_addr_i         ( dm_slave_addr        ),
    .slave_be_i           ( dm_slave_be          ),
    .slave_wdata_i        ( dm_slave_wdata       ),
    .slave_rdata_o        ( dm_slave_rdata       ),
    .master_req_o         ( dm_master_req        ),
    .master_add_o         ( dm_master_add        ),
    .master_we_o          ( dm_master_we         ),
    .master_wdata_o       ( dm_master_wdata      ),
    .master_be_o          ( dm_master_be         ),
    .master_gnt_i         ( dm_master_gnt        ),
    .master_r_valid_i     ( dm_master_r_valid    ),
    .master_r_rdata_i     ( dm_master_r_rdata    ),
    .dmi_rst_ni           ( rst_ni               ),
    .dmi_req_valid_i      ( debug_req_valid      ),
    .dmi_req_ready_o      ( debug_req_ready      ),
    .dmi_req_i            ( debug_req            ),
    .dmi_resp_valid_o     ( debug_resp_valid     ),
    .dmi_resp_ready_i     ( debug_resp_ready     ),
    .dmi_resp_o           ( debug_resp           )
  );
  AXI_BUS #(
      .AXI_ADDR_WIDTH ( AxiAddrWidth     ),
      .AXI_DATA_WIDTH ( AxiDataWidth     ),
      .AXI_ID_WIDTH   ( AxiIdWidth       ),
      .AXI_USER_WIDTH ( AxiUserWidth     )
  ) dm_master();
  axi2mem #(
      .AXI_ID_WIDTH   ( AxiIdWidth   ),
      .AXI_ADDR_WIDTH ( AxiAddrWidth ),
      .AXI_DATA_WIDTH ( AxiDataWidth ),
      .AXI_USER_WIDTH ( AxiUserWidth )
  ) i_dm_axi2mem (
      .clk_i      ( clk_i                     ),
      .rst_ni     ( rst_ni                    ),
      .slave      ( dm_master                 ),
      .req_o      ( dm_slave_req              ),
      .we_o       ( dm_slave_we               ),
      .addr_o     ( dm_slave_addr             ),
      .be_o       ( dm_slave_be               ),
      .data_o     ( dm_slave_wdata            ),
      .data_i     ( dm_slave_rdata            )
  );
  noc_axilite_bridge #(
    .SLAVE_RESP_BYTEWIDTH   ( 8             ),
    .SWAP_ENDIANESS         ( SwapEndianess )
  ) i_debug_axilite_bridge (
    .clk                    ( clk_i                         ),
    .rst                    ( ~rst_ni                       ),
    
    .splitter_bridge_val    ( buf_ariane_debug_noc2_valid_i ),
    .splitter_bridge_data   ( buf_ariane_debug_noc2_data_i  ),
    .bridge_splitter_rdy    ( ariane_debug_buf_noc2_ready_o ),
    .bridge_splitter_val    ( ariane_debug_buf_noc3_valid_o ),
    .bridge_splitter_data   ( ariane_debug_buf_noc3_data_o  ),
    .splitter_bridge_rdy    ( buf_ariane_debug_noc3_ready_i ),
    
    
    .m_axi_awaddr           ( dm_master.aw_addr             ),
    .m_axi_awvalid          ( dm_master.aw_valid            ),
    .m_axi_awready          ( dm_master.aw_ready            ),
    
    .m_axi_wdata            ( dm_master.w_data              ),
    .m_axi_wstrb            ( dm_master.w_strb              ),
    .m_axi_wvalid           ( dm_master.w_valid             ),
    .m_axi_wready           ( dm_master.w_ready             ),
    
    .m_axi_araddr           ( dm_master.ar_addr             ),
    .m_axi_arvalid          ( dm_master.ar_valid            ),
    .m_axi_arready          ( dm_master.ar_ready            ),
    
    .m_axi_rdata            ( dm_master.r_data              ),
    .m_axi_rresp            ( dm_master.r_resp              ),
    .m_axi_rvalid           ( dm_master.r_valid             ),
    .m_axi_rready           ( dm_master.r_ready             ),
    
    .m_axi_bresp            ( dm_master.b_resp              ),
    .m_axi_bvalid           ( dm_master.b_valid             ),
    .m_axi_bready           ( dm_master.b_ready             ),
    
    .w_reqbuf_size          (                               ),
    .r_reqbuf_size          (                               )
  );
  
  
  assign dm_master_gnt      = '0;
  assign dm_master_r_valid  = '0;
  assign dm_master_r_rdata  = '0;
  
  assign dm_master.aw_id     = '0;
  assign dm_master.aw_len    = '0;
  assign dm_master.aw_size   = 3'b11;
  assign dm_master.aw_burst  = '0;
  assign dm_master.aw_lock   = '0;
  assign dm_master.aw_cache  = '0;
  assign dm_master.aw_prot   = '0;
  assign dm_master.aw_qos    = '0;
  assign dm_master.aw_region = '0;
  assign dm_master.aw_atop   = '0;
  assign dm_master.w_last    = 1'b1;
  assign dm_master.ar_id     = '0;
  assign dm_master.ar_len    = '0;
  assign dm_master.ar_size   = 3'b11;
  assign dm_master.ar_burst  = '0;
  assign dm_master.ar_lock   = '0;
  assign dm_master.ar_cache  = '0;
  assign dm_master.ar_prot   = '0;
  assign dm_master.ar_qos    = '0;
  assign dm_master.ar_region = '0;
  
  
  
  logic                    rom_req;
  logic [AxiAddrWidth-1:0] rom_addr;
  logic [AxiDataWidth-1:0] rom_rdata, rom_rdata_bm, rom_rdata_linux;
  AXI_BUS #(
    .AXI_ID_WIDTH   ( AxiIdWidth   ),
    .AXI_ADDR_WIDTH ( AxiAddrWidth ),
    .AXI_DATA_WIDTH ( AxiDataWidth ),
    .AXI_USER_WIDTH ( AxiUserWidth )
  ) br_master();
  axi2mem #(
    .AXI_ID_WIDTH   ( AxiIdWidth    ),
    .AXI_ADDR_WIDTH ( AxiAddrWidth  ),
    .AXI_DATA_WIDTH ( AxiDataWidth  ),
    .AXI_USER_WIDTH ( AxiUserWidth  )
  ) i_axi2rom (
    .clk_i                ,
    .rst_ni               ,
    .slave  ( br_master  ),
    .req_o  ( rom_req    ),
    .we_o   (            ),
    .addr_o ( rom_addr   ),
    .be_o   (            ),
    .data_o (            ),
    .data_i ( rom_rdata  )
  );
  bootrom i_bootrom_bm (
    .clk_i                   ,
    .req_i      ( rom_req   ),
    .addr_i     ( rom_addr  ),
    .rdata_o    ( rom_rdata_bm )
  );
  bootrom_linux i_bootrom_linux (
    .clk_i                   ,
    .req_i      ( rom_req   ),
    .addr_i     ( rom_addr  ),
    .rdata_o    ( rom_rdata_linux )
  );
  
  assign rom_rdata = (ariane_boot_sel_i) ? rom_rdata_bm : rom_rdata_linux;
  noc_axilite_bridge #(
    .SLAVE_RESP_BYTEWIDTH   ( 8             ),
    .SWAP_ENDIANESS         ( SwapEndianess )
  ) i_bootrom_axilite_bridge (
    .clk                    ( clk_i                           ),
    .rst                    ( ~rst_ni                         ),
    
    .splitter_bridge_val    ( buf_ariane_bootrom_noc2_valid_i ),
    .splitter_bridge_data   ( buf_ariane_bootrom_noc2_data_i  ),
    .bridge_splitter_rdy    ( ariane_bootrom_buf_noc2_ready_o ),
    .bridge_splitter_val    ( ariane_bootrom_buf_noc3_valid_o ),
    .bridge_splitter_data   ( ariane_bootrom_buf_noc3_data_o  ),
    .splitter_bridge_rdy    ( buf_ariane_bootrom_noc3_ready_i ),
    
    
    .m_axi_awaddr           ( br_master.aw_addr               ),
    .m_axi_awvalid          ( br_master.aw_valid              ),
    .m_axi_awready          ( br_master.aw_ready              ),
    
    .m_axi_wdata            ( br_master.w_data                ),
    .m_axi_wstrb            ( br_master.w_strb                ),
    .m_axi_wvalid           ( br_master.w_valid               ),
    .m_axi_wready           ( br_master.w_ready               ),
    
    .m_axi_araddr           ( br_master.ar_addr               ),
    .m_axi_arvalid          ( br_master.ar_valid              ),
    .m_axi_arready          ( br_master.ar_ready              ),
    
    .m_axi_rdata            ( br_master.r_data                ),
    .m_axi_rresp            ( br_master.r_resp                ),
    .m_axi_rvalid           ( br_master.r_valid               ),
    .m_axi_rready           ( br_master.r_ready               ),
    
    .m_axi_bresp            ( br_master.b_resp                ),
    .m_axi_bvalid           ( br_master.b_valid               ),
    .m_axi_bready           ( br_master.b_ready               ),
    
    .w_reqbuf_size          (                                 ),
    .r_reqbuf_size          (                                 )
  );
  
  assign br_master.aw_id     = '0;
  assign br_master.aw_len    = '0;
  assign br_master.aw_size   = 3'b11;
  assign br_master.aw_burst  = '0;
  assign br_master.aw_lock   = '0;
  assign br_master.aw_cache  = '0;
  assign br_master.aw_prot   = '0;
  assign br_master.aw_qos    = '0;
  assign br_master.aw_region = '0;
  assign br_master.aw_atop   = '0;
  assign br_master.w_last    = 1'b1;
  assign br_master.ar_id     = '0;
  assign br_master.ar_len    = '0;
  assign br_master.ar_size   = 3'b11;
  assign br_master.ar_burst  = '0;
  assign br_master.ar_lock   = '0;
  assign br_master.ar_cache  = '0;
  assign br_master.ar_prot   = '0;
  assign br_master.ar_qos    = '0;
  assign br_master.ar_region = '0;
  
  
  
  ariane_axi::req_t    clint_axi_req;
  ariane_axi::resp_t   clint_axi_resp;
  clint #(
    .AXI_ADDR_WIDTH ( AxiAddrWidth ),
    .AXI_DATA_WIDTH ( AxiDataWidth ),
    .AXI_ID_WIDTH   ( AxiIdWidth   ),
    .NR_CORES       ( NumHarts     )
  ) i_clint (
    .clk_i                         ,
    .rst_ni                        ,
    .testmode_i                    ,
    .axi_req_i   ( clint_axi_req  ),
    .axi_resp_o  ( clint_axi_resp ),
    .rtc_i                         ,
    .timer_irq_o                   ,
    .ipi_o
  );
  noc_axilite_bridge #(
    .SLAVE_RESP_BYTEWIDTH   ( 8             ),
    .SWAP_ENDIANESS         ( SwapEndianess )
  ) i_clint_axilite_bridge (
    .clk                    ( clk_i                         ),
    .rst                    ( ~rst_ni                       ),
    
    .splitter_bridge_val    ( buf_ariane_clint_noc2_valid_i ),
    .splitter_bridge_data   ( buf_ariane_clint_noc2_data_i  ),
    .bridge_splitter_rdy    ( ariane_clint_buf_noc2_ready_o ),
    .bridge_splitter_val    ( ariane_clint_buf_noc3_valid_o ),
    .bridge_splitter_data   ( ariane_clint_buf_noc3_data_o  ),
    .splitter_bridge_rdy    ( buf_ariane_clint_noc3_ready_i ),
    
    
    .m_axi_awaddr           ( clint_axi_req.aw.addr         ),
    .m_axi_awvalid          ( clint_axi_req.aw_valid        ),
    .m_axi_awready          ( clint_axi_resp.aw_ready       ),
    
    .m_axi_wdata            ( clint_axi_req.w.data          ),
    .m_axi_wstrb            ( clint_axi_req.w.strb          ),
    .m_axi_wvalid           ( clint_axi_req.w_valid         ),
    .m_axi_wready           ( clint_axi_resp.w_ready        ),
    
    .m_axi_araddr           ( clint_axi_req.ar.addr         ),
    .m_axi_arvalid          ( clint_axi_req.ar_valid        ),
    .m_axi_arready          ( clint_axi_resp.ar_ready       ),
    
    .m_axi_rdata            ( clint_axi_resp.r.data         ),
    .m_axi_rresp            ( clint_axi_resp.r.resp         ),
    .m_axi_rvalid           ( clint_axi_resp.r_valid        ),
    .m_axi_rready           ( clint_axi_req.r_ready         ),
    
    .m_axi_bresp            ( clint_axi_resp.b.resp         ),
    .m_axi_bvalid           ( clint_axi_resp.b_valid        ),
    .m_axi_bready           ( clint_axi_req.b_ready         ),
    
    .w_reqbuf_size          (                               ),
    .r_reqbuf_size          (                               )
  );
  
  assign clint_axi_req.aw.id     = '0;
  assign clint_axi_req.aw.len    = '0;
  assign clint_axi_req.aw.size   = 3'b11;
  assign clint_axi_req.aw.burst  = '0;
  assign clint_axi_req.aw.lock   = '0;
  assign clint_axi_req.aw.cache  = '0;
  assign clint_axi_req.aw.prot   = '0;
  assign clint_axi_req.aw.qos    = '0;
  assign clint_axi_req.aw.region = '0;
  assign clint_axi_req.aw.atop   = '0;
  assign clint_axi_req.w.last    = 1'b1;
  assign clint_axi_req.ar.id     = '0;
  assign clint_axi_req.ar.len    = '0;
  assign clint_axi_req.ar.size   = 3'b11;
  assign clint_axi_req.ar.burst  = '0;
  assign clint_axi_req.ar.lock   = '0;
  assign clint_axi_req.ar.cache  = '0;
  assign clint_axi_req.ar.prot   = '0;
  assign clint_axi_req.ar.qos    = '0;
  assign clint_axi_req.ar.region = '0;
  
  
  
  AXI_BUS #(
    .AXI_ID_WIDTH   ( AxiIdWidth   ),
    .AXI_ADDR_WIDTH ( AxiAddrWidth ),
    .AXI_DATA_WIDTH ( AxiDataWidth ),
    .AXI_USER_WIDTH ( AxiUserWidth )
  ) plic_master();
  noc_axilite_bridge #(
    
    
    
    .SLAVE_RESP_BYTEWIDTH   ( 0             ),
    .SWAP_ENDIANESS         ( SwapEndianess ),
    
    .ALIGN_RDATA            ( 0             )
  ) i_plic_axilite_bridge (
    .clk                    ( clk_i                        ),
    .rst                    ( ~rst_ni                      ),
    
    .splitter_bridge_val    ( buf_ariane_plic_noc2_valid_i ),
    .splitter_bridge_data   ( buf_ariane_plic_noc2_data_i  ),
    .bridge_splitter_rdy    ( ariane_plic_buf_noc2_ready_o ),
    .bridge_splitter_val    ( ariane_plic_buf_noc3_valid_o ),
    .bridge_splitter_data   ( ariane_plic_buf_noc3_data_o  ),
    .splitter_bridge_rdy    ( buf_ariane_plic_noc3_ready_i ),
    
    
    .m_axi_awaddr           ( plic_master.aw_addr               ),
    .m_axi_awvalid          ( plic_master.aw_valid              ),
    .m_axi_awready          ( plic_master.aw_ready              ),
    
    .m_axi_wdata            ( plic_master.w_data                ),
    .m_axi_wstrb            ( plic_master.w_strb                ),
    .m_axi_wvalid           ( plic_master.w_valid               ),
    .m_axi_wready           ( plic_master.w_ready               ),
    
    .m_axi_araddr           ( plic_master.ar_addr               ),
    .m_axi_arvalid          ( plic_master.ar_valid              ),
    .m_axi_arready          ( plic_master.ar_ready              ),
    
    .m_axi_rdata            ( plic_master.r_data                ),
    .m_axi_rresp            ( plic_master.r_resp                ),
    .m_axi_rvalid           ( plic_master.r_valid               ),
    .m_axi_rready           ( plic_master.r_ready               ),
    
    .m_axi_bresp            ( plic_master.b_resp                ),
    .m_axi_bvalid           ( plic_master.b_valid               ),
    .m_axi_bready           ( plic_master.b_ready               ),
    
    .w_reqbuf_size          ( plic_master.aw_size               ),
    .r_reqbuf_size          ( plic_master.ar_size               )
  );
  
  assign plic_master.aw_id     = '0;
  assign plic_master.aw_len    = '0;
  assign plic_master.aw_burst  = '0;
  assign plic_master.aw_lock   = '0;
  assign plic_master.aw_cache  = '0;
  assign plic_master.aw_prot   = '0;
  assign plic_master.aw_qos    = '0;
  assign plic_master.aw_region = '0;
  assign plic_master.aw_atop   = '0;
  assign plic_master.w_last    = 1'b1;
  assign plic_master.ar_id     = '0;
  assign plic_master.ar_len    = '0;
  assign plic_master.ar_burst  = '0;
  assign plic_master.ar_lock   = '0;
  assign plic_master.ar_cache  = '0;
  assign plic_master.ar_prot   = '0;
  assign plic_master.ar_qos    = '0;
  assign plic_master.ar_region = '0;
  reg_intf::reg_intf_resp_d32 plic_resp;
  reg_intf::reg_intf_req_a32_d32 plic_req;
  enum logic [2:0] {Idle, WriteSecond, ReadSecond, WriteResp, ReadResp} state_d, state_q;
  logic [31:0] rword_d, rword_q;
  
  assign rword_d = (plic_req.valid && !plic_req.write) ? plic_resp.rdata : rword_q;
  assign plic_master.r_data = {plic_resp.rdata, rword_q};
  always_ff @(posedge clk_i or negedge rst_ni) begin : p_plic_regs
    if (!rst_ni) begin
      state_q <= Idle;
      rword_q <= '0;
    end else begin
      state_q <= state_d;
      rword_q <= rword_d;
    end
  end
  
  
  always_comb begin : p_plic_if
    automatic logic [31:0] waddr, raddr;
    
    waddr = plic_master.aw_addr[31:0] - 32'(PlicBase) + 32'hc000000;
    raddr = plic_master.ar_addr[31:0] - 32'(PlicBase) + 32'hc000000;
    
    plic_master.aw_ready = plic_resp.ready;
    plic_master.w_ready  = plic_resp.ready;
    plic_master.ar_ready = plic_resp.ready;
    plic_master.r_valid  = 1'b0;
    plic_master.r_resp   = '0;
    plic_master.b_valid  = 1'b0;
    plic_master.b_resp   = '0;
    
    plic_req.valid       = 1'b0;
    plic_req.wstrb       = '0;
    plic_req.write       = 1'b0;
    plic_req.wdata       = plic_master.w_data[31:0];
    plic_req.addr        = waddr;
    
    state_d              = state_q;
    unique case (state_q)
      Idle: begin
        if (plic_master.w_valid && plic_master.aw_valid && plic_resp.ready) begin
          plic_req.valid = 1'b1;
          plic_req.write = plic_master.w_strb[3:0];
          plic_req.wstrb = '1;
          
          if (plic_master.aw_size == 3'b11) begin
            state_d = WriteSecond;
          end else begin
            state_d = WriteResp;
          end
        end else if (plic_master.ar_valid && plic_resp.ready) begin
          plic_req.valid = 1'b1;
          plic_req.addr  = raddr;
          
          if (plic_master.ar_size == 3'b11) begin
            state_d = ReadSecond;
          end else begin
            state_d = ReadResp;
          end
        end
      end
      
      WriteSecond: begin
        plic_master.aw_ready = 1'b0;
        plic_master.w_ready  = 1'b0;
        plic_master.ar_ready = 1'b0;
        plic_req.addr        = waddr + 32'h4;
        plic_req.wdata       = plic_master.w_data[63:32];
        if (plic_resp.ready && plic_master.b_ready) begin
          plic_req.valid       = 1'b1;
          plic_req.write       = 1'b1;
          plic_req.wstrb       = '1;
          plic_master.b_valid  = 1'b1;
          state_d              = Idle;
        end
      end
      
      ReadSecond: begin
        plic_master.aw_ready = 1'b0;
        plic_master.w_ready  = 1'b0;
        plic_master.ar_ready = 1'b0;
        plic_req.addr        = raddr + 32'h4;
        if (plic_resp.ready && plic_master.r_ready) begin
          plic_req.valid      = 1'b1;
          plic_master.r_valid = 1'b1;
          state_d             = Idle;
        end
      end
      WriteResp: begin
        plic_master.aw_ready = 1'b0;
        plic_master.w_ready  = 1'b0;
        plic_master.ar_ready = 1'b0;
        if (plic_master.b_ready) begin
          plic_master.b_valid  = 1'b1;
          state_d              = Idle;
        end
      end
      ReadResp: begin
        plic_master.aw_ready = 1'b0;
        plic_master.w_ready  = 1'b0;
        plic_master.ar_ready = 1'b0;
        if (plic_master.r_ready) begin
          plic_master.r_valid = 1'b1;
          state_d             = Idle;
        end
      end
      default: state_d = Idle;
    endcase
  end
  plic_top #(
    .N_SOURCE    ( NumSources      ),
    .N_TARGET    ( 2*NumHarts      ),
    .MAX_PRIO    ( PlicMaxPriority )
  ) i_plic (
    .clk_i,
    .rst_ni,
    .req_i         ( plic_req    ),
    .resp_o        ( plic_resp   ),
    .le_i          ( irq_le_i    ), 
    .irq_sources_i,                 
    .eip_targets_o ( irq_o       )
  );
endmodule 
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
module dmbr(
    input clk,
    input rst,
    input func_en, 
    input stall_en, 
   
    
    input proc_ld,
    
    input [6-1:0] creditIn_0,
    input [6-1:0] creditIn_1,
    input [6-1:0] creditIn_2,
    input [6-1:0] creditIn_3,
    input [6-1:0] creditIn_4,
    input [6-1:0] creditIn_5,
    input [6-1:0] creditIn_6,
    input [6-1:0] creditIn_7,
    input [6-1:0] creditIn_8,
    input [6-1:0] creditIn_9,
    input [16-1:0] replenishCyclesIn,
    input [10-1:0] binScaleIn,
    
    input                     l1missIn,
    input [4-1:0] l1missTag,
    input                     l2responseIn,
    input                     l2missIn,
    input [4-1:0] l2missTag,
    output reg [6-1:0] curr_cred_bin_0,
output reg [6-1:0] curr_cred_bin_1,
output reg [6-1:0] curr_cred_bin_2,
output reg [6-1:0] curr_cred_bin_3,
output reg [6-1:0] curr_cred_bin_4,
output reg [6-1:0] curr_cred_bin_5,
output reg [6-1:0] curr_cred_bin_6,
output reg [6-1:0] curr_cred_bin_7,
output reg [6-1:0] curr_cred_bin_8,
output reg [6-1:0] curr_cred_bin_9,
   
    
    output reg stallOut
);
  
reg rep_en;
reg add_counter_reset;
reg [9-1:0] sat_counter;
reg [9-1:0] add_counter;
reg [9:0] curInterval;
reg [16-1:0] stall_cycles;
reg [16-1:0] total_stall_cycles;
reg [6-1:0] curCredit_0;
reg [6-1:0] next_credit_0;
reg [6-1:0] repCredit_0;
reg req_en_0;
reg add_en_0;
reg [6-1:0] curCredit_1;
reg [6-1:0] next_credit_1;
reg [6-1:0] repCredit_1;
reg req_en_1;
reg add_en_1;
reg [6-1:0] curCredit_2;
reg [6-1:0] next_credit_2;
reg [6-1:0] repCredit_2;
reg req_en_2;
reg add_en_2;
reg [6-1:0] curCredit_3;
reg [6-1:0] next_credit_3;
reg [6-1:0] repCredit_3;
reg req_en_3;
reg add_en_3;
reg [6-1:0] curCredit_4;
reg [6-1:0] next_credit_4;
reg [6-1:0] repCredit_4;
reg req_en_4;
reg add_en_4;
reg [6-1:0] curCredit_5;
reg [6-1:0] next_credit_5;
reg [6-1:0] repCredit_5;
reg req_en_5;
reg add_en_5;
reg [6-1:0] curCredit_6;
reg [6-1:0] next_credit_6;
reg [6-1:0] repCredit_6;
reg req_en_6;
reg add_en_6;
reg [6-1:0] curCredit_7;
reg [6-1:0] next_credit_7;
reg [6-1:0] repCredit_7;
reg req_en_7;
reg add_en_7;
reg [6-1:0] curCredit_8;
reg [6-1:0] next_credit_8;
reg [6-1:0] repCredit_8;
reg req_en_8;
reg add_en_8;
reg [6-1:0] curCredit_9;
reg [6-1:0] next_credit_9;
reg [6-1:0] repCredit_9;
reg req_en_9;
reg add_en_9;
reg [3:0] bin_used_0;
reg [9:0] interval_0;
reg [9-1:0] bin_number_0;
reg [9:0] sum_counter_0;
reg [3:0] bin_used_1;
reg [9:0] interval_1;
reg [9-1:0] bin_number_1;
reg [9:0] sum_counter_1;
reg [3:0] bin_used_2;
reg [9:0] interval_2;
reg [9-1:0] bin_number_2;
reg [9:0] sum_counter_2;
reg [3:0] bin_used_3;
reg [9:0] interval_3;
reg [9-1:0] bin_number_3;
reg [9:0] sum_counter_3;
reg [3:0] bin_used_4;
reg [9:0] interval_4;
reg [9-1:0] bin_number_4;
reg [9:0] sum_counter_4;
reg [3:0] bin_used_5;
reg [9:0] interval_5;
reg [9-1:0] bin_number_5;
reg [9:0] sum_counter_5;
reg [3:0] bin_used_6;
reg [9:0] interval_6;
reg [9-1:0] bin_number_6;
reg [9:0] sum_counter_6;
reg [3:0] bin_used_7;
reg [9:0] interval_7;
reg [9-1:0] bin_number_7;
reg [9:0] sum_counter_7;
reg [3:0] bin_used_8;
reg [9:0] interval_8;
reg [9-1:0] bin_number_8;
reg [9:0] sum_counter_8;
reg [3:0] bin_used_9;
reg [9:0] interval_9;
reg [9-1:0] bin_number_9;
reg [9:0] sum_counter_9;
reg [3:0] bin_used_10;
reg [9:0] interval_10;
reg [9-1:0] bin_number_10;
reg [9:0] sum_counter_10;
reg [3:0] bin_used_11;
reg [9:0] interval_11;
reg [9-1:0] bin_number_11;
reg [9:0] sum_counter_11;
reg [3:0] bin_used_12;
reg [9:0] interval_12;
reg [9-1:0] bin_number_12;
reg [9:0] sum_counter_12;
reg [3:0] bin_used_13;
reg [9:0] interval_13;
reg [9-1:0] bin_number_13;
reg [9:0] sum_counter_13;
reg [3:0] bin_used_14;
reg [9:0] interval_14;
reg [9-1:0] bin_number_14;
reg [9:0] sum_counter_14;
reg [3:0] bin_used_15;
reg [9:0] interval_15;
reg [9-1:0] bin_number_15;
reg [9:0] sum_counter_15;
reg [6-1:0] curCredit_mux;
reg [6-1:0] repCredit_mux;
reg [6-1:0] curCredit_mux2;
reg [6-1:0] repCredit_mux2;
reg [9:0] add_interval;
reg [10-1:0] binScale;
wire [9-1:0] max_interval = (10 << binScale) + 1'b1;
wire [9-1:0] next_sat_counter = l1missIn ? {9{1'b0}} : (sat_counter < max_interval) ? sat_counter + 1'b1 : sat_counter;
wire [9-1:0] add_interval2 = add_interval > max_interval ? max_interval : add_interval[9-1:0];
wire [9-1:0] next_add_counter = (l2responseIn && add_counter_reset) ? add_interval2 : (l2responseIn && !l2missIn) ? 
                          ((add_counter + add_interval2 < max_interval) ? add_counter + add_interval2 : max_interval) :  
                              add_counter_reset ? {9{1'b0}}  : add_counter;
reg [16-1:0] repInterval;
reg rep_reset;
wire [16-1:0] next_repInterval = rep_reset ?  {16{1'b0}} : repInterval + 1'b1;
reg [16-1:0] replenishCycles;
reg stall;
reg [3:0]  bin_number;
reg [3:0]  add_bin;
wire [16-1:0] next_total_stall_cycles = stall_cycles > 0  ? total_stall_cycles + stall_cycles :
                                      total_stall_cycles > 0 ? total_stall_cycles - 1'b1 : {16{1'b0}};
wire [6-1:0] cur_credit_minus_one = curCredit_mux > 0 ? curCredit_mux - 1 : curCredit_mux;
wire [6-1:0] input2 = rep_en ? repCredit_mux2 : curCredit_mux2;
wire [9:0] sum_counter = sat_counter + add_counter;
wire [6-1:0] req_out = rep_en ? repCredit_mux : cur_credit_minus_one;
wire [6-1:0] add_out = input2 < {6{1'b1}} ? input2 + 1'b1 : input2;
always @*
begin
    rep_en = 1'b0;
    req_en_0 = 1'b0;
    req_en_1 = 1'b0; 
    req_en_2 = 1'b0;
    req_en_3 = 1'b0;
    req_en_4 = 1'b0;
    req_en_5 = 1'b0;
    req_en_6 = 1'b0;
    req_en_7 = 1'b0;
    req_en_8 = 1'b0;
    req_en_9 = 1'b0;
    stall = 1'b0;
    rep_reset = 1'b0;
    stall_cycles = 0;
    curInterval = {9+1{1'b0}} ;
    bin_number = 4'b0;
    stallOut = 1'b0;
    if (stall_en && total_stall_cycles > 0) begin
        stallOut = 1'b1;
    end
    if (repInterval == replenishCycles)
    begin
        rep_en = 1'b1;
        rep_reset = 1'b1;
    end
    if (l1missIn) begin
        curInterval = sum_counter;
        add_counter_reset = 1'b1;
    end
    else begin
        add_counter_reset = 1'b0;
        curInterval = 0;
    end
            
    if (l1missIn) begin
        if (curInterval >= 8'd9 << binScale && curCredit_9 > 0)
        begin
            req_en_9 = 1'b1;
            stall = 1'b0;
            bin_number = 9;
        end
        else if (curInterval >= 8'd8 << binScale && curCredit_8 > 0)
        begin
            req_en_8 = 1'b1;
            stall = 1'b0;
            bin_number = 8;
        end
        else if (curInterval >= 8'd7 << binScale && curCredit_7 > 0)
        begin
            req_en_7 = 1'b1;
            stall = 1'b0;
            bin_number = 7;
        end
        else if (curInterval >= 8'd6 << binScale && curCredit_6 > 0)
        begin
            req_en_6 = 1'b1;
            stall = 1'b0;
            bin_number = 6;
        end
        else if (curInterval >= 8'd5 << binScale && curCredit_5 > 0)
        begin
            req_en_5 = 1'b1;
            stall = 1'b0;
            bin_number = 5;
        end
        else if (curInterval >= 8'd4 << binScale && curCredit_4 > 0)
        begin
            req_en_4 = 1'b1;
            stall = 1'b0;
            bin_number = 4;
        end
        else if (curInterval >= 8'd3 << binScale && curCredit_3 > 0)
        begin
            req_en_3 = 1'b1;
            stall = 1'b0;
            bin_number = 3;
        end
        else if (curInterval >= 8'd2 << binScale && curCredit_2 > 0)
        begin
            req_en_2 = 1'b1;
            stall = 1'b0;
            bin_number = 2;
        end
        else if (curInterval >= 8'd1 << binScale && curCredit_1 > 0)
        begin
            req_en_1 = 1'b1;
            stall = 1'b0;
            bin_number = 1;
        end
        else if (curCredit_0 > 0)
        begin
            req_en_0 = 1'b1;
            stall = 1'b0;
            bin_number = 0;
        end
    
        else begin
            stall = 1'b1;
            if (curCredit_1 > 0)
            begin
                req_en_1 = 1'b1;
                stall_cycles = (8'd1 << binScale) - curInterval;
                bin_number = 1;
            end
            else if (curCredit_2 > 0)
            begin
                req_en_2 = 1'b1;
                stall_cycles = (8'd2 << binScale) - curInterval;
                bin_number = 2;
            end
            else if (curCredit_3 > 0)
            begin
                req_en_3 = 1'b1;
                stall_cycles = (8'd3 << binScale) - curInterval;
                bin_number = 3;
            end
            else if (curCredit_4 > 0)
            begin
                req_en_4 = 1'b1;
                stall_cycles = (8'd4 << binScale) - curInterval;
                bin_number = 4;
            end
            else if (curCredit_5 > 0)
            begin
                req_en_5 = 1'b1;
                stall_cycles = (8'd5 << binScale) - curInterval;
                bin_number = 5;
            end
            else if (curCredit_6 > 0)
            begin
                req_en_6 = 1'b1;
                stall_cycles = (8'd6 << binScale) - curInterval;
                bin_number = 6;
            end
            else if (curCredit_7 > 0)
            begin
                req_en_7 = 1'b1;
                stall_cycles = (8'd7 << binScale) - curInterval;
                bin_number = 7;
            end
            else if (curCredit_8 > 0)
            begin
                req_en_8 = 1'b1;
                stall_cycles = (8'd8 << binScale) - curInterval;
                bin_number = 8;
            end
            else if (curCredit_9 > 0)
            begin
                req_en_9 = 1'b1;
                stall_cycles = (8'd9 << binScale) - curInterval;
                bin_number = 9;
            end
            else
            begin
                req_en_0 = 1'b1;
                stall_cycles = replenishCycles - repInterval;
                bin_number = 10;
            end
        end
    end
end
always @ *
begin
    bin_number_0 = bin_used_0;
    bin_number_1 = bin_used_1;
    bin_number_2 = bin_used_2;
    bin_number_3 = bin_used_3;
    bin_number_4 = bin_used_4;
    bin_number_5 = bin_used_5;
    bin_number_6 = bin_used_6;
    bin_number_7 = bin_used_7;
    bin_number_8 = bin_used_8;
    bin_number_9 = bin_used_9;
    bin_number_10 = bin_used_10;
    bin_number_11 = bin_used_11;
    bin_number_12 = bin_used_12;
    bin_number_13 = bin_used_13;
    bin_number_14 = bin_used_14;
    bin_number_15 = bin_used_15;
    sum_counter_0 = interval_0;
    sum_counter_1 = interval_1;
    sum_counter_2 = interval_2;
    sum_counter_3 = interval_3;
    sum_counter_4 = interval_4;
    sum_counter_5 = interval_5;
    sum_counter_6 = interval_6;
    sum_counter_7 = interval_7;
    sum_counter_8 = interval_8;
    sum_counter_9 = interval_9;
    sum_counter_10 = interval_10;
    sum_counter_11 = interval_11;
    sum_counter_12 = interval_12;
    sum_counter_13 = interval_13;
    sum_counter_14 = interval_14;
    sum_counter_15 = interval_15;
    if (l1missIn) begin
        case (l1missTag) 
            4'd0: begin
                bin_number_0 = bin_number;
                sum_counter_0 = sum_counter;
            end
            4'd1: begin 
                bin_number_1 = bin_number;
                sum_counter_1 = sum_counter;
            end
            4'd2: begin
                bin_number_2 = bin_number;
                sum_counter_2 = sum_counter;
            end
            4'd3: begin
                bin_number_3 = bin_number;
                sum_counter_3 = sum_counter;
            end
            4'd4: begin
                bin_number_4 = bin_number;
                sum_counter_4 = sum_counter;
            end
            4'd5: begin 
                bin_number_5 = bin_number;
                sum_counter_5 = sum_counter;
            end
            4'd6: begin
                bin_number_6 = bin_number;
                sum_counter_6 = sum_counter;
            end
            4'd7: begin
                bin_number_7 = bin_number;
                sum_counter_7 = sum_counter;
            end
            4'd8: begin
                bin_number_8 = bin_number;
                sum_counter_8 = sum_counter;
            end
            4'd9: begin 
                bin_number_9 = bin_number;
                sum_counter_9 = sum_counter;
            end
            4'd10: begin
                bin_number_10 = bin_number;
                sum_counter_10 = sum_counter;
            end
            4'd11: begin
                bin_number_11 = bin_number;
                sum_counter_11 = sum_counter;
            end
            4'd12: begin
                bin_number_12 = bin_number;
                sum_counter_12 = sum_counter;
            end
            4'd13: begin 
                bin_number_13 = bin_number;
                sum_counter_13 = sum_counter;
            end
            4'd14: begin
                bin_number_14 = bin_number;
                sum_counter_14 = sum_counter;
            end
            4'd15: begin
                bin_number_15 = bin_number;
                sum_counter_15 = sum_counter;
            end
            default:;
        endcase
    end
end
always @ *
begin
    add_bin = 0;
    add_interval = 0;
    if (l2responseIn) begin
        if (!l2missIn) begin
            case (l2missTag)
                4'd0: begin
                    add_bin = bin_used_0;
                    add_interval = interval_0;
                end
                4'd1: begin
                    add_bin = bin_used_1;
                    add_interval = interval_1;
                end
                4'd2: begin
                    add_bin = bin_used_2;
                    add_interval = interval_2;
                end
                4'd3: begin
                    add_bin = bin_used_3;
                    add_interval = interval_3;
                end
                4'd4: begin
                    add_bin = bin_used_4;
                    add_interval = interval_4;
                end
                4'd5: begin
                    add_bin = bin_used_5;
                    add_interval = interval_5;
                end
                4'd6: begin
                    add_bin = bin_used_6;
                    add_interval = interval_6;
                end
                4'd7: begin
                    add_bin = bin_used_7;
                    add_interval = interval_7;
                end
                4'd8: begin
                    add_bin = bin_used_8;
                    add_interval = interval_8;
                end
                4'd9: begin
                    add_bin = bin_used_9;
                    add_interval = interval_9;
                end
                4'd10: begin
                    add_bin = bin_used_10;
                    add_interval = interval_10;
                end
                4'd11: begin
                    add_bin = bin_used_11;
                    add_interval = interval_11;
                end
                4'd12: begin
                    add_bin = bin_used_12;
                    add_interval = interval_12;
                end
                4'd13: begin
                    add_bin = bin_used_13;
                    add_interval = interval_13;
                end
                4'd14: begin
                    add_bin = bin_used_14;
                    add_interval = interval_14;
                end
                4'd15: begin
                    add_bin = bin_used_15;
                    add_interval = interval_15;
                end
                default: begin
                    add_bin = 10;
                    add_interval = 0;
                end
            endcase
        end
    end
end
always @ *
begin
    add_en_0 = 1'b0;
    add_en_1 = 1'b0; 
    add_en_2 = 1'b0;
    add_en_3 = 1'b0;
    add_en_4 = 1'b0;
    add_en_5 = 1'b0;
    add_en_6 = 1'b0;
    add_en_7 = 1'b0;
    add_en_8 = 1'b0;
    add_en_9 = 1'b0;
    if (l2responseIn) begin
        if (!l2missIn) begin
            case (add_bin)
               4'd0: add_en_0 = 1'b1;
               4'd1: add_en_1 = 1'b1;
               4'd2: add_en_2 = 1'b1;
               4'd3: add_en_3 = 1'b1;
               4'd4: add_en_4 = 1'b1;
               4'd5: add_en_5 = 1'b1;
               4'd6: add_en_6 = 1'b1;
               4'd7: add_en_7 = 1'b1;
               4'd8: add_en_8 = 1'b1;
               4'd9: add_en_9 = 1'b1;
               default: begin
                    add_en_0 = 1'b0;
                    add_en_1 = 1'b0; 
                    add_en_2 = 1'b0;
                    add_en_3 = 1'b0;
                    add_en_4 = 1'b0;
                    add_en_5 = 1'b0;
                    add_en_6 = 1'b0;
                    add_en_7 = 1'b0;
                    add_en_8 = 1'b0;
                    add_en_9 = 1'b0;
               end
           endcase
        end
    end 
end
always @ *
begin
    curCredit_mux = ({6{req_en_0}} & curCredit_0) | ({6{req_en_1}} & curCredit_1) | ({6{req_en_2}} & curCredit_2) | ({6{req_en_3}} & curCredit_3) | ({6{req_en_4}} & curCredit_4) | ({6{req_en_5}} & curCredit_5) | ({6{req_en_6}} & curCredit_6) | ({6{req_en_7}} & curCredit_7) | ({6{req_en_8}} & curCredit_8) | ({6{req_en_9}} & curCredit_9);
    repCredit_mux = ({6{req_en_0}} & repCredit_0) | ({6{req_en_1}} & repCredit_1) | ({6{req_en_2}} & repCredit_2) | ({6{req_en_3}} & repCredit_3) | ({6{req_en_4}} & repCredit_4) | ({6{req_en_5}} & repCredit_5) | ({6{req_en_6}} & repCredit_6) | ({6{req_en_7}} & repCredit_7) | ({6{req_en_8}} & repCredit_8) | ({6{req_en_9}} & repCredit_9);
end
always @ *
begin
    curCredit_mux2 = ({6{add_en_0}} & curCredit_0) | ({6{add_en_1}} & curCredit_1) | ({6{add_en_2}} & curCredit_2) | ({6{add_en_3}} & curCredit_3) | ({6{add_en_4}} & curCredit_4) | ({6{add_en_5}} & curCredit_5) | ({6{add_en_6}} & curCredit_6) | ({6{add_en_7}} & curCredit_7) | ({6{add_en_8}} & curCredit_8) | ({6{add_en_9}} & curCredit_9);
    repCredit_mux2 = ({6{add_en_0}} & repCredit_0) | ({6{add_en_1}} & repCredit_1) | ({6{add_en_2}} & repCredit_2) | ({6{add_en_3}} & repCredit_3) | ({6{add_en_4}} & repCredit_4) | ({6{add_en_5}} & repCredit_5) | ({6{add_en_6}} & repCredit_6) | ({6{add_en_7}} & repCredit_7) | ({6{add_en_8}} & repCredit_8) | ({6{add_en_9}} & repCredit_9);
end
always @ *
begin
    next_credit_0 = curCredit_0;
    case({req_en_0, rep_en, add_en_0})
        3'b001: next_credit_0  = add_out;
        3'b010: next_credit_0 = repCredit_0;
        3'b011: next_credit_0 = add_out;
        3'b100: next_credit_0 = req_out;
        3'b110: next_credit_0 = req_out;
        3'b111: next_credit_0 = repCredit_0;
        3'b000: next_credit_0 = curCredit_0;
        3'b101: next_credit_0 = curCredit_0;
        default:;
    endcase
end
always @ *
begin
    next_credit_1 = curCredit_1;
    case({req_en_1, rep_en, add_en_1})
        3'b001: next_credit_1 = add_out;
        3'b010: next_credit_1 = repCredit_1;
        3'b011: next_credit_1 = add_out;
        3'b100: next_credit_1 = req_out;
        3'b110: next_credit_1 = req_out;
        3'b111: next_credit_1 = repCredit_1;
        3'b000: next_credit_1 = curCredit_1;
        3'b101: next_credit_1 = curCredit_1;
        default:;
    endcase
end
always @ *
begin
    next_credit_2 = curCredit_2;
    case({req_en_2, rep_en, add_en_2})
        3'b001: next_credit_2  = add_out;
        3'b010: next_credit_2 = repCredit_2;
        3'b011: next_credit_2 = add_out;
        3'b100: next_credit_2 = req_out;
        3'b110: next_credit_2 = req_out;
        3'b111: next_credit_2 = repCredit_2;
        3'b000: next_credit_2 = curCredit_2;
        3'b101: next_credit_2 = curCredit_2;
        default:;
    endcase
end
always @ *
begin
    next_credit_3 = curCredit_3;
    case({req_en_3, rep_en, add_en_3})
        3'b001: next_credit_3  = add_out;
        3'b010: next_credit_3 = repCredit_3;
        3'b011: next_credit_3 = add_out;
        3'b100: next_credit_3 = req_out;
        3'b110: next_credit_3 = req_out;
        3'b111: next_credit_3 = repCredit_3;
        3'b000: next_credit_3 = curCredit_3;
        3'b101: next_credit_3 = curCredit_3;
        default:;
    endcase
end
always @ *
begin
    next_credit_4 = curCredit_4;
    case({req_en_4, rep_en, add_en_4})
        3'b001: next_credit_4  = add_out;
        3'b010: next_credit_4 = repCredit_4;
        3'b011: next_credit_4 = add_out;
        3'b100: next_credit_4 = req_out;
        3'b110: next_credit_4 = req_out;
        3'b111: next_credit_4 = repCredit_4;
        3'b000: next_credit_4 = curCredit_4;
        3'b101: next_credit_4 = curCredit_4;
        default:;
    endcase
end
always @ *
begin
    next_credit_5 = curCredit_5;
    case({req_en_5, rep_en, add_en_5})
        3'b001: next_credit_5 = add_out;
        3'b010: next_credit_5 = repCredit_5;
        3'b011: next_credit_5 = add_out;
        3'b100: next_credit_5 = req_out;
        3'b110: next_credit_5 = req_out;
        3'b111: next_credit_5 = repCredit_5;
        3'b000: next_credit_5 = curCredit_5;
        3'b101: next_credit_5 = curCredit_5;
        default:;
    endcase
end
always @ *
begin
    next_credit_6 = curCredit_6;
    case({req_en_6, rep_en, add_en_6})
        3'b001: next_credit_6 = add_out;
        3'b010: next_credit_6 = repCredit_6;
        3'b011: next_credit_6 = add_out;
        3'b100: next_credit_6 = req_out;
        3'b110: next_credit_6 = req_out;
        3'b111: next_credit_6 = repCredit_6;
        3'b000: next_credit_6 = curCredit_6;
        3'b101: next_credit_6 = curCredit_6;
        default:;
    endcase
end
always @ *
begin
    next_credit_7 = curCredit_7;
    case({req_en_7, rep_en, add_en_7})
        3'b001: next_credit_7 = add_out;
        3'b010: next_credit_7 = repCredit_7;
        3'b011: next_credit_7 = add_out;
        3'b100: next_credit_7 = req_out;
        3'b110: next_credit_7 = req_out;
        3'b111: next_credit_7 = repCredit_7;
        3'b000: next_credit_7 = curCredit_7;
        3'b101: next_credit_7 = curCredit_7;
        default:;
    endcase
end
always @ *
begin
    next_credit_8 = curCredit_8;
    case({req_en_8, rep_en, add_en_8})
        3'b001: next_credit_8 = add_out;
        3'b010: next_credit_8 = repCredit_8;
        3'b011: next_credit_8 = add_out;
        3'b100: next_credit_8 = req_out;
        3'b110: next_credit_8 = req_out;
        3'b111: next_credit_8 = repCredit_8;
        3'b000: next_credit_8 = curCredit_8;
        3'b101: next_credit_8 = curCredit_8;
        default:;
    endcase
end
always @ *
begin
    next_credit_9 = curCredit_9;
    case({req_en_9, rep_en, add_en_9})
        3'b001: next_credit_9 = add_out;
        3'b010: next_credit_9 = repCredit_9;
        3'b011: next_credit_9 = add_out;
        3'b100: next_credit_9 = req_out;
        3'b110: next_credit_9 = req_out;
        3'b111: next_credit_9 = repCredit_9;
        3'b000: next_credit_9 = curCredit_9;
        3'b101: next_credit_9 = curCredit_9;
        default:;
    endcase
end
always @*
begin
    curr_cred_bin_0 = curCredit_0;
curr_cred_bin_1 = curCredit_1;
curr_cred_bin_2 = curCredit_2;
curr_cred_bin_3 = curCredit_3;
curr_cred_bin_4 = curCredit_4;
curr_cred_bin_5 = curCredit_5;
curr_cred_bin_6 = curCredit_6;
curr_cred_bin_7 = curCredit_7;
curr_cred_bin_8 = curCredit_8;
curr_cred_bin_9 = curCredit_9;
 
end
always @ (posedge clk)
begin
    if (rst)
    begin
        repCredit_0 <= {6{1'b0}};
        repCredit_1 <= {6{1'b0}};
        repCredit_2 <= {6{1'b0}};
        repCredit_3 <= {6{1'b0}};
        repCredit_4 <= {6{1'b0}};
        repCredit_5 <= {6{1'b0}};
        repCredit_6 <= {6{1'b0}};
        repCredit_7 <= {6{1'b0}};
        repCredit_8 <= {6{1'b0}};
        repCredit_9 <= {6{1'b0}};
        repInterval <= {16{1'b0}};
        total_stall_cycles <= {16{1'b0}};
        interval_0 <= {9+1{1'b0}};
        interval_1 <= {9+1{1'b0}};
        interval_2 <= {9+1{1'b0}};
        interval_3 <= {9+1{1'b0}};
        interval_4 <= {9+1{1'b0}};
        interval_5 <= {9+1{1'b0}};
        interval_6 <= {9+1{1'b0}};
        interval_7 <= {9+1{1'b0}};
        interval_8 <= {9+1{1'b0}};
        interval_9 <= {9+1{1'b0}};
        interval_10 <= {9+1{1'b0}};
        interval_11 <= {9+1{1'b0}};
        interval_12 <= {9+1{1'b0}};
        interval_13 <= {9+1{1'b0}};
        interval_14 <= {9+1{1'b0}};
        interval_15 <= {9+1{1'b0}};
        bin_used_0 <= 4'b0;
        bin_used_1 <= 4'b0;
        bin_used_2 <= 4'b0;
        bin_used_3 <= 4'b0;
        bin_used_4 <= 4'b0;
        bin_used_5 <= 4'b0;
        bin_used_6 <= 4'b0;
        bin_used_7 <= 4'b0;
        bin_used_8 <= 4'b0;
        bin_used_9 <= 4'b0;
        bin_used_10 <= 4'b0;
        bin_used_11 <= 4'b0;
        bin_used_12 <= 4'b0;
        bin_used_13 <= 4'b0;
        bin_used_14 <= 4'b0;
        bin_used_15 <= 4'b0;
        sat_counter <= {9{1'b0}};
        add_counter <= {9{1'b0}};
        replenishCycles <= {16{1'b0}};
        binScale <= {10{1'b0}};
    end
    else if (func_en)
    begin
        if (proc_ld) begin
            repCredit_0 <= creditIn_0;
            repCredit_1 <= creditIn_1;
            repCredit_2 <= creditIn_2;
            repCredit_3 <= creditIn_3;
            repCredit_4 <= creditIn_4;
            repCredit_5 <= creditIn_5;
            repCredit_6 <= creditIn_6;
            repCredit_7 <= creditIn_7;
            repCredit_8 <= creditIn_8;
            repCredit_9 <= creditIn_9;
            replenishCycles <= replenishCyclesIn;
            binScale <= binScaleIn;
        end
        sat_counter <= next_sat_counter; 
        add_counter <= next_add_counter;
        bin_used_0 <= bin_number_0;
        bin_used_1 <= bin_number_1;
        bin_used_2 <= bin_number_2;
        bin_used_3 <= bin_number_3;
        bin_used_4 <= bin_number_4;
        bin_used_5 <= bin_number_5;
        bin_used_6 <= bin_number_6;
        bin_used_7 <= bin_number_7;
        bin_used_8 <= bin_number_8;
        bin_used_9 <= bin_number_9;
        bin_used_10 <= bin_number_10;
        bin_used_11 <= bin_number_11;
        bin_used_12 <= bin_number_12;
        bin_used_13 <= bin_number_13;
        bin_used_14 <= bin_number_14;
        bin_used_15 <= bin_number_15;
        interval_0 <= sum_counter_0;
        interval_1 <= sum_counter_1;
        interval_2 <= sum_counter_2;
        interval_3 <= sum_counter_3;
        interval_4 <= sum_counter_4;
        interval_5 <= sum_counter_5;
        interval_6 <= sum_counter_6;
        interval_7 <= sum_counter_7;
        interval_8 <= sum_counter_8;
        interval_9 <= sum_counter_9;
        interval_10 <= sum_counter_10;
        interval_11 <= sum_counter_11;
        interval_12 <= sum_counter_12;
        interval_13 <= sum_counter_13;
        interval_14 <= sum_counter_14;
        interval_15 <= sum_counter_15;
        total_stall_cycles <= next_total_stall_cycles;
        repInterval <= next_repInterval;
        
    end
end
always @ (posedge clk)
begin
    if (rst) begin 
        curCredit_0 <= 1;
        curCredit_1 <= 1;
        curCredit_2 <= 1;
        curCredit_3 <= 1;
        curCredit_4 <= 1;
        curCredit_5 <= 1;
        curCredit_6 <= 1;
        curCredit_7 <= 1;
        curCredit_8 <= 1;
        curCredit_9 <= 1;
    end
    else if (proc_ld && func_en) begin
        curCredit_0 <= creditIn_0;
        curCredit_1 <= creditIn_1;
        curCredit_2 <= creditIn_2;
        curCredit_3 <= creditIn_3;
        curCredit_4 <= creditIn_4;
        curCredit_5 <= creditIn_5;
        curCredit_6 <= creditIn_6;
        curCredit_7 <= creditIn_7;
        curCredit_8 <= creditIn_8;
        curCredit_9 <= creditIn_9;
    end
    else if (func_en) begin
        curCredit_0 <= next_credit_0;
        curCredit_1 <= next_credit_1;
        curCredit_2 <= next_credit_2;
        curCredit_3 <= next_credit_3;
        curCredit_4 <= next_credit_4;
        curCredit_5 <= next_credit_5;
        curCredit_6 <= next_credit_6;
        curCredit_7 <= next_credit_7;
        curCredit_8 <= next_credit_8;
        curCredit_9 <= next_credit_9;
    end
end
  
    
endmodule
module bus_compare_equal (a, b, bus_equal);
    parameter WIDTH = 8;
    parameter BHC = 10;
    input [WIDTH-1:0] a, b;
    output wire bus_equal;
    assign bus_equal = (a==b) ? 1'b1 : 1'b0;
endmodule
module flip_bus (in, out);
    parameter WIDTH = 8;
    parameter BHC = 10;
    input [WIDTH-1:0] in;
    output wire [WIDTH-1:0] out;
    
    assign out = ~in;
endmodule
module one_of_eight(in0,in1,in2,in3,in4,in5,in6,in7,sel,out);
    parameter WIDTH = 8;
    parameter BHC = 10;
    input [2:0] sel;
    input [WIDTH-1:0] in0,in1,in2,in3,in4,in5,in6,in7;
    output reg [WIDTH-1:0] out;
    always@ (*)
    begin
        out={WIDTH{1'b0}};
        case(sel)
            3'd0:out=in0;
            3'd1:out=in1;
            3'd2:out=in2;
            3'd3:out=in3;
            3'd4:out=in4;
            3'd5:out=in5;
            3'd6:out=in6;
            3'd7:out=in7;
            default:; 
        endcase
    end
endmodule
module one_of_five(in0,in1,in2,in3,in4,sel,out);
    parameter WIDTH = 8;
    parameter BHC = 10;
    input [2:0] sel;
    input [WIDTH-1:0] in0,in1,in2,in3,in4;
    output reg [WIDTH-1:0] out;
    always@(*)
    begin
        out={WIDTH{1'b0}};
        case(sel)
            3'd0:out=in0;
            3'd1:out=in1;
            3'd2:out=in2;
            3'd3:out=in3;
            3'd4:out=in4;
            default:; 
        endcase
    end
endmodule
module net_dff #(parameter WIDTH=8, parameter BHC=10) 
    (input wire [WIDTH-1:0] d, 
    output reg [WIDTH-1:0] q,
    input wire clk);
always @ (posedge clk)
begin
    q <= d;
end
endmodule
module one_of_n(
  
  in0,
  in1,
  sel,
  out);
    parameter WIDTH = 8;
    parameter BHC = 10;
    input [0:0] sel;
    input [WIDTH-1:0] in0,in1;
    output reg [WIDTH-1:0] out;
    always@(*)
    begin
        out={WIDTH{1'b0}};
        case(sel)
        
            1'd0:out=in0;
            1'd1:out=in1;
            default:; 
        endcase
    end
endmodule
module one_of_n_plus_3(
  
  in0,
  in1,
  in2,
  in3,
  in4,
  sel,
  out);
    parameter WIDTH = 8;
    parameter BHC = 10;
    input [2:0] sel;
    
    input [WIDTH-1:0] in0,in1,in2,in3,in4;
    output reg [WIDTH-1:0] out;
    always@(*)
    begin
        out={WIDTH{1'b0}};
        case(sel)
        
            3'd0:out=in0;
            3'd1:out=in1;
            3'd2:out=in2;
            3'd3:out=in3;
            3'd4:out=in4;
            default:; 
        endcase
    end
endmodule
module fpga_bridge_rcv_32 (
    rst, 
    wr_clk,
    rd_clk,
    credit_rd_clk,
    bout_data_1,
    bout_val_1,
    bout_rdy_1,
    bout_data_2,
    bout_val_2,
    bout_rdy_2,
    bout_data_3,
    bout_val_3,
    bout_rdy_3,
    data_from_chip,
    data_channel,
    credit_to_chip
); 
input rst;
input wr_clk;
input rd_clk;
input credit_rd_clk;
input bout_rdy_1;
input bout_rdy_2;
input bout_rdy_3;
input [31:0] data_from_chip;
input [ 1:0] data_channel;
output [63:0]   bout_data_1;
output          bout_val_1;
output [63:0]   bout_data_2;
output          bout_val_2;
output [63:0]   bout_data_3;
output          bout_val_3;
output [2:0]    credit_to_chip;
wire sort_rdy_1;
wire sort_rdy_2;
wire sort_rdy_3;
wire [63:0] sort_data_1;
wire [63:0] sort_data_2;
wire [63:0] sort_data_3;
wire sort_val_1;
wire sort_val_2;
wire sort_val_3;
wire fifo1_full;
wire fifo2_full;
wire fifo3_full;
wire credit_fifo_full;
reg [31:0] data_from_chip_f ;
reg  [1:0] data_channel_f ;
reg [31:0] data_from_chip_ff; 
reg  [1:0] data_channel_ff; 
reg [31:0] data_from_chip_fff; 
reg  [1:0] data_channel_fff; 
reg [31:0] channel_buffer;
reg [0:0]  channel_buffer_count;
wire [63:0] buffered_data;
reg [1:0] buffered_channel;
reg wr_rst_f;
reg wr_rst_ff;
reg rd_rst_f;
reg rd_rst_ff;
reg credit_rd_rst_f;
reg credit_rd_rst_ff;
always @ (posedge wr_clk)
begin
    wr_rst_f <= rst;
    wr_rst_ff <= wr_rst_f;
end
always @ (posedge rd_clk)
begin
    rd_rst_f <= rst;
    rd_rst_ff <= rd_rst_f;
end
always @ (posedge credit_rd_clk)
begin
    credit_rd_rst_f <= rst;
    credit_rd_rst_ff <= credit_rd_rst_f;
end
assign sort_data_1 = (buffered_channel == 2'b01 && buffered_channel == data_channel_fff && channel_buffer_count == 1'b1) ? buffered_data : 64'd0;
assign sort_data_2 = (buffered_channel == 2'b10 && buffered_channel == data_channel_fff && channel_buffer_count == 1'b1) ? buffered_data : 64'd0;
assign sort_data_3 = (buffered_channel == 2'b11 && buffered_channel == data_channel_fff && channel_buffer_count == 1'b1) ? buffered_data : 64'd0;
assign sort_val_1  = (buffered_channel == 2'b01 && buffered_channel == data_channel_fff && channel_buffer_count == 1'b1) ? 1'b1 : 1'b0;
assign sort_val_2  = (buffered_channel == 2'b10 && buffered_channel == data_channel_fff && channel_buffer_count == 1'b1) ? 1'b1 : 1'b0;
assign sort_val_3  = (buffered_channel == 2'b11 && buffered_channel == data_channel_fff && channel_buffer_count == 1'b1) ? 1'b1 : 1'b0;
assign buffered_data = {data_from_chip_fff, channel_buffer};
always @(posedge wr_clk) begin
    data_from_chip_f <= data_from_chip;
    data_from_chip_ff <= data_from_chip_f;
    data_from_chip_fff <= data_from_chip_ff;
end
always @(posedge wr_clk) begin
    if(wr_rst_ff) begin
        buffered_channel <= 2'd0;
        channel_buffer_count <= 0;
        data_channel_f <= 2'd0;
        data_channel_ff <= 2'd0;
        data_channel_fff <= 2'd0;
    end
    else begin
        if(!channel_buffer_count && data_channel_fff != 0) begin 
            channel_buffer <= data_from_chip_fff;
            buffered_channel <= data_channel_fff;
            channel_buffer_count <= channel_buffer_count + 1'b1;
        end
        else if (channel_buffer_count && buffered_channel == data_channel_fff) begin
            channel_buffer_count <= 1'b0;
            buffered_channel <= 2'b00;
        end
        data_channel_f <= data_channel;
        data_channel_ff <= data_channel_f;
        data_channel_fff <= data_channel_ff;
    end
end
wire          bout_val_pre1;
wire          bout_val_pre2;
wire          bout_val_pre3;
reg           bout_val_buf1;
reg           bout_val_buf2;
reg           bout_val_buf3;
wire fifo1_empty;
    async_fifo #(
    .DSIZE(64),
    .ASIZE(9),
    .MEMSIZE(256) )
    async_fifo_1(
        .rreset(rd_rst_ff),
        .wreset(wr_rst_ff),
        .wclk(wr_clk),
        .rclk(rd_clk),
        .ren(bout_rdy_1 & ~credit_fifo_full),
        .wval(sort_val_1),
        .wdata(sort_data_1),
        .rdata(bout_data_1),
        .wfull(fifo1_full), 
        .rempty(fifo1_empty)
    );
assign bout_val_1 = ~fifo1_empty & ~credit_fifo_full;
wire fifo2_empty;
    async_fifo #(
    .DSIZE(64),
    .ASIZE(9),
    .MEMSIZE(256) )
    async_fifo_2(
        .rreset(rd_rst_ff),
        .wreset(wr_rst_ff),
        .wclk(wr_clk),
        .rclk(rd_clk),
        .ren(bout_rdy_2 & ~credit_fifo_full),
        .wval(sort_val_2),
        .wdata(sort_data_2),
        .rdata(bout_data_2),
        .wfull(fifo2_full), 
        .rempty(fifo2_empty)
    );
assign bout_val_2 = ~fifo2_empty & ~credit_fifo_full;
wire fifo3_empty;
    async_fifo #(
    .DSIZE(64),
    .ASIZE(9),
    .MEMSIZE(256) )
    async_fifo_3(
        .rreset(rd_rst_ff),
        .wreset(wr_rst_ff),
        .wclk(wr_clk),
        .rclk(rd_clk),
        .ren(bout_rdy_3 & ~credit_fifo_full),
        .wval(sort_val_3),
        .wdata(sort_data_3),
        .rdata(bout_data_3),
        .wfull(fifo3_full), 
        .rempty(fifo3_empty)
    );
assign bout_val_3 = ~fifo3_empty & ~credit_fifo_full;
wire [2:0] credit_gather;
wire credit_val;
wire [2:0] credit_fifo_out;
reg  [2:0] credit_to_chip_r ;
reg  [2:0] credit_fifo_out_f;
wire credit_empty;
    async_fifo #(
    .DSIZE(3),
    .ASIZE(11),
    .MEMSIZE(1024) )
    async_credit_fifo(
        .rreset(credit_rd_rst_ff),
        .wreset(rd_rst_ff),
        .wclk(rd_clk),
        .rclk(credit_rd_clk),
        .ren(~credit_rd_rst_ff),
        .wval(~rd_rst_ff & (| credit_gather)),
        .wdata(credit_gather),
        .rdata(credit_fifo_out),
        .wfull(credit_fifo_full),   
        .rempty(credit_empty)
    );
assign credit_val = ~ credit_empty;
assign credit_to_chip = credit_to_chip_r;
assign credit_gather[0] = bout_val_1 & bout_rdy_1;
assign credit_gather[1] = bout_val_2 & bout_rdy_2;
assign credit_gather[2] = bout_val_3 & bout_rdy_3;
always@(posedge credit_rd_clk) begin
   if(credit_rd_rst_ff) begin
        credit_to_chip_r <= 3'b000;
        credit_fifo_out_f <= 3'b000;
   end
   else begin
       credit_to_chip_r <= credit_fifo_out_f;
       if(credit_val) begin 
           credit_fifo_out_f <= credit_fifo_out;
       end
       else
           credit_fifo_out_f <= 3'b000;
   end 
end
endmodule
module fpga_bridge_send_32 (
    rst, 
    wr_clk,
    rd_clk,
    credit_wr_clk,
    bin_data_1,
    bin_val_1,
    bin_rdy_1,
    bin_data_2,
    bin_val_2,
    bin_rdy_2,
    bin_data_3,
    bin_val_3,
    bin_rdy_3,
    data_to_chip,
    data_channel,
    credit_from_chip
);  
parameter FULL_THRESHOLD = 9'd255;
input rst;
input wr_clk;
input rd_clk;
input credit_wr_clk;
output          bin_rdy_1;
output          bin_rdy_2;
output          bin_rdy_3;
output [31:0]   data_to_chip;
output [ 1:0]    data_channel;
input [63:0]    bin_data_1;
input           bin_val_1;
input [63:0]    bin_data_2;
input           bin_val_2;
input [63:0]    bin_data_3;
input           bin_val_3;
input [2:0]     credit_from_chip;
wire network_rdy_1;
wire network_rdy_2;
wire network_rdy_3;
wire fifo1_full;
wire fifo2_full;
wire fifo3_full;
wire [63:0] network_data_1;
wire [63:0] network_data_2;
wire [63:0] network_data_3;
wire network_val_1;
wire network_val_2;
wire network_val_3;
wire network_empty_1;
wire network_empty_2;
wire network_empty_3;
wire [63:0] data_to_serial_buffer;
reg  [31:0] serial_buffer_data; 
reg  [31:0] serial_buffer_data_f ;
reg  [31:0] serial_buffer_data_next;
reg   [0:0] serial_buffer_data_counter;
wire  [1:0] channel_to_serial_buffer;
reg   [1:0] serial_buffer_channel; 
reg   [1:0] serial_buffer_channel_f ;
reg   [2:0] credit_from_chip_f ;
reg   [2:0] credit_from_chip_ff; 
reg         credit_fifo_wren_f;
wire  [2:0] credit_fifo_out;
wire        credit_fifo_full;
wire        credit_fifo_empty;
reg   [2:0] credit_fifo_out_f;
reg wr_rst_f;
reg wr_rst_ff;
reg rd_rst_f;
reg rd_rst_ff;
reg credit_wr_rst_f;
reg credit_wr_rst_ff;
always @ (posedge wr_clk)
begin
    wr_rst_f <= rst;
    wr_rst_ff <= wr_rst_f;
end
always @ (posedge rd_clk)
begin
    rd_rst_f <= rst;
    rd_rst_ff <= rd_rst_f;
end
always @ (posedge credit_wr_clk)
begin
    credit_wr_rst_f <= rst;
    credit_wr_rst_ff <= credit_wr_rst_f;
end
assign bin_rdy_1 = ~fifo1_full; 
assign bin_rdy_2 = ~fifo2_full; 
assign bin_rdy_3 = ~fifo3_full; 
assign data_to_chip = serial_buffer_data_f;
assign data_channel = serial_buffer_channel_f;
bridge_network_chooser_32 #(
    .FULL_THRESHOLD(FULL_THRESHOLD)
)separator(
    .rst    (rd_rst_ff),
    .clk    (rd_clk),
    .data_out(data_to_serial_buffer),
    .data_channel(channel_to_serial_buffer),
    .val_1  (network_val_1),
    .val_2  (network_val_2),
    .val_3  (network_val_3),
    .din_1  (network_data_1),
    .din_2  (network_data_2),
    .din_3  (network_data_3),
    .rdy_1  (network_rdy_1),
    .rdy_2  (network_rdy_2),
    .rdy_3  (network_rdy_3),
    .credit_from_chip(credit_fifo_out_f)
);
    async_fifo #(
    .DSIZE(64),
    .ASIZE(9),
    .MEMSIZE(256) )
    async_fifo_1(
        .rreset(rd_rst_ff),
        .wreset(wr_rst_ff),
        .wclk(wr_clk),
        .rclk(rd_clk),
        .ren(network_rdy_1),
        .wval(bin_val_1),
        .wdata(bin_data_1),
        .rdata(network_data_1),
        .wfull(fifo1_full),
        .rempty(network_empty_1)
    );
    async_fifo #(
    .DSIZE(64),
    .ASIZE(9),
    .MEMSIZE(256) )
    async_fifo_2(
        .rreset(rd_rst_ff),
        .wreset(wr_rst_ff),
        .wclk(wr_clk),
        .rclk(rd_clk),
        .ren(network_rdy_2),
        .wval(bin_val_2),
        .wdata(bin_data_2),
        .rdata(network_data_2),
        .wfull(fifo2_full),
        .rempty(network_empty_2)
    );
    async_fifo #(
    .DSIZE(64),
    .ASIZE(9),
    .MEMSIZE(256) )
    async_fifo_3(
        .rreset(rd_rst_ff),
        .wreset(wr_rst_ff),
        .wclk(wr_clk),
        .rclk(rd_clk),
        .ren(network_rdy_3),
        .wval(bin_val_3),
        .wdata(bin_data_3),
        .rdata(network_data_3),
        .wfull(fifo3_full),
        .rempty(network_empty_3)
    );
assign network_val_1 = ~network_empty_1;
assign network_val_2 = ~network_empty_2;
assign network_val_3 = ~network_empty_3;
always @(posedge rd_clk) begin
    if(rd_rst_ff) begin
        serial_buffer_channel <= 2'd0;
        serial_buffer_data_counter <= 1'b1;
        serial_buffer_channel_f <= 2'd0;
    end
    else begin
        if( channel_to_serial_buffer != 0 && serial_buffer_data_counter == 1) begin
            
            serial_buffer_data <= data_to_serial_buffer[31:0];
            serial_buffer_data_next <= data_to_serial_buffer[63:32];
            serial_buffer_channel <= channel_to_serial_buffer;
            serial_buffer_data_counter <= serial_buffer_data_counter + 1'b1;
        end
        else if( serial_buffer_channel != 0 && serial_buffer_data_counter != 1'b1) begin
            serial_buffer_data <= serial_buffer_data_next;
            
            serial_buffer_data_counter <= serial_buffer_data_counter + 1'b1;
        end
        else begin
            serial_buffer_data_counter <= 1'b1;
            serial_buffer_channel <= channel_to_serial_buffer;
        end
        serial_buffer_data_f <= serial_buffer_data;
        serial_buffer_channel_f <= serial_buffer_channel;
    end
end
    async_fifo #(
    .DSIZE(3),
    .ASIZE(11),
    .MEMSIZE(1024) )
    async_credit_fifo(
        .rreset(rd_rst_ff),
        .wreset(credit_wr_rst_ff),
        .wclk(credit_wr_clk),
        .rclk(rd_clk),
        .ren(~rd_rst_ff),
        .wval(~credit_wr_rst_ff & credit_fifo_wren_f),
        .wdata(credit_from_chip_ff),
        .rdata(credit_fifo_out),
        .wfull(credit_fifo_full),
        .rempty(credit_fifo_empty)
    );
always @(posedge credit_wr_clk) begin
    if(credit_wr_rst_ff) begin
       credit_fifo_wren_f <= 1'b0; 
    end
    else begin
        credit_fifo_wren_f <= |credit_from_chip_f;
    end
end
always @ (posedge credit_wr_clk) begin
    
    credit_from_chip_f <= credit_from_chip;
    credit_from_chip_ff <= credit_from_chip_f; 
end
always @(posedge rd_clk) begin
    if(rd_rst_ff) begin
        credit_fifo_out_f <= 3'd0;
    end
    else begin
        if (~credit_fifo_empty)
            credit_fifo_out_f <= credit_fifo_out;
        else
            credit_fifo_out_f <= 3'd0;
    end
end
endmodule
module bridge_network_chooser_32 (
    rst,
    clk,
    data_out,
    data_channel,
    din_1,
    rdy_1,
    val_1,
    din_2,
    rdy_2,
    val_2,
    din_3,
    rdy_3,
    val_3,
    credit_from_chip
);
input rst;
input clk;
input [63:0] din_1;
input [63:0] din_2;
input [63:0] din_3;
input        val_1;
input        val_2;
input        val_3;
input [ 2:0] credit_from_chip;
output [63:0] data_out;
output [ 1:0] data_channel;
output        rdy_1;
output        rdy_2;
output        rdy_3;
reg [8:0] credit_1; 
reg [8:0] credit_2;
reg [8:0] credit_3;
wire [1:0] select;
reg  [1:0] select_reg;
reg  [0:0] select_counter;
reg sel_23;
reg sel_13;
reg sel_12;
reg [1:0] sel_123;
parameter FULL_THRESHOLD = 9'd255;
reg rdy_1_f;
reg rdy_2_f;
reg rdy_3_f;
wire rdy_1_next;
wire rdy_2_next;
wire rdy_3_next;
assign data_out =   rdy_1_f ? din_1 :
                    rdy_2_f ? din_2 :
                    rdy_3_f ? din_3 : 64'd0;
assign data_channel = select_reg; 
assign rdy_1 = rdy_1_f;
assign rdy_2 = rdy_2_f;
assign rdy_3 = rdy_3_f;
assign rdy_1_next = (select == 2'b01 && select_counter == 1'b0) ? 1'b1 : 1'b0;
assign rdy_2_next = (select == 2'b10 && select_counter == 1'b0) ? 1'b1 : 1'b0;
assign rdy_3_next = (select == 2'b11 && select_counter == 1'b0) ? 1'b1 : 1'b0;
assign select = ( (select_counter != 1'b0         ) )   ? select_reg :
                ( (credit_1 == FULL_THRESHOLD || ~val_1) &&            
                  (credit_2 == FULL_THRESHOLD || ~val_2) && 
                  (credit_3 == FULL_THRESHOLD || ~val_3) )   ? 2'b00  :
                ( (credit_2 == FULL_THRESHOLD || ~val_2) &&            
                  (credit_3 == FULL_THRESHOLD || ~val_3) )   ? 2'b01  :
                ( (credit_1 == FULL_THRESHOLD || ~val_1) &&
                  (credit_3 == FULL_THRESHOLD || ~val_3) )   ? 2'b10  :
                ( (credit_1 == FULL_THRESHOLD || ~val_1) &&
                  (credit_2 == FULL_THRESHOLD || ~val_2) )   ? 2'b11  :
                ( (credit_1 == FULL_THRESHOLD || ~val_1) )   ? (sel_23 ? 2'b11 : 2'b10) : 
                ( (credit_2 == FULL_THRESHOLD || ~val_2) )   ? (sel_13 ? 2'b11 : 2'b01) :
                ( (credit_3 == FULL_THRESHOLD || ~val_3) )   ? (sel_12 ? 2'b10 : 2'b01) :
                                                sel_123; 
always @(posedge clk) begin
    if(rst) begin
        rdy_1_f <= 1'b0;
        rdy_2_f <= 1'b0;
        rdy_3_f <= 1'b0;
    end
    else begin
        rdy_1_f <= rdy_1_next;
        rdy_2_f <= rdy_2_next;
        rdy_3_f <= rdy_3_next;
    end
end
always @(posedge clk) begin
    if(rst) begin
        select_reg <= 2'd0;
    end
    else begin
        select_reg <= select;
    end
end
always @(posedge clk) begin
    if(rst) begin
        credit_1 <= 9'd0;
        credit_2 <= 9'd0;
        credit_3 <= 9'd0;
        sel_23 <= 0;
        sel_13 <= 0;
        sel_12 <= 0;
        sel_123 <= 0;
        select_counter <= 0;
    end
    else begin
        
        if(select == 0) begin
            select_counter <= 0;
        end
        else begin
            select_counter <= select_counter + 2'b01; 
        end
        
        if(credit_from_chip[0] & ~(rdy_1 & val_1)) begin
            credit_1 <= credit_1 - 9'd1;
        end
        if(credit_from_chip[1] & ~(rdy_2 & val_2)) begin
            credit_2 <= credit_2 - 9'd1;
        end
        if(credit_from_chip[2] & ~(rdy_3 & val_3)) begin
            credit_3 <= credit_3 - 9'd1;
        end
        
        if((credit_1 < FULL_THRESHOLD) &&
           (credit_2 < FULL_THRESHOLD) &&
           (credit_3 < FULL_THRESHOLD) &&
           (sel_123 == 0)         )
            sel_123 <= 2'b01;
        
        if(rdy_1 & val_1) begin
            sel_13 <= 1;
            sel_12 <= 1;
            if (sel_123 == 2'b01) begin
                sel_123 <= 2'b10;
            end
            if(~credit_from_chip[0]) begin
                credit_1 <= credit_1 + 9'd1;
            end
        end 
        if(rdy_2 & val_2) begin
            sel_23 <= 1;
            sel_12 <= 0;
            if (sel_123 == 2'b10) begin
                sel_123 <= 2'b11;
            end
            if( ~credit_from_chip[1]) begin
                credit_2 <= credit_2 + 9'd1;
            end
        end
        if(rdy_3 & val_3) begin
            sel_23 <= 0;
            sel_13 <= 0;
            if (sel_123 == 2'b11) begin
                sel_123 <= 2'b01;
            end
            if (~credit_from_chip[2]) begin
                credit_3 <= credit_3 + 9'd1;
            end
        end
    end
end 
endmodule
module io_xbar_bus_compare_equal (a, b, bus_equal);
    parameter WIDTH = 8;
    parameter BHC = 10;
    input [WIDTH-1:0] a, b;
    output wire bus_equal;
    assign bus_equal = (a==b) ? 1'b1 : 1'b0;
endmodule
module io_xbar_flip_bus (in, out);
    parameter WIDTH = 8;
    parameter BHC = 10;
    input [WIDTH-1:0] in;
    output wire [WIDTH-1:0] out;
    
    assign out = ~in;
endmodule
module io_xbar_net_dff #(parameter WIDTH=8, parameter BHC=10) 
    (input wire [WIDTH-1:0] d, 
    output reg [WIDTH-1:0] q,
    input wire clk);
always @ (posedge clk)
begin
    q <= d;
end
endmodule
module io_xbar_one_of_n(
  
  in0,
  in1,
  in2,
  in3,
  in4,
  in5,
  sel,
  out);
    parameter WIDTH = 8;
    parameter BHC = 10;
    input [2:0] sel;
    input [WIDTH-1:0] in0,in1,in2,in3,in4,in5;
    output reg [WIDTH-1:0] out;
    always@(*)
    begin
        out={WIDTH{1'b0}};
        case(sel)
        
            3'd0:out=in0;
            3'd1:out=in1;
            3'd2:out=in2;
            3'd3:out=in3;
            3'd4:out=in4;
            3'd5:out=in5;
            default:; 
        endcase
    end
endmodule
module io_xbar_one_of_n_plus_3(
  
  in0,
  in1,
  in2,
  in3,
  in4,
  in5,
  in6,
  in7,
  in8,
  sel,
  out);
    parameter WIDTH = 8;
    parameter BHC = 10;
    input [3:0] sel;
    
    input [WIDTH-1:0] in0,in1,in2,in3,in4,in5,in6,in7,in8;
    output reg [WIDTH-1:0] out;
    always@(*)
    begin
        out={WIDTH{1'b0}};
        case(sel)
        
            4'd0:out=in0;
            4'd1:out=in1;
            4'd2:out=in2;
            4'd3:out=in3;
            4'd4:out=in4;
            4'd5:out=in5;
            4'd6:out=in6;
            4'd7:out=in7;
            4'd8:out=in8;
            default:; 
        endcase
    end
endmodule
 
 
 
 
 
 
 
module io_xbar_input_control(thanks_all_temp_out,
                             route_req_0_out, route_req_1_out, route_req_2_out, route_req_3_out, route_req_4_out, route_req_5_out, 
                             default_ready_0, default_ready_1, default_ready_2, default_ready_3, default_ready_4, default_ready_5, 
                             tail_out, clk, reset,
                             my_loc_x_in, my_loc_y_in, my_chip_id_in,
                             abs_x, abs_y, abs_chip_id, final_bits, valid_in,
                             thanks_0, thanks_1, thanks_2, thanks_3, thanks_4, thanks_5, 
                             length);
output thanks_all_temp_out;
output route_req_0_out;
output route_req_1_out;
output route_req_2_out;
output route_req_3_out;
output route_req_4_out;
output route_req_5_out;
output default_ready_0;
output default_ready_1;
output default_ready_2;
output default_ready_3;
output default_ready_4;
output default_ready_5;
output tail_out;
input clk;
input reset;
input [8-1:0] my_loc_x_in;
input [8-1:0] my_loc_y_in;
input [14-1:0] my_chip_id_in;
input [8-1:0] abs_x;
input [8-1:0] abs_y;
input [14-1:0] abs_chip_id;
input [2:0] final_bits;
input valid_in;
input thanks_0;
input thanks_1;
input thanks_2;
input thanks_3;
input thanks_4;
input thanks_5;
input [8-1:0] length;
reg [8-1:0] count_f;
reg header_last_f;
reg thanks_all_f;
reg count_zero_f;
reg count_one_f;
reg tail_last_f;
reg [8-1:0] count_temp;
wire header_last_temp;
wire thanks_all_temp;
wire count_zero_temp;
wire count_one_temp;
wire tail_last_temp;
wire header;
wire [8-1:0] count_minus_one;
wire length_zero; 
                  
wire tail;
reg header_temp;
assign thanks_all_temp = thanks_0 | thanks_1 | thanks_2 | thanks_3 | thanks_4 | thanks_5;
assign header = valid_in & header_temp;
assign count_zero_temp = count_temp == 0;
assign count_one_temp = count_temp == 1;
assign thanks_all_temp_out = thanks_all_temp;
assign tail_out = tail;
assign count_minus_one = count_f - 1;
assign length_zero = length == 0;
assign header_last_temp = header_temp;
assign tail = (header & length_zero) | ((~thanks_all_f) & tail_last_f) | (thanks_all_f & count_one_f);
assign tail_last_temp = tail;
io_xbar_route_request_calc tail_calc(.route_req_0(route_req_0_out),
                                           .route_req_1(route_req_1_out),
                                           .route_req_2(route_req_2_out),
                                           .route_req_3(route_req_3_out),
                                           .route_req_4(route_req_4_out),
                                           .route_req_5(route_req_5_out),
                                           .default_ready_0(default_ready_0),
                                           .default_ready_1(default_ready_1),
                                           .default_ready_2(default_ready_2),
                                           .default_ready_3(default_ready_3),
                                           .default_ready_4(default_ready_4),
                                           .default_ready_5(default_ready_5),
                                           .my_loc_x_in(my_loc_x_in),
                                           .my_loc_y_in(my_loc_y_in),
                                           .my_chip_id_in(my_chip_id_in),
                                           .abs_x(abs_x),
                                           .abs_y(abs_y),
                                           .abs_chip_id(abs_chip_id),
                                           .final_bits(final_bits),
                                           .length(length),
                                           .header_in(header));
always @ (header_last_f or thanks_all_f or count_zero_f)
begin
        case({header_last_f, count_zero_f, thanks_all_f})
        3'b000: header_temp <= 1'b0;
        3'b001: header_temp <= 1'b0;
        3'b010: header_temp <= 1'b0;
        3'b011: header_temp <= 1'b1;
        3'b100: header_temp <= 1'b1;
        
        3'b101: header_temp <= 1'b0;
        3'b110: header_temp <= 1'b1;
        3'b111: header_temp <= 1'b1;
        default:
                header_temp <= 1'b1;
        endcase
end
always @ (header or thanks_all_f or count_f or count_minus_one or length)
begin
        if(header)
        begin
                count_temp <= length;
        end
        else
        begin
                if(thanks_all_f)
                begin
                        count_temp <= count_minus_one;
                end
                else
                begin
                        count_temp <= count_f;
                end
        end
end
always @ (posedge clk)
begin
        if(reset)
        begin
                count_f <= 5'd0;
                header_last_f <= 1'b1;
                thanks_all_f <= 1'b0;
                count_zero_f <= 1'b1; 
                count_one_f <= 1'b0;
                tail_last_f <= 1'b0;
        end
        else
        begin
                count_f <= count_temp;
                header_last_f <= header_last_temp;
                thanks_all_f <= thanks_all_temp;
                count_zero_f <= count_zero_temp;
                count_one_f <= count_one_temp;
                tail_last_f <= tail_last_temp;
        end
end
endmodule
 
 
 
 
 
 
 
module io_xbar_route_request_calc(route_req_0, route_req_1, route_req_2, route_req_3, route_req_4, route_req_5, 
                                        default_ready_0, default_ready_1, default_ready_2, default_ready_3, default_ready_4, default_ready_5, 
                                        my_loc_x_in, my_loc_y_in, my_chip_id_in, abs_x, abs_y, abs_chip_id, final_bits, length, header_in);
output route_req_0;
output route_req_1;
output route_req_2;
output route_req_3;
output route_req_4;
output route_req_5;
output default_ready_0;
output default_ready_1;
output default_ready_2;
output default_ready_3;
output default_ready_4;
output default_ready_5;
input [8-1:0] my_loc_x_in;
input [8-1:0] my_loc_y_in;
input [14-1:0] my_chip_id_in;
input [8-1:0] abs_x;
input [8-1:0] abs_y;
input [14-1:0] abs_chip_id;
input [2:0] final_bits;
input [8-1:0] length;
input header_in;
wire off_chip;
wire [8*3+3-1:0]              stub;
assign off_chip = abs_chip_id != my_chip_id_in;
assign route_req_1 = header_in & (!off_chip) & (abs_x == 8'd1);
assign route_req_2 = header_in & (!off_chip) & (abs_x == 8'd2);
assign route_req_3 = header_in & (!off_chip) & (abs_x == 8'd3);
assign route_req_4 = header_in & (!off_chip) & (abs_x == 8'd4);
assign route_req_5 = header_in & (!off_chip) & (abs_x == 8'd5);
assign route_req_0 = (header_in & (!off_chip) & (abs_x == 8'd0)) | (header_in & (off_chip)) ;
assign default_ready_0 = route_req_0;
assign default_ready_1 = route_req_1;
assign default_ready_2 = route_req_2;
assign default_ready_3 = route_req_3;
assign default_ready_4 = route_req_4;
assign default_ready_5 = route_req_5;
assign stub = {my_loc_x_in, my_loc_y_in, abs_y, final_bits};
endmodule
   
 
 
 
 
 
 
 
module io_xbar_input_top_16(route_req_0_out, route_req_1_out, route_req_2_out, route_req_3_out, route_req_4_out, route_req_5_out, default_ready_0_out, default_ready_1_out, default_ready_2_out, default_ready_3_out, default_ready_4_out, default_ready_5_out, tail_out, yummy_out, data_out, valid_out, clk, reset, my_loc_x_in, my_loc_y_in, my_chip_id_in, valid_in, data_in,thanks_0, thanks_1, thanks_2, thanks_3, thanks_4, thanks_5);
output route_req_0_out;
output route_req_1_out;
output route_req_2_out;
output route_req_3_out;
output route_req_4_out;
output route_req_5_out;
output default_ready_0_out;
output default_ready_1_out;
output default_ready_2_out;
output default_ready_3_out;
output default_ready_4_out;
output default_ready_5_out;
output tail_out;
output yummy_out;
output [64-1:0] data_out;
output valid_out;
input clk;
input reset;
input [8-1:0] my_loc_x_in;
input [8-1:0] my_loc_y_in;
input [14-1:0] my_chip_id_in;
input valid_in;
input [64-1:0] data_in;
input thanks_0;
input thanks_1;
input thanks_2;
input thanks_3;
input thanks_4;
input thanks_5;
   
wire thanks_all_temp;
wire valid_out_internal;
wire [64-1:0] data_out_internal;
wire [64-1:0] data_out_internal_pre;
assign valid_out = valid_out_internal;
assign data_out = data_out_internal;
network_input_blk_multi_out #(.LOG2_NUMBER_FIFO_ELEMENTS(4)) NIB(.clk(clk), .reset(reset), .data_in(data_in), .valid_in(valid_in), .yummy_out(yummy_out), .thanks_in(thanks_all_temp), .data_val(data_out_internal_pre), .data_val1(), .data_avail(valid_out_internal));
assign data_out_internal = data_out_internal_pre;
io_xbar_input_control control(.thanks_all_temp_out(thanks_all_temp), .route_req_0_out(route_req_0_out), .route_req_1_out(route_req_1_out), .route_req_2_out(route_req_2_out), .route_req_3_out(route_req_3_out), .route_req_4_out(route_req_4_out), .route_req_5_out(route_req_5_out), .default_ready_0(default_ready_0_out), .default_ready_1(default_ready_1_out), .default_ready_2(default_ready_2_out), .default_ready_3(default_ready_3_out), .default_ready_4(default_ready_4_out), .default_ready_5(default_ready_5_out), .tail_out(tail_out), .clk(clk), .reset(reset), .my_loc_x_in(my_loc_x_in), .my_loc_y_in(my_loc_y_in), 
    .my_chip_id_in(my_chip_id_in), .abs_x(data_out_internal[64-14-1:64-14-8]), .abs_y(data_out_internal[64-14-8-1:64-14-2*8]), .abs_chip_id(data_out_internal[64-1:64-14]),.final_bits(data_out_internal[64-14-2*8-2:64-14-2*8-4]), .valid_in(valid_out_internal), .thanks_0(thanks_0), .thanks_1(thanks_1), .thanks_2(thanks_2), .thanks_3(thanks_3), .thanks_4(thanks_4), .thanks_5(thanks_5), .length(data_out_internal[64-14-2*8-5:64-14-2*8-4-8]));
endmodule
 
 
 
 
 
 
 
module io_xbar_input_top_4(route_req_0_out, route_req_1_out, route_req_2_out, route_req_3_out, route_req_4_out, route_req_5_out, 
                           default_ready_0_out, default_ready_1_out, default_ready_2_out, default_ready_3_out, default_ready_4_out, default_ready_5_out, 
                           tail_out, yummy_out, data_out, valid_out, clk, reset,
                           my_loc_x_in, my_loc_y_in, my_chip_id_in,  valid_in, data_in,
                           thanks_0, thanks_1, thanks_2, thanks_3, thanks_4, thanks_5);
output route_req_0_out;
output route_req_1_out;
output route_req_2_out;
output route_req_3_out;
output route_req_4_out;
output route_req_5_out;
output default_ready_0_out;
output default_ready_1_out;
output default_ready_2_out;
output default_ready_3_out;
output default_ready_4_out;
output default_ready_5_out;
output tail_out;
output yummy_out;
output [64-1:0] data_out;
output valid_out;
input clk;
input reset;
input [8-1:0] my_loc_x_in;
input [8-1:0] my_loc_y_in;
input [14-1:0] my_chip_id_in;
input valid_in;
input [64-1:0] data_in;
input thanks_0;
input thanks_1;
input thanks_2;
input thanks_3;
input thanks_4;
input thanks_5;
wire thanks_all_temp;
wire [64-1:0] data_internal;
wire valid_out_internal;
assign valid_out = valid_out_internal;
network_input_blk_multi_out #(.LOG2_NUMBER_FIFO_ELEMENTS(2)) NIB(.clk(clk),
                                      .reset(reset),
                                      .data_in(data_in),
                                      .valid_in(valid_in),
                                      .yummy_out(yummy_out),
                                      .thanks_in(thanks_all_temp),
                                      .data_val(data_out),
                                      .data_val1(data_internal), 
                                      .data_avail(valid_out_internal));
io_xbar_input_control control(.thanks_all_temp_out(thanks_all_temp),
                              .route_req_0_out(route_req_0_out), .route_req_1_out(route_req_1_out), .route_req_2_out(route_req_2_out), .route_req_3_out(route_req_3_out), .route_req_4_out(route_req_4_out), .route_req_5_out(route_req_5_out), 
                              .default_ready_0(default_ready_0_out), .default_ready_1(default_ready_1_out), .default_ready_2(default_ready_2_out), .default_ready_3(default_ready_3_out), .default_ready_4(default_ready_4_out), .default_ready_5(default_ready_5_out), 
                              .tail_out(tail_out),
                              .clk(clk), .reset(reset),
                              .my_loc_x_in(my_loc_x_in), 
                              .my_loc_y_in(my_loc_y_in), 
                              .my_chip_id_in(my_chip_id_in),
                              .abs_x(data_internal[64-14-1:64-14-8]), 
                              .abs_y(data_internal[64-14-8-1:64-14-2*8]), 
                              .abs_chip_id(data_internal[64-1:64-14]),
                              .final_bits(data_internal[64-14-2*8-2:64-14-2*8-4]),
                              .valid_in(valid_out_internal),
                              .thanks_0(thanks_0), .thanks_1(thanks_1), .thanks_2(thanks_2), .thanks_3(thanks_3), .thanks_4(thanks_4), .thanks_5(thanks_5), 
                              .length(data_internal[64-14-2*8-5:64-14-2*8-4-8]));
endmodule
 
 
 
 
 
 
 
module io_xbar_output_control(thanks_0, thanks_1, thanks_2, thanks_3, thanks_4, thanks_5, 
                              valid_out, current_route, ec_wants_to_send_but_cannot, clk, reset, 
                              route_req_0_in, route_req_1_in, route_req_2_in, route_req_3_in, route_req_4_in, route_req_5_in, 
                              tail_0_in, tail_1_in, tail_2_in, tail_3_in, tail_4_in, tail_5_in, 
                              valid_out_temp, default_ready, space_avail);
output thanks_0;
output thanks_1;
output thanks_2;
output thanks_3;
output thanks_4;
output thanks_5;
output valid_out;
output [2:0] current_route;
output    ec_wants_to_send_but_cannot;
input clk;
input reset;
input route_req_0_in;
input route_req_1_in;
input route_req_2_in;
input route_req_3_in;
input route_req_4_in;
input route_req_5_in;
input tail_0_in;
input tail_1_in;
input tail_2_in;
input tail_3_in;
input tail_4_in;
input tail_5_in;
input valid_out_temp;
input default_ready;
input space_avail;
reg [2:0]current_route_f;
reg planned_f;
wire [2:0] current_route_temp;
wire planned_or_default;
wire route_req_all_or_with_planned;
wire route_req_all_but_default;
wire valid_out_internal;
reg new_route_needed;
reg planned_temp;
reg [2:0] new_route;
reg tail_current_route;
reg route_req_0_mask;
reg route_req_1_mask;
reg route_req_2_mask;
reg route_req_3_mask;
reg route_req_4_mask;
reg route_req_5_mask;
reg thanks_0;
reg thanks_1;
reg thanks_2;
reg thanks_3;
reg thanks_4;
reg thanks_5;
reg    ec_wants_to_send_but_cannot;
assign planned_or_default = planned_f | default_ready;
assign valid_out_internal = valid_out_temp & planned_or_default & space_avail;
always @(posedge clk)
  begin
     ec_wants_to_send_but_cannot <= valid_out_temp & planned_or_default & ~space_avail;
  end
assign current_route_temp = (new_route_needed) ? new_route : current_route_f;
assign current_route = current_route_f;
assign route_req_all_or_with_planned = (route_req_0_in & route_req_0_mask) | (route_req_1_in & route_req_1_mask) | (route_req_2_in & route_req_2_mask) | (route_req_3_in & route_req_3_mask) | (route_req_4_in & route_req_4_mask) | (route_req_5_in & route_req_5_mask);
assign route_req_all_but_default = (route_req_1_in) | (route_req_2_in) | (route_req_3_in) | (route_req_4_in) | (route_req_5_in);
assign valid_out = valid_out_internal;
always @ (current_route_f or tail_0_in or tail_1_in or tail_2_in or tail_3_in or tail_4_in or tail_5_in)
begin
	case(current_route_f) 
	
	3'b000:
	begin
		tail_current_route <= tail_0_in;
	end
	3'b001:
	begin
		tail_current_route <= tail_1_in;
	end
	3'b010:
	begin
		tail_current_route <= tail_2_in;
	end
	3'b011:
	begin
		tail_current_route <= tail_3_in;
	end
	3'b100:
	begin
		tail_current_route <= tail_4_in;
	end
	3'b101:
	begin
		tail_current_route <= tail_5_in;
	end
	default:
	begin
		tail_current_route <= 1'bx; 
					    
					    
					    
					    
	end
	endcase
end
always @ (current_route_f or valid_out_internal)
begin
	case(current_route_f)
	
	
	3'b000:
	begin
		thanks_0 <= valid_out_internal;
		thanks_1 <= 1'b0;
		thanks_2 <= 1'b0;
		thanks_3 <= 1'b0;
		thanks_4 <= 1'b0;
		thanks_5 <= 1'b0;
	end
	3'b001:
	begin
		thanks_0 <= 1'b0;
		thanks_1 <= valid_out_internal;
		thanks_2 <= 1'b0;
		thanks_3 <= 1'b0;
		thanks_4 <= 1'b0;
		thanks_5 <= 1'b0;
	end
	3'b010:
	begin
		thanks_0 <= 1'b0;
		thanks_1 <= 1'b0;
		thanks_2 <= valid_out_internal;
		thanks_3 <= 1'b0;
		thanks_4 <= 1'b0;
		thanks_5 <= 1'b0;
	end
	3'b011:
	begin
		thanks_0 <= 1'b0;
		thanks_1 <= 1'b0;
		thanks_2 <= 1'b0;
		thanks_3 <= valid_out_internal;
		thanks_4 <= 1'b0;
		thanks_5 <= 1'b0;
	end
	3'b100:
	begin
		thanks_0 <= 1'b0;
		thanks_1 <= 1'b0;
		thanks_2 <= 1'b0;
		thanks_3 <= 1'b0;
		thanks_4 <= valid_out_internal;
		thanks_5 <= 1'b0;
	end
	3'b101:
	begin
		thanks_0 <= 1'b0;
		thanks_1 <= 1'b0;
		thanks_2 <= 1'b0;
		thanks_3 <= 1'b0;
		thanks_4 <= 1'b0;
		thanks_5 <= valid_out_internal;
	end
	default:
	begin
	
		thanks_0 <= 1'bx;
		thanks_1 <= 1'bx;
		thanks_2 <= 1'bx;
		thanks_3 <= 1'bx;
		thanks_4 <= 1'bx;
		thanks_5 <= 1'bx;
	
					
					
					
	end
	endcase
end
always @(current_route_f or route_req_0_in or route_req_1_in or route_req_2_in or route_req_3_in or route_req_4_in or route_req_5_in)
begin
	case(current_route_f)
	
	
	3'b000:
	begin
		new_route <= (route_req_1_in)?3'b001:((route_req_2_in)?3'b010:((route_req_3_in)?3'b011:((route_req_4_in)?3'b100:((route_req_5_in)?3'b101:3'b000))));
	end
	3'b001:
	begin
		new_route <= (route_req_2_in)?3'b010:((route_req_3_in)?3'b011:((route_req_4_in)?3'b100:((route_req_5_in)?3'b101:((route_req_0_in)?3'b000:3'b000))));
	end
	3'b010:
	begin
		new_route <= (route_req_3_in)?3'b011:((route_req_4_in)?3'b100:((route_req_5_in)?3'b101:((route_req_0_in)?3'b000:((route_req_1_in)?3'b001:3'b000))));
	end
	3'b011:
	begin
		new_route <= (route_req_4_in)?3'b100:((route_req_5_in)?3'b101:((route_req_0_in)?3'b000:((route_req_1_in)?3'b001:((route_req_2_in)?3'b010:3'b000))));
	end
	3'b100:
	begin
		new_route <= (route_req_5_in)?3'b101:((route_req_0_in)?3'b000:((route_req_1_in)?3'b001:((route_req_2_in)?3'b010:((route_req_3_in)?3'b011:3'b000))));
	end
	3'b101:
	begin
		new_route <= (route_req_0_in)?3'b000:((route_req_1_in)?3'b001:((route_req_2_in)?3'b010:((route_req_3_in)?3'b011:((route_req_4_in)?3'b100:3'b000))));
	end
	default:
	begin
		new_route <= 3'b000;
			
	end
	endcase
end
always @(current_route_f or planned_f)
begin
	if(planned_f)
	begin
		case(current_route_f)
		
		3'b000:
			begin
				route_req_0_mask <= 1'b0;
				route_req_1_mask <= 1'b1;
				route_req_2_mask <= 1'b1;
				route_req_3_mask <= 1'b1;
				route_req_4_mask <= 1'b1;
				route_req_5_mask <= 1'b1;
			end
		3'b001:
			begin
				route_req_0_mask <= 1'b1;
				route_req_1_mask <= 1'b0;
				route_req_2_mask <= 1'b1;
				route_req_3_mask <= 1'b1;
				route_req_4_mask <= 1'b1;
				route_req_5_mask <= 1'b1;
			end
		3'b010:
			begin
				route_req_0_mask <= 1'b1;
				route_req_1_mask <= 1'b1;
				route_req_2_mask <= 1'b0;
				route_req_3_mask <= 1'b1;
				route_req_4_mask <= 1'b1;
				route_req_5_mask <= 1'b1;
			end
		3'b011:
			begin
				route_req_0_mask <= 1'b1;
				route_req_1_mask <= 1'b1;
				route_req_2_mask <= 1'b1;
				route_req_3_mask <= 1'b0;
				route_req_4_mask <= 1'b1;
				route_req_5_mask <= 1'b1;
			end
		3'b100:
			begin
				route_req_0_mask <= 1'b1;
				route_req_1_mask <= 1'b1;
				route_req_2_mask <= 1'b1;
				route_req_3_mask <= 1'b1;
				route_req_4_mask <= 1'b0;
				route_req_5_mask <= 1'b1;
			end
		3'b101:
			begin
				route_req_0_mask <= 1'b1;
				route_req_1_mask <= 1'b1;
				route_req_2_mask <= 1'b1;
				route_req_3_mask <= 1'b1;
				route_req_4_mask <= 1'b1;
				route_req_5_mask <= 1'b0;
			end
		default:
			begin
				route_req_0_mask <= 1'b1;
				route_req_1_mask <= 1'b1;
				route_req_2_mask <= 1'b1;
				route_req_3_mask <= 1'b1;
				route_req_4_mask <= 1'b1;
				route_req_5_mask <= 1'b1;
			end
		
		endcase
	end
	else
	begin
	
		route_req_0_mask <= 1'b1;
		route_req_1_mask <= 1'b1;
		route_req_2_mask <= 1'b1;
		route_req_3_mask <= 1'b1;
		route_req_4_mask <= 1'b1;
		route_req_5_mask <= 1'b1;
	
	end
end
always @ (planned_f or tail_current_route or valid_out_internal or default_ready)
begin
	case({default_ready, valid_out_internal, tail_current_route, planned_f}) 
	4'b0000:	new_route_needed <= 1'b1;
	4'b0001:	new_route_needed <= 1'b0;
	4'b0010:	new_route_needed <= 1'b1;
	4'b0011:	new_route_needed <= 1'b0;
	4'b0100:	new_route_needed <= 1'b0;	
	4'b0101:	new_route_needed <= 1'b0;	
	4'b0110:	new_route_needed <= 1'b1;
	4'b0111:	new_route_needed <= 1'b1;
	4'b1000:	new_route_needed <= 1'b1;
	4'b1001:	new_route_needed <= 1'b0;
	4'b1010:	new_route_needed <= 1'b1;	
    
	4'b1011:	new_route_needed <= 1'b0;
	4'b1100:	new_route_needed <= 1'b0;
	4'b1101:	new_route_needed <= 1'b0;
	4'b1110:	new_route_needed <= 1'b1;
	4'b1111:	new_route_needed <= 1'b1;
	default:	new_route_needed <= 1'b1;
			
	endcase
end
always @ (planned_f or tail_current_route or valid_out_internal or default_ready or route_req_all_or_with_planned or route_req_all_but_default)
begin
	case({route_req_all_or_with_planned, default_ready, valid_out_internal, tail_current_route, planned_f}) 
	5'b00000:	planned_temp <= 1'b0;
	5'b00001:	planned_temp <= 1'b1;
	5'b00010:	planned_temp <= 1'b0;
	5'b00011:	planned_temp <= 1'b1;
	5'b00100:	planned_temp <= 1'b0;	
	5'b00101:	planned_temp <= 1'b1;
	5'b00110:	planned_temp <= 1'b0;	
	5'b00111:	planned_temp <= 1'b0;
	5'b01000:	planned_temp <= 1'b0;	
	5'b01001:	planned_temp <= 1'b1;
	5'b01010:	planned_temp <= 1'b0;	
	5'b01011:	planned_temp <= 1'b1;
	5'b01100:	planned_temp <= 1'b0;	
	5'b01101:	planned_temp <= 1'b1;
	5'b01110:	planned_temp <= 1'b0;	
	5'b01111:	planned_temp <= 1'b0;	
						
						
						
						
						
	5'b10000:	planned_temp <= 1'b1;
	5'b10001:	planned_temp <= 1'b1;
	5'b10010:	planned_temp <= 1'b1;
	5'b10011:	planned_temp <= 1'b1;
	5'b10100:	planned_temp <= 1'b1;
	5'b10101:	planned_temp <= 1'b1;
	5'b10110:	planned_temp <= 1'b1;
	5'b10111:	planned_temp <= 1'b1;
	5'b11000:	planned_temp <= 1'b1;
	5'b11001:	planned_temp <= 1'b1;
	5'b11010:	planned_temp <= 1'b1;
	5'b11011:	planned_temp <= 1'b1;
	5'b11100:	planned_temp <= 1'b1;
	5'b11101:	planned_temp <= 1'b1;
						
						
						
						
						
	5'b11110:	planned_temp <= route_req_all_but_default;
	5'b11111:	planned_temp <= 1'b1;
	default:	planned_temp <= 1'b0;
	endcase
end
always @(posedge clk)
begin
	if(reset)
	begin
		current_route_f <= 3'd0;
		planned_f <= 1'd0;
	end
	else
	begin
		current_route_f <= current_route_temp;
		planned_f <= planned_temp;
	end
end
endmodule
 
 
 
 
 
 
 
module io_xbar_output_datapath(data_out, valid_out_temp, data_0_in, data_1_in, data_2_in, data_3_in, data_4_in, data_5_in, valid_0_in, valid_1_in, valid_2_in, valid_3_in, valid_4_in, valid_5_in, current_route_in);
output [64-1:0] data_out;
output valid_out_temp;
input [64-1:0] data_0_in;
input [64-1:0] data_1_in;
input [64-1:0] data_2_in;
input [64-1:0] data_3_in;
input [64-1:0] data_4_in;
input [64-1:0] data_5_in;
input valid_0_in;
input valid_1_in;
input valid_2_in;
input valid_3_in;
input valid_4_in;
input valid_5_in;
input [2:0] current_route_in;
io_xbar_one_of_n #(64) data_mux(.in0(data_0_in), .in1(data_1_in), .in2(data_2_in), .in3(data_3_in), .in4(data_4_in), .in5(data_5_in), .sel(current_route_in), .out(data_out));
io_xbar_one_of_n #(1) valid_mux(.in0(valid_0_in), .in1(valid_1_in), .in2(valid_2_in), .in3(valid_3_in), .in4(valid_4_in), .in5(valid_5_in), .sel(current_route_in), .out(valid_out_temp));
endmodule
 
 
 
 
 
 
 
module io_xbar_output_top(data_out, 
                          thanks_0_out, thanks_1_out, thanks_2_out, thanks_3_out, thanks_4_out, thanks_5_out, 
                          valid_out, popped_interrupt_mesg_out, popped_memory_ack_mesg_out, popped_memory_ack_mesg_out_sender, ec_wants_to_send_but_cannot, clk, reset, 
                          route_req_0_in, route_req_1_in, route_req_2_in, route_req_3_in, route_req_4_in, route_req_5_in, 
                          tail_0_in, tail_1_in, tail_2_in, tail_3_in, tail_4_in, tail_5_in, 
                          data_0_in, data_1_in, data_2_in, data_3_in, data_4_in, data_5_in, 
                          valid_0_in, valid_1_in, valid_2_in, valid_3_in, valid_4_in, valid_5_in, 
                          default_ready_in, yummy_in);
parameter KILL_HEADERS = 1'b0;
output [64-1:0] data_out;
output thanks_0_out;
output thanks_1_out;
output thanks_2_out;
output thanks_3_out;
output thanks_4_out;
output thanks_5_out;
output valid_out;
output popped_interrupt_mesg_out;
output popped_memory_ack_mesg_out;
output [9:0] popped_memory_ack_mesg_out_sender;
output ec_wants_to_send_but_cannot;
input clk;
input reset;
input route_req_0_in;
input route_req_1_in;
input route_req_2_in;
input route_req_3_in;
input route_req_4_in;
input route_req_5_in;
input tail_0_in;
input tail_1_in;
input tail_2_in;
input tail_3_in;
input tail_4_in;
input tail_5_in;
input [64-1:0] data_0_in;
input [64-1:0] data_1_in;
input [64-1:0] data_2_in;
input [64-1:0] data_3_in;
input [64-1:0] data_4_in;
input [64-1:0] data_5_in;
input valid_0_in;
input valid_1_in;
input valid_2_in;
input valid_3_in;
input valid_4_in;
input valid_5_in;
input default_ready_in;
input yummy_in;
wire valid_out_temp_connection;
wire [2:0] current_route_connection;
wire space_avail_connection;
wire valid_out_pre;
wire data_out_len_zero;
wire data_out_interrupt_user_bits_set;
wire data_out_memory_ack_user_bits_set;
wire [64-1:0] data_out_internal;
wire valid_out_internal;
reg current_route_req;
assign valid_out_internal = valid_out_pre & ~(KILL_HEADERS & current_route_req);
assign data_out_len_zero = data_out_internal[64-14-2*8-4:64-14-2*8-3-8] == 8'd0;
assign data_out_interrupt_user_bits_set = data_out_internal[23:20] == 4'b1111;
assign data_out_memory_ack_user_bits_set = data_out_internal[23:20] == 4'b1110;
assign popped_interrupt_mesg_out = data_out_interrupt_user_bits_set & data_out_len_zero & valid_out_pre & (KILL_HEADERS & current_route_req);
assign popped_memory_ack_mesg_out = data_out_memory_ack_user_bits_set & data_out_len_zero & valid_out_pre & (KILL_HEADERS & current_route_req);
assign popped_memory_ack_mesg_out_sender = data_out_internal[19:10] & { 10 { KILL_HEADERS} };
assign data_out = data_out_internal;
assign valid_out = valid_out_internal;
io_xbar_space_avail_top space(.valid(valid_out_internal), .clk(clk), .reset(reset), .yummy(yummy_in),.spc_avail(space_avail_connection));
io_xbar_output_datapath datapath(.data_out(data_out_internal), .valid_out_temp(valid_out_temp_connection), .data_0_in(data_0_in), .data_1_in(data_1_in), .data_2_in(data_2_in), .data_3_in(data_3_in), .data_4_in(data_4_in), .data_5_in(data_5_in), .valid_0_in(valid_0_in), .valid_1_in(valid_1_in), .valid_2_in(valid_2_in), .valid_3_in(valid_3_in), .valid_4_in(valid_4_in), .valid_5_in(valid_5_in), .current_route_in(current_route_connection));
io_xbar_output_control control(.thanks_0(thanks_0_out), .thanks_1(thanks_1_out), .thanks_2(thanks_2_out), .thanks_3(thanks_3_out), .thanks_4(thanks_4_out), .thanks_5(thanks_5_out), 
                               .valid_out(valid_out_pre), .current_route(current_route_connection), .ec_wants_to_send_but_cannot(ec_wants_to_send_but_cannot), .clk(clk), .reset(reset), 
                               .route_req_0_in(route_req_0_in), .route_req_1_in(route_req_1_in), .route_req_2_in(route_req_2_in), .route_req_3_in(route_req_3_in), .route_req_4_in(route_req_4_in), .route_req_5_in(route_req_5_in), 
                               .tail_0_in(tail_0_in), .tail_1_in(tail_1_in), .tail_2_in(tail_2_in), .tail_3_in(tail_3_in), .tail_4_in(tail_4_in), .tail_5_in(tail_5_in), 
                               .valid_out_temp(valid_out_temp_connection), .default_ready(default_ready_in), .space_avail(space_avail_connection));
always @ (current_route_connection or route_req_0_in or route_req_1_in or route_req_2_in or route_req_3_in or route_req_4_in or route_req_5_in)
begin
	case(current_route_connection)
    
	3'b000:    current_route_req <= route_req_0_in;
	3'b001:    current_route_req <= route_req_1_in;
	3'b010:    current_route_req <= route_req_2_in;
	3'b011:    current_route_req <= route_req_3_in;
	3'b100:    current_route_req <= route_req_4_in;
	3'b101:    current_route_req <= route_req_5_in;
    
	default:	current_route_req <= 1'bx;
	endcase
end
endmodule
module clk_gating_latch (
    input wire clk,
    input wire clk_en,
    output wire clk_out
);
 
  wire clk_en_sync;
  reg clk_en_sync_latch;
  assign clk_out = clk & clk_en_sync_latch;
  synchronizer sync(
      .clk            (clk),
      .presyncdata    (clk_en),
      .syncdata       (clk_en_sync)
  );
  
  
  always @ (clk or clk_en_sync)
      if (~clk) clk_en_sync_latch = clk_en_sync;
endmodule 
 
 
 
 
 
 
 
module credit_to_valrdy (
   clk,
   reset,
   
   data_in,
   valid_in,
   yummy_in,
            
   
   data_out,
   valid_out,
   ready_out
);
   input	 clk;
   input	 reset;
   input [64-1:0]	 data_in;
   input	 valid_in;
   input     ready_out;
    
   output	 yummy_in;
   output	 valid_out;
   output [64-1:0] data_out;
   
   wire	 thanksIn;
   wire valid_out_temp;
   assign valid_out = valid_out_temp;
   network_input_blk_multi_out #(.LOG2_NUMBER_FIFO_ELEMENTS(2)) data(
      .clk(clk),
      .reset(reset),
      .data_in(data_in),
      .valid_in(valid_in),
      .thanks_in(valid_out & ready_out),
      .yummy_out(yummy_in),
      .data_val(data_out),
      .data_val1(),
      .data_avail(valid_out_temp));
endmodule
module zznor64_32 ( znor64, znor32, a );
  input  [63:0] a;
  output        znor64;
  output        znor32;
  assign znor32 =  ~(a[0]  | a[1]  | a[2]  | a[3]  | a[4]  | a[5]  | a[6]  | a[7]
		   | a[8]  | a[9]  | a[10] | a[11] | a[12] | a[13] | a[14] | a[15]
		   | a[16] | a[17] | a[18] | a[19] | a[20] | a[21] | a[22] | a[23]
		   | a[24] | a[25] | a[26] | a[27] | a[28] | a[29] | a[30] | a[31]); 
  assign znor64 =  ~(a[0]  | a[1]  | a[2]  | a[3]  | a[4]  | a[5]  | a[6]  | a[7]
		   | a[8]  | a[9]  | a[10] | a[11] | a[12] | a[13] | a[14] | a[15]
		   | a[16] | a[17] | a[18] | a[19] | a[20] | a[21] | a[22] | a[23]
		   | a[24] | a[25] | a[26] | a[27] | a[28] | a[29] | a[30] | a[31] 
		   | a[32] | a[33] | a[34] | a[35] | a[36] | a[37] | a[38] | a[39] 
		   | a[40] | a[41] | a[42] | a[43] | a[44] | a[45] | a[46] | a[47] 
		   | a[48] | a[49] | a[50] | a[51] | a[52] | a[53] | a[54] | a[55] 
		   | a[56] | a[57] | a[58] | a[59] | a[60] | a[61] | a[62] | a[63]);
endmodule 
module zzor36 ( z, a );
  input  [35:0] a;
  output        z;
  assign z =  (a[0]  | a[1]  | a[2]  | a[3]  | a[4]  | a[5]  | a[6]  | a[7]
	     | a[8]  | a[9]  | a[10] | a[11] | a[12] | a[13] | a[14] | a[15]
	     | a[16] | a[17] | a[18] | a[19] | a[20] | a[21] | a[22] | a[23]
	     | a[24] | a[25] | a[26] | a[27] | a[28] | a[29] | a[30] | a[31]
	     | a[32] | a[33] | a[34] | a[35]); 
   
endmodule 
module zzor32 ( z, a );
  input  [31:0] a;
  output        z;
  assign z =  (a[0]  | a[1]  | a[2]  | a[3]  | a[4]  | a[5]  | a[6]  | a[7]
	     | a[8]  | a[9]  | a[10] | a[11] | a[12] | a[13] | a[14] | a[15]
	     | a[16] | a[17] | a[18] | a[19] | a[20] | a[21] | a[22] | a[23]
	     | a[24] | a[25] | a[26] | a[27] | a[28] | a[29] | a[30] | a[31]); 
endmodule 
module zznor24 ( z, a );
  input  [23:0] a;
  output        z;
  assign z =  ~(a[0]  | a[1]  | a[2]  | a[3]  | a[4]  | a[5]  | a[6]  | a[7]
	      | a[8]  | a[9]  | a[10] | a[11] | a[12] | a[13] | a[14] | a[15]
	      | a[16] | a[17] | a[18] | a[19] | a[20] | a[21] | a[22] | a[23]); 
endmodule 
module zznor16 ( z, a );
  input  [15:0] a;
  output        z;
  assign z =  ~(a[0] | a[1] | a[2]  | a[3]  | a[4]  | a[5]  | a[6]  | a[7]
	      | a[8] | a[9] | a[10] | a[11] | a[12] | a[13] | a[14] | a[15]); 
endmodule 
module zzor8 ( z, a );
  input  [7:0] a;
  output       z;
  assign z =  (a[0] | a[1] | a[2] | a[3] | a[4] | a[5] | a[6] | a[7]); 
   
endmodule 
module zzadd13 ( rs1_data, rs2_data, cin, adder_out );
  input  [12:0] rs1_data;   
  input  [12:0] rs2_data;   
  input         cin;        
  output [12:0] adder_out;  
  assign adder_out = rs1_data + rs2_data + cin;
endmodule 
module zzadd56 ( rs1_data, rs2_data, cin, adder_out );
  input  [55:0] rs1_data;   
  input  [55:0] rs2_data;   
  input         cin;        
  output [55:0] adder_out;  
  assign adder_out = rs1_data + rs2_data + cin;
endmodule 
module zzadd48 ( rs1_data, rs2_data, cin, adder_out );
  input  [47:0] rs1_data;   
  input  [47:0] rs2_data;   
  input         cin;        
  output [47:0] adder_out;  
  assign adder_out = rs1_data + rs2_data + cin;
endmodule 
module zzadd34c ( rs1_data, rs2_data, cin, adder_out );
  input  [33:0] rs1_data;
  input  [33:0] rs2_data;
  input         cin;
  output [33:0] adder_out;
  assign adder_out = rs1_data + rs2_data + cin;
endmodule 
module zzadd32 ( rs1_data, rs2_data, cin, adder_out, cout );
  input  [31:0] rs1_data;   
  input  [31:0] rs2_data;   
  input         cin;        
  output [31:0] adder_out;  
  output 	cout;       
  assign {cout, adder_out} = rs1_data + rs2_data + cin;
endmodule 
module zzadd18 ( rs1_data, rs2_data, cin, adder_out, cout );
  input  [17:0] rs1_data;   
  input  [17:0] rs2_data;   
  input         cin;        
  output [17:0] adder_out;  
  output 	cout;       
  assign {cout, adder_out} = rs1_data + rs2_data + cin;
endmodule 
module zzadd8 ( rs1_data, rs2_data, cin, adder_out, cout );
  input  [7:0] rs1_data;   
  input  [7:0] rs2_data;   
  input        cin;        
  output [7:0] adder_out;  
  output       cout;       
  assign {cout, adder_out} = rs1_data + rs2_data + cin;
endmodule 
module zzadd32op4 ( rs1_data, rs2_data, rs3_data, rs4_data, adder_out );
  input  [31:0] rs1_data;   
  input  [31:0] rs2_data;   
  input  [31:0] rs3_data;   
  input  [31:0] rs4_data;   
  output [31:0] adder_out;  
  assign adder_out = rs1_data + rs2_data + rs3_data + rs4_data;
endmodule 
module zzadd64 ( rs1_data, rs2_data, cin, adder_out, cout32, cout64 );
   input [63:0]  rs1_data;   
   input [63:0]  rs2_data;   
   input         cin;        
   output [63:0] adder_out;  
   output        cout32;     
   output        cout64;     
   assign {cout32, adder_out[31:0]}  = rs1_data[31:0]  + rs2_data[31:0]  + cin;
   assign {cout64, adder_out[63:32]} = rs1_data[63:32] + rs2_data[63:32] + cout32;
endmodule 
module zzadd32v (
   
   z,
   
   a, b, cin, add32
   ) ;
   input [31:0] a;
   input [31:0] b;
   input        cin;
   input        add32;
   output [31:0] z;
   wire          cout15; 
   wire          cin16; 
   wire          cout31; 
   assign        cin16 = (add32)? cout15: cin;
   assign      {cout15, z[15:0]} = a[15:0]+b[15:0]+ cin;
   assign      {cout31, z[31:16]} = a[31:16]+b[31:16]+ cin16;
endmodule 
module zzinc64 ( in, out );
  input  [63:0] in;
  output [63:0] out;   
  assign out = in + 1'b1;
endmodule 
module zzinc48 ( in, out, overflow );
  input  [47:0] in;
  output [47:0] out;      
  output        overflow; 
  assign out      = in + 1'b1;
  assign overflow = ~in[47] & out[47];
endmodule 
module zzinc32 ( in, out );
  input  [31:0] in;
  output [31:0] out;   
  assign out = in + 1'b1;
endmodule 
module zzecc_exu_chkecc2 ( q,ce, ue, ne, d, p, vld );
   input [63:0] d;
   input [7:0]  p;
   input        vld;
   output [6:0] q;
   output       ce,
                ue,
                ne;
   wire       parity;
   assign     ce = vld & parity;
   assign ue = vld & ~parity & (q[6] | q[5] | q[4] | q[3] | q[2] | q[1] | q[0]);
   assign ne = ~vld | ~(parity | q[6] | q[5] | q[4] | q[3] | q[2] | q[1] | q[0]);
   assign q[0] = d[0]  ^ d[1]  ^ d[3]  ^ d[4]  ^ d[6]  ^ d[8]  ^ d[10]
               ^ d[11] ^ d[13] ^ d[15] ^ d[17] ^ d[19] ^ d[21] ^ d[23]
               ^ d[25] ^ d[26] ^ d[28] ^ d[30] ^ d[32] ^ d[34] ^ d[36]
               ^ d[38] ^ d[40] ^ d[42] ^ d[44] ^ d[46] ^ d[48] ^ d[50]
               ^ d[52] ^ d[54] ^ d[56] ^ d[57] ^ d[59] ^ d[61] ^ d[63]
               ^ p[0]  ;
   assign q[1] = d[0]  ^ d[2]  ^ d[3]  ^ d[5]  ^ d[6]  ^ d[9]  ^ d[10]
               ^ d[12] ^ d[13] ^ d[16] ^ d[17] ^ d[20] ^ d[21] ^ d[24]
               ^ d[25] ^ d[27] ^ d[28] ^ d[31] ^ d[32] ^ d[35] ^ d[36]
               ^ d[39] ^ d[40] ^ d[43] ^ d[44] ^ d[47] ^ d[48] ^ d[51]
               ^ d[52] ^ d[55] ^ d[56] ^ d[58] ^ d[59] ^ d[62] ^ d[63]
               ^ p[1]  ;
   assign q[2] = d[1]  ^ d[2]  ^ d[3]  ^ d[7]  ^ d[8]  ^ d[9]  ^ d[10]
               ^ d[14] ^ d[15] ^ d[16] ^ d[17] ^ d[22] ^ d[23] ^ d[24]
               ^ d[25] ^ d[29] ^ d[30] ^ d[31] ^ d[32] ^ d[37] ^ d[38]
               ^ d[39] ^ d[40] ^ d[45] ^ d[46] ^ d[47] ^ d[48] ^ d[53]
               ^ d[54] ^ d[55] ^ d[56] ^ d[60] ^ d[61] ^ d[62] ^ d[63]
               ^ p[2]  ;
   assign q[3] = d[4]  ^ d[5]  ^ d[6]  ^ d[7]  ^ d[8]  ^ d[9]  ^ d[10]
               ^ d[18] ^ d[19] ^ d[20] ^ d[21] ^ d[22] ^ d[23] ^ d[24]
               ^ d[25] ^ d[33] ^ d[34] ^ d[35] ^ d[36] ^ d[37] ^ d[38]
               ^ d[39] ^ d[40] ^ d[49] ^ d[50] ^ d[51] ^ d[52] ^ d[53]
               ^ d[54] ^ d[55] ^ d[56] ^ p[3]  ;
   assign q[4] = d[11] ^ d[12] ^ d[13] ^ d[14] ^ d[15] ^ d[16] ^ d[17]
               ^ d[18] ^ d[19] ^ d[20] ^ d[21] ^ d[22] ^ d[23] ^ d[24]
               ^ d[25] ^ d[41] ^ d[42] ^ d[43] ^ d[44] ^ d[45] ^ d[46]
               ^ d[47] ^ d[48] ^ d[49] ^ d[50] ^ d[51] ^ d[52] ^ d[53]
               ^ d[54] ^ d[55] ^ d[56] ^ p[4]  ;
   assign q[5] = d[26] ^ d[27] ^ d[28] ^ d[29] ^ d[30] ^ d[31] ^ d[32]
               ^ d[33] ^ d[34] ^ d[35] ^ d[36] ^ d[37] ^ d[38] ^ d[39]
               ^ d[40] ^ d[41] ^ d[42] ^ d[43] ^ d[44] ^ d[45] ^ d[46]
               ^ d[47] ^ d[48] ^ d[49] ^ d[50] ^ d[51] ^ d[52] ^ d[53]
               ^ d[54] ^ d[55] ^ d[56] ^ p[5]  ;
   assign q[6] = d[57] ^ d[58] ^ d[59] ^ d[60] ^ d[61] ^ d[62] ^ d[63] ^ p[6] ;
   assign parity = d[0]  ^ d[1]  ^ d[2]  ^ d[3]  ^ d[4]  ^ d[5]  ^ d[6]  ^ d[7]
                 ^ d[8]  ^ d[9]  ^ d[10] ^ d[11] ^ d[12] ^ d[13] ^ d[14] ^ d[15]
                 ^ d[16] ^ d[17] ^ d[18] ^ d[19] ^ d[20] ^ d[21] ^ d[22] ^ d[23]
                 ^ d[24] ^ d[25] ^ d[26] ^ d[27] ^ d[28] ^ d[29] ^ d[30] ^ d[31]
                 ^ d[32] ^ d[33] ^ d[34] ^ d[35] ^ d[36] ^ d[37] ^ d[38] ^ d[39]
                 ^ d[40] ^ d[41] ^ d[42] ^ d[43] ^ d[44] ^ d[45] ^ d[46] ^ d[47]
                 ^ d[48] ^ d[49] ^ d[50] ^ d[51] ^ d[52] ^ d[53] ^ d[54] ^ d[55]
                 ^ d[56] ^ d[57] ^ d[58] ^ d[59] ^ d[60] ^ d[61] ^ d[62] ^ d[63]
                 ^ p[0]  ^ p[1]  ^ p[2]  ^ p[3]  ^ p[4]  ^ p[5]  ^ p[6]  ^ p[7];
endmodule 
module zzecc_sctag_24b_gen ( din, dout, parity ) ;
input  [23:0] din ;
output [23:0] dout ;
output [5:0]  parity ;
wire   [23:0] dout ;
wire   [5:0]  parity ;
wire          p1 ;
wire          p2 ;
wire          p4 ;
wire          p8 ;
wire          p16 ;
wire          p30 ;
assign p1  = din[0]  ^ din[1]  ^ din[3]  ^ din[4]  ^ din[6]  ^ din[8]  ^
             din[10] ^ din[11] ^ din[13] ^ din[15] ^ din[17] ^ din[19] ^
             din[21] ^ din[23] ;
assign p2  = din[0]  ^ din[2]  ^ din[3]  ^ din[5]  ^ din[6]  ^ din[9]  ^
             din[10] ^ din[12] ^ din[13] ^ din[16] ^ din[17] ^ din[20] ^
             din[21] ;
assign p4  = din[1]  ^ din[2]  ^ din[3]  ^ din[7]  ^ din[8]  ^ din[9]  ^
             din[10] ^ din[14] ^ din[15] ^ din[16] ^ din[17] ^ din[22] ^
             din[23] ;
assign p8  = din[4]  ^ din[5]  ^ din[6]  ^ din[7]  ^ din[8]  ^ din[9]  ^
             din[10] ^ din[18] ^ din[19] ^ din[20] ^ din[21] ^ din[22] ^
             din[23] ;
assign p16 = din[11] ^ din[12] ^ din[13] ^ din[14] ^ din[15] ^ din[16] ^
             din[17] ^ din[18] ^ din[19] ^ din[20] ^ din[21] ^ din[22] ^
             din[23] ;
assign p30 = din[0]  ^ din[1]  ^ din[2]  ^ din[4]  ^ din[5]  ^
             din[7]  ^ din[10] ^ din[11] ^ din[12] ^ din[14] ^
             din[17] ^ din[18] ^ din[21] ^ din[23] ;
assign dout   = din ;
assign parity = {p30, p16, p8, p4, p2, p1} ;
endmodule
module zzecc_sctag_30b_cor ( din, parity, dout, corrected_bit ) ;
input  [23:0] din ;
input  [4:0]  parity ;
output [23:0] dout ;
output [4:0]  corrected_bit ;
wire   [23:0] dout ;
wire   [4:0]  corrected_bit ;
wire          p1 ;
wire          p2 ;
wire          p4 ;
wire          p8 ;
wire          p16 ;
wire [23:0]   error_bit ;
assign p1  = parity[0] ^
             din[0]  ^ din[1]  ^ din[3]  ^ din[4]  ^ din[6]  ^ din[8]  ^
             din[10] ^ din[11] ^ din[13] ^ din[15] ^ din[17] ^ din[19] ^
             din[21] ^ din[23] ;
assign p2  = parity[1] ^
             din[0]  ^ din[2]  ^ din[3]  ^ din[5]  ^ din[6]  ^ din[9]  ^
             din[10] ^ din[12] ^ din[13] ^ din[16] ^ din[17] ^ din[20] ^
             din[21] ;
assign p4  = parity[2] ^
             din[1]  ^ din[2]  ^ din[3]  ^ din[7]  ^ din[8]  ^ din[9]  ^
             din[10] ^ din[14] ^ din[15] ^ din[16] ^ din[17] ^ din[22] ^
             din[23] ;
assign p8  = parity[3] ^
             din[4]  ^ din[5]  ^ din[6]  ^ din[7]  ^ din[8]  ^ din[9]  ^
             din[10] ^ din[18] ^ din[19] ^ din[20] ^ din[21] ^ din[22] ^
             din[23] ;
assign p16 = parity[4] ^
             din[11] ^ din[12] ^ din[13] ^ din[14] ^ din[15] ^ din[16] ^
             din[17] ^ din[18] ^ din[19] ^ din[20] ^ din[21] ^ din[22] ^
             din[23] ;
assign  error_bit[0]  = !p16 & !p8 & !p4 &  p2 &  p1 ; 
assign  error_bit[1]  = !p16 & !p8 &  p4 & !p2 &  p1 ; 
assign  error_bit[2]  = !p16 & !p8 &  p4 &  p2 & !p1 ; 
assign  error_bit[3]  = !p16 & !p8 &  p4 &  p2 &  p1 ; 
assign  error_bit[4]  = !p16 &  p8 & !p4 & !p2 &  p1 ; 
assign  error_bit[5]  = !p16 &  p8 & !p4 &  p2 & !p1 ; 
assign  error_bit[6]  = !p16 &  p8 & !p4 &  p2 &  p1 ; 
assign  error_bit[7]  = !p16 &  p8 &  p4 & !p2 & !p1 ; 
assign  error_bit[8]  = !p16 &  p8 &  p4 & !p2 &  p1 ; 
assign  error_bit[9]  = !p16 &  p8 &  p4 &  p2 & !p1 ; 
assign  error_bit[10] = !p16 &  p8 &  p4 &  p2 &  p1 ; 
assign  error_bit[11] =  p16 & !p8 & !p4 & !p2 &  p1 ; 
assign  error_bit[12] =  p16 & !p8 & !p4 &  p2 & !p1 ; 
assign  error_bit[13] =  p16 & !p8 & !p4 &  p2 &  p1 ; 
assign  error_bit[14] =  p16 & !p8 &  p4 & !p2 & !p1 ; 
assign  error_bit[15] =  p16 & !p8 &  p4 & !p2 &  p1 ; 
assign  error_bit[16] =  p16 & !p8 &  p4 &  p2 & !p1 ; 
assign  error_bit[17] =  p16 & !p8 &  p4 &  p2 &  p1 ; 
assign  error_bit[18] =  p16 &  p8 & !p4 & !p2 & !p1 ; 
assign  error_bit[19] =  p16 &  p8 & !p4 & !p2 &  p1 ; 
assign  error_bit[20] =  p16 &  p8 & !p4 &  p2 & !p1 ; 
assign  error_bit[21] =  p16 &  p8 & !p4 &  p2 &  p1 ; 
assign  error_bit[22] =  p16 &  p8 &  p4 & !p2 & !p1 ; 
assign  error_bit[23] =  p16 &  p8 &  p4 & !p2 &  p1 ; 
assign  dout          = din ^ error_bit ;
assign  corrected_bit = {p16, p8, p4, p2, p1} ;
endmodule
module zzecc_sctag_ecc39 ( dout, cflag, pflag, parity, din);
   
   output[31:0] dout;
   output [5:0] cflag;
   output 	pflag;
   
   
   input [31:0] din;
   input [6:0]	parity;
   wire 	c0,c1,c2,c3,c4,c5;
   wire [31:0] 	err_bit_pos;
   
   
   assign c0= parity[0]^(din[0]^din[1])^(din[3]^din[4])^(din[6]^din[8])
                     ^(din[10]^din[11])^(din[13]^din[15])^(din[17]^din[19])
		     ^(din[21]^din[23])^(din[25]^din[26])^(din[28]^din[30]);
   
   assign c1= parity[1]^(din[0]^din[2])^(din[3]^din[5])^(din[6]^din[9])
                     ^(din[10]^din[12])^(din[13]^din[16])^(din[17]^din[20])
		     ^(din[21]^din[24])^(din[25]^din[27])^(din[28]^din[31]);
   
   assign c2= parity[2]^(din[1]^din[2])^(din[3]^din[7])^(din[8]^din[9])
                     ^(din[10]^din[14])^(din[15]^din[16])^(din[17]^din[22])
		     ^(din[23]^din[24])^(din[25]^din[29])^(din[30]^din[31]);
   
   assign c3= parity[3]^(din[4]^din[5])^(din[6]^din[7])^(din[8]^din[9])
                     ^(din[10]^din[18])^(din[19]^din[20])^(din[21]^din[22])
		     ^(din[23]^din[24])^din[25];
   
   assign c4= parity[4]^(din[11]^din[12])^(din[13]^din[14])^
                    (din[15]^din[16])^(din[17]^din[18])^(din[19]^din[20])^
                    (din[21]^din[22])^(din[23]^din[24])^din[25];
   assign c5= parity[5]^(din[26]^din[27])^(din[28]^din[29])^
		    (din[30]^din[31]);
   
   assign pflag= c0 ^
		(( (((parity[1]^parity[2])^(parity[3]^parity[4])) ^
		 ((parity[5]^parity[6])^(din[2]^din[5]))) ^		 
		 (((din[7]^din[9])^(din[12]^din[14])) ^
		 ((din[16]^din[18])^(din[20]^din[22]))) ) ^
		 ((din[24]^din[27])^(din[29]^din[31])) );
   
   assign cflag= {c5,c4,c3,c2,c1,c0};
   
   
   assign err_bit_pos[0] = (c0)&(c1)&(~c2)&(~c3)&(~c4)&(~c5);
   assign err_bit_pos[1] = (c0)&(~c1)&(c2)&(~c3)&(~c4)&(~c5);
   assign err_bit_pos[2] = (~c0)&(c1)&(c2)&(~c3)&(~c4)&(~c5);
   assign err_bit_pos[3] = (c0)&(c1)&(c2)&(~c3)&(~c4)&(~c5);
   assign err_bit_pos[4] = (c0)&(~c1)&(~c2)&(c3)&(~c4)&(~c5);
   assign err_bit_pos[5] = (~c0)&(c1)&(~c2)&(c3)&(~c4)&(~c5);
   assign err_bit_pos[6] = (c0)&(c1)&(~c2)&(c3)&(~c4)&(~c5);
   assign err_bit_pos[7] = (~c0)&(~c1)&(c2)&(c3)&(~c4)&(~c5);
   assign err_bit_pos[8] = (c0)&(~c1)&(c2)&(c3)&(~c4)&(~c5);
   assign err_bit_pos[9] = (~c0)&(c1)&(c2)&(c3)&(~c4)&(~c5);
   assign err_bit_pos[10] = (c0)&(c1)&(c2)&(c3)&(~c4)&(~c5);
   assign err_bit_pos[11] = (c0)&(~c1)&(~c2)&(~c3)&(c4)&(~c5);
   assign err_bit_pos[12] = (~c0)&(c1)&(~c2)&(~c3)&(c4)&(~c5);
   assign err_bit_pos[13] = (c0)&(c1)&(~c2)&(~c3)&(c4)&(~c5);
   assign err_bit_pos[14] = (~c0)&(~c1)&(c2)&(~c3)&(c4)&(~c5);
   assign err_bit_pos[15] = (c0)&(~c1)&(c2)&(~c3)&(c4)&(~c5);
   assign err_bit_pos[16] = (~c0)&(c1)&(c2)&(~c3)&(c4)&(~c5);
   assign err_bit_pos[17] = (c0)&(c1)&(c2)&(~c3)&(c4)&(~c5);
   assign err_bit_pos[18] = (~c0)&(~c1)&(~c2)&(c3)&(c4)&(~c5);
   assign err_bit_pos[19] = (c0)&(~c1)&(~c2)&(c3)&(c4)&(~c5);
   assign err_bit_pos[20] = (~c0)&(c1)&(~c2)&(c3)&(c4)&(~c5);
   assign err_bit_pos[21] = (c0)&(c1)&(~c2)&(c3)&(c4)&(~c5);
   assign err_bit_pos[22] = (~c0)&(~c1)&(c2)&(c3)&(c4)&(~c5);
   assign err_bit_pos[23] = (c0)&(~c1)&(c2)&(c3)&(c4)&(~c5);
   assign err_bit_pos[24] = (~c0)&(c1)&(c2)&(c3)&(c4)&(~c5);
   assign err_bit_pos[25] = (c0)&(c1)&(c2)&(c3)&(c4)&(~c5);
   assign err_bit_pos[26] = (c0)&(~c1)&(~c2)&(~c3)&(~c4)&(c5);
   assign err_bit_pos[27] = (~c0)&(c1)&(~c2)&(~c3)&(~c4)&(c5);
   assign err_bit_pos[28] = (c0)&(c1)&(~c2)&(~c3)&(~c4)&(c5);
   assign err_bit_pos[29] = (~c0)&(~c1)&(c2)&(~c3)&(~c4)&(c5);
   assign err_bit_pos[30] = (c0)&(~c1)&(c2)&(~c3)&(~c4)&(c5);
   assign err_bit_pos[31] = (~c0)&(c1)&(c2)&(~c3)&(~c4)&(c5);
   
   
   assign dout = din ^ err_bit_pos;
endmodule 
module zzecc_sctag_pgen_32b ( dout, parity, din);
   
   output[31:0] dout;
   output [6:0] parity;
   
   input [31:0] din;
   
   assign dout = din ;
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   assign parity[0] = (din[0]^din[1])^(din[3]^din[4])^(din[6]^din[8])
                     ^(din[10]^din[11])^(din[13]^din[15])^(din[17]^din[19])
		     ^(din[21]^din[23])^(din[25]^din[26])^(din[28]^din[30]);
   
   assign parity[1] = (din[0]^din[2])^(din[3]^din[5])^(din[6]^din[9])
                     ^(din[10]^din[12])^(din[13]^din[16])^(din[17]^din[20])
		     ^(din[21]^din[24])^(din[25]^din[27])^(din[28]^din[31]);
   
   assign parity[2] = (din[1]^din[2])^(din[3]^din[7])^(din[8]^din[9])
                     ^(din[10]^din[14])^(din[15]^din[16])^(din[17]^din[22])
		     ^(din[23]^din[24])^(din[25]^din[29])^(din[30]^din[31]);
   
   assign parity[3] = (din[4]^din[5])^(din[6]^din[7])^(din[8]^din[9])
                     ^(din[10]^din[18])^(din[19]^din[20])^(din[21]^din[22])
		     ^(din[23]^din[24])^din[25];
   
   assign parity[4] = (din[11]^din[12])^(din[13]^din[14])^(din[15]^din[16])
                     ^(din[17]^din[18])^(din[19]^din[20])^(din[21]^din[22])
		     ^(din[23]^din[24])^din[25];
   
   assign parity[5] = (din[26]^din[27])^(din[28]^din[29])^(din[30]^din[31]);
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   assign parity[6] =  din[0] ^ din[1]  ^ din[2]  ^ din[4]  ^ din[5] ^ din[7]
		    ^ din[10] ^ din[11] ^ din[12] ^ din[14] ^ din[17]
		    ^ din[18] ^ din[21] ^ din[23] ^ din[24] ^ din[26]
		    ^ din[27] ^ din[29];
   
endmodule 
module zzpar34 ( z, d );
   input  [33:0] d;
   output        z;
   assign  z =  d[0]  ^ d[1]  ^ d[2]  ^ d[3]  ^ d[4]  ^ d[5]  ^ d[6]  ^ d[7]
	      ^ d[8]  ^ d[9]  ^ d[10] ^ d[11] ^ d[12] ^ d[13] ^ d[14] ^ d[15]
	      ^ d[16] ^ d[17] ^ d[18] ^ d[19] ^ d[20] ^ d[21] ^ d[22] ^ d[23]
	      ^ d[24] ^ d[25] ^ d[26] ^ d[27] ^ d[28] ^ d[29] ^ d[30] ^ d[31]
	      ^ d[32] ^ d[33]; 
endmodule 
module zzpar32 ( z, d );
   input  [31:0] d;
   output        z;
   assign  z =  d[0]  ^ d[1]  ^ d[2]  ^ d[3]  ^ d[4]  ^ d[5]  ^ d[6]  ^ d[7]
	      ^ d[8]  ^ d[9]  ^ d[10] ^ d[11] ^ d[12] ^ d[13] ^ d[14] ^ d[15]
	      ^ d[16] ^ d[17] ^ d[18] ^ d[19] ^ d[20] ^ d[21] ^ d[22] ^ d[23]
	      ^ d[24] ^ d[25] ^ d[26] ^ d[27] ^ d[28] ^ d[29] ^ d[30] ^ d[31]; 
endmodule 
module zzpar28 ( z, d );
   input  [27:0] d;
   output        z;
   assign  z =  d[0]  ^ d[1]  ^ d[2]  ^ d[3]  ^ d[4]  ^ d[5]  ^ d[6]  ^ d[7]
	      ^ d[8]  ^ d[9]  ^ d[10] ^ d[11] ^ d[12] ^ d[13] ^ d[14] ^ d[15]
	      ^ d[16] ^ d[17] ^ d[18] ^ d[19] ^ d[20] ^ d[21] ^ d[22] ^ d[23]
	      ^ d[24] ^ d[25] ^ d[26] ^ d[27]; 
endmodule 
module zzpar16 ( z, d );
   input  [15:0] d;
   output        z;
   assign z = d[0] ^ d[1] ^ d[2]  ^ d[3]  ^ d[4]  ^ d[5]  ^ d[6]  ^ d[7]
	    ^ d[8] ^ d[9] ^ d[10] ^ d[11] ^ d[12] ^ d[13] ^ d[14] ^ d[15]; 
   
endmodule 
module zzpar8 ( z, d );
   input  [7:0] d;
   output       z;
   assign  z =  d[0] ^ d[1] ^ d[2] ^ d[3] ^ d[4] ^ d[5] ^ d[6] ^ d[7]; 
endmodule 
module zzpenc64 (
   
   z, 
   
  a 
   );
   input [63:0] a;
   output [5:0] z;
   integer      i;
   reg  [5:0]   z;
     always @ (a)
     begin
          z = 6'b0;
          for (i=0;i<64;i=i+1)
               if (a[i])
                      z = i;
     end
endmodule 
module zzbufh_60x4 (
   
   z,
   
  a
   );
   input [3:0] a;
   output [3:0] z;
   assign z = a;
endmodule 
module zzadd64_lv ( rs1_data, rs2_data, cin, adder_out, cout32, cout64 );
   input [63:0]  rs1_data;   
   input [63:0]  rs2_data;   
   input         cin;        
   output [63:0] adder_out;  
   output        cout32;     
   output        cout64;     
   assign {cout32, adder_out[31:0]}  = rs1_data[31:0]  + rs2_data[31:0]  + cin;
   assign {cout64, adder_out[63:32]} = rs1_data[63:32] + rs2_data[63:32] + cout32;
endmodule 
module zzpar8_lv ( z, d );
   input  [7:0] d;
   output       z;
   assign  z =  d[0] ^ d[1] ^ d[2] ^ d[3] ^ d[4] ^ d[5] ^ d[6] ^ d[7]; 
endmodule 
module zzpar32_lv ( z, d );
   input  [31:0] d;
   output        z;
   assign  z =  d[0]  ^ d[1]  ^ d[2]  ^ d[3]  ^ d[4]  ^ d[5]  ^ d[6]  ^ d[7]
              ^ d[8]  ^ d[9]  ^ d[10] ^ d[11] ^ d[12] ^ d[13] ^ d[14] ^ d[15]
              ^ d[16] ^ d[17] ^ d[18] ^ d[19] ^ d[20] ^ d[21] ^ d[22] ^ d[23]
              ^ d[24] ^ d[25] ^ d[26] ^ d[27] ^ d[28] ^ d[29] ^ d[30] ^ d[31];
endmodule 
module zznor64_32_lv ( znor64, znor32, a );
  input  [63:0] a;
  output        znor64;
  output        znor32;
  assign znor32 =  ~(a[0]  | a[1]  | a[2]  | a[3]  | a[4]  | a[5]  | a[6]  | a[7]
		   | a[8]  | a[9]  | a[10] | a[11] | a[12] | a[13] | a[14] | a[15]
		   | a[16] | a[17] | a[18] | a[19] | a[20] | a[21] | a[22] | a[23]
		   | a[24] | a[25] | a[26] | a[27] | a[28] | a[29] | a[30] | a[31]); 
  assign znor64 =  ~(a[0]  | a[1]  | a[2]  | a[3]  | a[4]  | a[5]  | a[6]  | a[7]
		   | a[8]  | a[9]  | a[10] | a[11] | a[12] | a[13] | a[14] | a[15]
		   | a[16] | a[17] | a[18] | a[19] | a[20] | a[21] | a[22] | a[23]
		   | a[24] | a[25] | a[26] | a[27] | a[28] | a[29] | a[30] | a[31] 
		   | a[32] | a[33] | a[34] | a[35] | a[36] | a[37] | a[38] | a[39] 
		   | a[40] | a[41] | a[42] | a[43] | a[44] | a[45] | a[46] | a[47] 
		   | a[48] | a[49] | a[50] | a[51] | a[52] | a[53] | a[54] | a[55] 
		   | a[56] | a[57] | a[58] | a[59] | a[60] | a[61] | a[62] | a[63]);
endmodule 
module zzpenc64_lv (
   
   z,
   
  a
   );
   input [63:0] a;
   output [5:0] z;
   integer      i;
   reg  [5:0]   z;
     always @ (a)
     begin
          z = 6'b0;
          for (i=0;i<64;i=i+1)
               if (a[i])
                      z = i;
     end
endmodule 
module zzor36_lv ( z, a );
  input  [35:0] a;
  output        z;
  assign z =  (a[0]  | a[1]  | a[2]  | a[3]  | a[4]  | a[5]  | a[6]  | a[7]
             | a[8]  | a[9]  | a[10] | a[11] | a[12] | a[13] | a[14] | a[15]
             | a[16] | a[17] | a[18] | a[19] | a[20] | a[21] | a[22] | a[23]
             | a[24] | a[25] | a[26] | a[27] | a[28] | a[29] | a[30] | a[31]
             | a[32] | a[33] | a[34] | a[35]);
endmodule 
module zzpar34_lv ( z, d );
   input  [33:0] d;
   output        z;
   assign  z =  d[0]  ^ d[1]  ^ d[2]  ^ d[3]  ^ d[4]  ^ d[5]  ^ d[6]  ^ d[7]
              ^ d[8]  ^ d[9]  ^ d[10] ^ d[11] ^ d[12] ^ d[13] ^ d[14] ^ d[15]
              ^ d[16] ^ d[17] ^ d[18] ^ d[19] ^ d[20] ^ d[21] ^ d[22] ^ d[23]
              ^ d[24] ^ d[25] ^ d[26] ^ d[27] ^ d[28] ^ d[29] ^ d[30] ^ d[31]
              ^ d[32] ^ d[33];
endmodule 
module mul64 (rs1_l, rs2, valid, areg, accreg, x2, out, rclk, si, so, se, mul_rst_l, mul_step);
input  [63:0]  	rs1_l;			
input  [63:0]  	rs2;			
input	       	valid;			
input  [96:0]  	areg;			
input  [135:129] accreg;		
input	       	x2;			
input	       	rclk, si, se, mul_rst_l, mul_step;
output  	so;
output [135:0] 	out;
wire	       	cyc1, cyc2, cyc3;	
wire [2:0]	b0, b1, b2,  b3,  b4,  b5,  b6,  b7;
wire [2:0]	b8, b9, b10, b11, b12, b13, b14, b15;
wire	    	b16;
wire [63:0]	op1_l, op1;
wire [81:0]	a0sum, a1sum, a0s, a1s; 
wire [81:4]	a0cout, a1cout, a0c, a1c;
wire		pcoutx2, psumx2;
wire 		x2_c1, x2_c2, x2_c3, x2_c2c3;
wire [98:0]	psum, pcout;
wire [98:30]	pcout_in, pc;
wire [98:31]	psum_in, ps;
wire [96:0]	ary2_cout, addin_cout;
wire [97:0]	ary2_sum,  addin_sum ;
wire		add_cin, addin_cin, add_co31, add_co96;
wire [103:0]	addout;
wire		clk_enb0, clk_enb1;
wire 		rst;
wire		clk;
wire		tm_l;
  assign clk = rclk;
  assign rst = ~mul_rst_l; 
  assign tm_l = ~se;
  clken_buf	ckbuf_0(.clk(clk_enb0), .rclk(clk), .enb_l(~mul_step), .tmb_l(tm_l));
  
  
  
  dffr_s  cyc1_dff(.din(valid), .clk(clk_enb0), .q(cyc1), .rst(rst), .se(se), .si(), .so());
  dffr_s  cyc2_dff(.din(cyc1),  .clk(clk_enb0), .q(cyc2), .rst(rst), .se(se), .si(), .so());
  dffr_s  cyc3_dff(.din(cyc2),  .clk(clk_enb0), .q(cyc3), .rst(rst), .se(se), .si(), .so());
  dffr_s  x2c1_dff(.din(x2),    .clk(clk_enb0), .q(x2_c1), .rst(rst), .se(se), .si(), .so());
  dffr_s  x2c2_dff(.din(x2_c1), .clk(clk_enb0), .q(x2_c2), .rst(rst), .se(se), .si(), .so());
  dffr_s  x2c3_dff(.din(x2_c2), .clk(clk_enb0), .q(x2_c3), .rst(rst), .se(se), .si(), .so());
  assign x2_c2c3 =  x2_c2 | x2_c3 ;
	
  
  
  
  clken_buf	ckbuf_1(.clk(clk_enb1), .rclk(clk), .enb_l(~(valid & mul_step)), .tmb_l(tm_l));
  dff_s #(64)  	ffrs1  (.din(rs1_l[63:0]), .clk(clk_enb1), .q(op1_l[63:0]),
			.se(se), .si(), .so());
  assign op1[63:0] = ~op1_l[63:0];
  mul_booth	 booth (.head (valid),
			.b_in (rs2),
			.b0   (b0),
			.b1   (b1),
			.b2   (b2),
			.b3   (b3),
			.b4   (b4),
			.b5   (b5),
			.b6   (b6),
			.b7   (b7),
			.b8   (b8),
			.b9   (b9),
			.b10  (b10),
			.b11  (b11),
			.b12  (b12),
			.b13  (b13),
			.b14  (b14),
			.b15  (b15),
			.b16  (b16),
			.clk  (clk), .se(se), .si(), .so(), .mul_step(mul_step), .tm_l(tm_l));
			
  
  
  
  mul_array1	ary1_a0(.cout (a0cout[81:4]),
			.sum  (a0sum[81:0]),
			.a    (op1),
			.b0   (b0),
			.b1   (b1),
			.b2   (b2),
			.b3   (b3),
			.b4   (b4),
			.b5   (b5),
			.b6   (b6),
			.b7   (b7),
			.b8   (3'b000),
			.head (cyc1),
			.bot  (1'b0)); 
 
  dff_s #(78)  a0cot_dff (.din(a0cout[81:4]), .clk(clk_enb0), .q(a0c[81:4]),
			.se(se), .si(), .so());
  dff_s #(82)  a0sum_dff (.din(a0sum[81:0]), .clk(clk_enb0), .q(a0s[81:0]),
			.se(se), .si(), .so());
  mul_array1	ary1_a1(.cout (a1cout[81:4]),
			.sum  (a1sum[81:0]),
			.a    (op1),
			.b0   (b8),
			.b1   (b9),
			.b2   (b10),
			.b3   (b11),
			.b4   (b12),
			.b5   (b13),
			.b6   (b14),
			.b7   (b15),
			.b8   ({1'b0,b16,1'b0}),
			.head (1'b0),	
			.bot  (cyc2)); 
  dff_s #(78)  a1cot_dff (.din(a1cout[81:4]), .clk(clk_enb0), .q(a1c[81:4]),
			.se(se), .si(), .so());
  dff_s #(82)  a1sum_dff (.din(a1sum[81:0]), .clk(clk_enb0), .q(a1s[81:0]),
			.se(se), .si(), .so());
  
  
  
  mul_array2 	 array2(.pcoutx2 (pcoutx2),
			.psumx2  (psumx2),
			.pcout 	 (pcout[98:0]),
			.psum    (psum[98:0]), 
			.a0c     (a0c[81:4]),
			.a0s     (a0s[81:0]),
			.a1c     (a1c[81:4]),
			.a1s     (a1s[81:0]),
			.pc	 (pc[98:30]),
			.ps	 (ps[98:31]),
			.areg    (areg[96:0]),
			.bot     (cyc3),
			.x2      (x2_c2c3));
 
  
  dp_mux2es #(97)  ary2_cmux (.dout(ary2_cout[96:0]),
                              .in0(pcout[96:0]),
                              .in1({pcout[95:0],pcoutx2}),
                              .sel(x2_c2c3));
  dff_s #(97)  a2cot_dff (.din(ary2_cout[96:0]), .clk(clk_enb0), .q(addin_cout[96:0]), 
              		.se(se), .si(), .so());
  dp_mux2es #(98) ary2_smux (.dout(ary2_sum[97:0]),
                             .in0(psum[97:0]),
                             .in1({psum[96:0],psumx2}),
                             .sel(x2_c2c3));
  dff_s #(98)  a2sum_dff (.din(ary2_sum[97:0]), .clk(clk_enb0), .q(addin_sum[97:0]), 
			.se(se), .si(), .so());
  
  assign psum_in[98:32]  = psum[98:32] & {67{cyc2}} ;
  assign psum_in[31]     = psum[31] & x2_c2 ;
  assign pcout_in[98:31] = pcout[98:31] & {68{cyc2}} ;
  assign pcout_in[30]    = pcout[30] & x2_c2 ;
  
  dff_s #(68)  psum_dff  (.din(psum_in[98:31]), .clk(clk_enb0), .q(ps[98:31]),
                	.se(se), .si(), .so());
  dff_s #(69)  pcout_dff (.din(pcout_in[98:30]), .clk(clk_enb0), .q(pc[98:30]),
            		.se(se), .si(), .so());
  
  
  
  assign 	add_cin = add_co31 & cyc3 ;
  assign {add_co31,addout[31:0]} =   {{1'b0},addin_sum[31:0]} 
		     		   + {{1'b0},addin_cout[30:0],addin_cin} ;
  assign {add_co96,addout[96:32]} =  addin_sum[97:32]	
				  + addin_cout[96:31]
				  + {{65'b0},add_co31} ;
  assign 	addout[103:97] =  accreg[135:129] + {{6'b0},add_co96} ;
  
  
  
  dff_s  	      co31_dff (.din(add_cin), .clk(clk_enb0), .q(addin_cin),
       			.se(se), .si(), .so());
  dff_s #(104)   out_dff (.din(addout[103:0]), .clk(clk_enb0), .q(out[135:32]),
              		.se(se), .si(), .so());
  dff_s #(32)    pip_dff (.din(out[63:32]), .clk(clk_enb0), .q(out[31:0]),
               		.se(se), .si(), .so());
endmodule 
module mul_array1 ( cout, sum, a, b0, b1, b2, b3, b4, b5, b6, b7, b8,
     bot, head );
input  bot, head;
output [81:4]  cout;
output [81:0]  sum;
input [2:0]  b6;
input [2:0]  b3;
input [2:0]  b8;
input [2:0]  b2;
input [2:0]  b1;
input [2:0]  b7;
input [63:0]  a;
input [2:0]  b0;
input [2:0]  b4;
input [2:0]  b5;
wire  [1:0]  b5n;
wire  [1:0]  b2n;
wire  [68:1]  c0;
wire  [69:0]  s1;
wire  [68:1]  c1;
wire  [69:0]  s2;
wire  [68:1]  c2;
wire  [70:4]  s_1;
wire  [69:2]  s0;
wire  [76:10]  s_2;
wire  [70:2]  c_1;
wire  [76:10]  c_2;
wire  [75:11]  co;
mul_negen p1n ( .b(b5[2:0]), .n1(b5n[1]), .n0(b5n[0]));
mul_negen p0n ( .b(b2[2:0]), .n1(b2n[1]), .n0(b2n[0]));
mul_csa42  sc3_71_ ( .c(s_2[71]), .cin(co[70]), .a(c_1[70]),
     .b(c_2[70]), .cout(co[71]), .sum(sum[71]), .d(s1[65]),
     .carry(cout[71]));
mul_csa42  sc3_75_ ( .c(s_2[75]), .cin(co[74]), .a(1'b0),
     .b(c_2[74]), .cout(co[75]), .sum(sum[75]), .d(s1[69]),
     .carry(cout[75]));
mul_csa42  sc3_74_ ( .c(s_2[74]), .cin(co[73]), .a(1'b0),
     .b(c_2[73]), .cout(co[74]), .sum(sum[74]), .d(s1[68]),
     .carry(cout[74]));
mul_csa42  sc3_73_ ( .c(s_2[73]), .cin(co[72]), .a(1'b0),
     .b(c_2[72]), .cout(co[73]), .sum(sum[73]), .d(s1[67]),
     .carry(cout[73]));
mul_csa42  sc3_72_ ( .c(s_2[72]), .cin(co[71]), .a(1'b0),
     .b(c_2[71]), .cout(co[72]), .sum(sum[72]), .d(s1[66]),
     .carry(cout[72]));
mul_csa42  sc3_76_ ( .c(s_2[76]), .cin(co[75]), .a(1'b0),
     .b(c_2[75]), .cout(), .sum(sum[76]), .d(1'b0),
     .carry(cout[76]));
mul_csa42  sc3_70_ ( .c(s_2[70]), .cin(co[69]), .a(c_1[69]),
     .b(c_2[69]), .cout(co[70]), .sum(sum[70]), .d(s_1[70]),
     .carry(cout[70]));
mul_csa42  sc3_69_ ( .c(s_2[69]), .cin(co[68]), .a(c_1[68]),
     .b(c_2[68]), .cout(co[69]), .sum(sum[69]), .d(s_1[69]),
     .carry(cout[69]));
mul_csa42  sc3_68_ ( .c(s_2[68]), .cin(co[67]), .a(c_1[67]),
     .b(c_2[67]), .cout(co[68]), .sum(sum[68]), .d(s_1[68]),
     .carry(cout[68]));
mul_csa42  sc3_67_ ( .c(s_2[67]), .cin(co[66]), .a(c_1[66]),
     .b(c_2[66]), .cout(co[67]), .sum(sum[67]), .d(s_1[67]),
     .carry(cout[67]));
mul_csa42  sc3_66_ ( .c(s_2[66]), .cin(co[65]), .a(c_1[65]),
     .b(c_2[65]), .cout(co[66]), .sum(sum[66]), .d(s_1[66]),
     .carry(cout[66]));
mul_csa42  sc3_65_ ( .c(s_2[65]), .cin(co[64]), .a(c_1[64]),
     .b(c_2[64]), .cout(co[65]), .sum(sum[65]), .d(s_1[65]),
     .carry(cout[65]));
mul_csa42  sc3_64_ ( .c(s_2[64]), .cin(co[63]), .a(c_1[63]),
     .b(c_2[63]), .cout(co[64]), .sum(sum[64]), .d(s_1[64]),
     .carry(cout[64]));
mul_csa42  sc3_63_ ( .c(s_2[63]), .cin(co[62]), .a(c_1[62]),
     .b(c_2[62]), .cout(co[63]), .sum(sum[63]), .d(s_1[63]),
     .carry(cout[63]));
mul_csa42  sc3_62_ ( .c(s_2[62]), .cin(co[61]), .a(c_1[61]),
     .b(c_2[61]), .cout(co[62]), .sum(sum[62]), .d(s_1[62]),
     .carry(cout[62]));
mul_csa42  sc3_61_ ( .c(s_2[61]), .cin(co[60]), .a(c_1[60]),
     .b(c_2[60]), .cout(co[61]), .sum(sum[61]), .d(s_1[61]),
     .carry(cout[61]));
mul_csa42  sc3_60_ ( .c(s_2[60]), .cin(co[59]), .a(c_1[59]),
     .b(c_2[59]), .cout(co[60]), .sum(sum[60]), .d(s_1[60]),
     .carry(cout[60]));
mul_csa42  sc3_59_ ( .c(s_2[59]), .cin(co[58]), .a(c_1[58]),
     .b(c_2[58]), .cout(co[59]), .sum(sum[59]), .d(s_1[59]),
     .carry(cout[59]));
mul_csa42  sc3_58_ ( .c(s_2[58]), .cin(co[57]), .a(c_1[57]),
     .b(c_2[57]), .cout(co[58]), .sum(sum[58]), .d(s_1[58]),
     .carry(cout[58]));
mul_csa42  sc3_57_ ( .c(s_2[57]), .cin(co[56]), .a(c_1[56]),
     .b(c_2[56]), .cout(co[57]), .sum(sum[57]), .d(s_1[57]),
     .carry(cout[57]));
mul_csa42  sc3_56_ ( .c(s_2[56]), .cin(co[55]), .a(c_1[55]),
     .b(c_2[55]), .cout(co[56]), .sum(sum[56]), .d(s_1[56]),
     .carry(cout[56]));
mul_csa42  sc3_55_ ( .c(s_2[55]), .cin(co[54]), .a(c_1[54]),
     .b(c_2[54]), .cout(co[55]), .sum(sum[55]), .d(s_1[55]),
     .carry(cout[55]));
mul_csa42  sc3_54_ ( .c(s_2[54]), .cin(co[53]), .a(c_1[53]),
     .b(c_2[53]), .cout(co[54]), .sum(sum[54]), .d(s_1[54]),
     .carry(cout[54]));
mul_csa42  sc3_53_ ( .c(s_2[53]), .cin(co[52]), .a(c_1[52]),
     .b(c_2[52]), .cout(co[53]), .sum(sum[53]), .d(s_1[53]),
     .carry(cout[53]));
mul_csa42  sc3_52_ ( .c(s_2[52]), .cin(co[51]), .a(c_1[51]),
     .b(c_2[51]), .cout(co[52]), .sum(sum[52]), .d(s_1[52]),
     .carry(cout[52]));
mul_csa42  sc3_51_ ( .c(s_2[51]), .cin(co[50]), .a(c_1[50]),
     .b(c_2[50]), .cout(co[51]), .sum(sum[51]), .d(s_1[51]),
     .carry(cout[51]));
mul_csa42  sc3_50_ ( .c(s_2[50]), .cin(co[49]), .a(c_1[49]),
     .b(c_2[49]), .cout(co[50]), .sum(sum[50]), .d(s_1[50]),
     .carry(cout[50]));
mul_csa42  sc3_49_ ( .c(s_2[49]), .cin(co[48]), .a(c_1[48]),
     .b(c_2[48]), .cout(co[49]), .sum(sum[49]), .d(s_1[49]),
     .carry(cout[49]));
mul_csa42  sc3_48_ ( .c(s_2[48]), .cin(co[47]), .a(c_1[47]),
     .b(c_2[47]), .cout(co[48]), .sum(sum[48]), .d(s_1[48]),
     .carry(cout[48]));
mul_csa42  sc3_47_ ( .c(s_2[47]), .cin(co[46]), .a(c_1[46]),
     .b(c_2[46]), .cout(co[47]), .sum(sum[47]), .d(s_1[47]),
     .carry(cout[47]));
mul_csa42  sc3_46_ ( .c(s_2[46]), .cin(co[45]), .a(c_1[45]),
     .b(c_2[45]), .cout(co[46]), .sum(sum[46]), .d(s_1[46]),
     .carry(cout[46]));
mul_csa42  sc3_45_ ( .c(s_2[45]), .cin(co[44]), .a(c_1[44]),
     .b(c_2[44]), .cout(co[45]), .sum(sum[45]), .d(s_1[45]),
     .carry(cout[45]));
mul_csa42  sc3_44_ ( .c(s_2[44]), .cin(co[43]), .a(c_1[43]),
     .b(c_2[43]), .cout(co[44]), .sum(sum[44]), .d(s_1[44]),
     .carry(cout[44]));
mul_csa42  sc3_43_ ( .c(s_2[43]), .cin(co[42]), .a(c_1[42]),
     .b(c_2[42]), .cout(co[43]), .sum(sum[43]), .d(s_1[43]),
     .carry(cout[43]));
mul_csa42  sc3_42_ ( .c(s_2[42]), .cin(co[41]), .a(c_1[41]),
     .b(c_2[41]), .cout(co[42]), .sum(sum[42]), .d(s_1[42]),
     .carry(cout[42]));
mul_csa42  sc3_41_ ( .c(s_2[41]), .cin(co[40]), .a(c_1[40]),
     .b(c_2[40]), .cout(co[41]), .sum(sum[41]), .d(s_1[41]),
     .carry(cout[41]));
mul_csa42  sc3_40_ ( .c(s_2[40]), .cin(co[39]), .a(c_1[39]),
     .b(c_2[39]), .cout(co[40]), .sum(sum[40]), .d(s_1[40]),
     .carry(cout[40]));
mul_csa42  sc3_39_ ( .c(s_2[39]), .cin(co[38]), .a(c_1[38]),
     .b(c_2[38]), .cout(co[39]), .sum(sum[39]), .d(s_1[39]),
     .carry(cout[39]));
mul_csa42  sc3_38_ ( .c(s_2[38]), .cin(co[37]), .a(c_1[37]),
     .b(c_2[37]), .cout(co[38]), .sum(sum[38]), .d(s_1[38]),
     .carry(cout[38]));
mul_csa42  sc3_37_ ( .c(s_2[37]), .cin(co[36]), .a(c_1[36]),
     .b(c_2[36]), .cout(co[37]), .sum(sum[37]), .d(s_1[37]),
     .carry(cout[37]));
mul_csa42  sc3_36_ ( .c(s_2[36]), .cin(co[35]), .a(c_1[35]),
     .b(c_2[35]), .cout(co[36]), .sum(sum[36]), .d(s_1[36]),
     .carry(cout[36]));
mul_csa42  sc3_35_ ( .c(s_2[35]), .cin(co[34]), .a(c_1[34]),
     .b(c_2[34]), .cout(co[35]), .sum(sum[35]), .d(s_1[35]),
     .carry(cout[35]));
mul_csa42  sc3_34_ ( .c(s_2[34]), .cin(co[33]), .a(c_1[33]),
     .b(c_2[33]), .cout(co[34]), .sum(sum[34]), .d(s_1[34]),
     .carry(cout[34]));
mul_csa42  sc3_33_ ( .c(s_2[33]), .cin(co[32]), .a(c_1[32]),
     .b(c_2[32]), .cout(co[33]), .sum(sum[33]), .d(s_1[33]),
     .carry(cout[33]));
mul_csa42  sc3_32_ ( .c(s_2[32]), .cin(co[31]), .a(c_1[31]),
     .b(c_2[31]), .cout(co[32]), .sum(sum[32]), .d(s_1[32]),
     .carry(cout[32]));
mul_csa42  sc3_31_ ( .c(s_2[31]), .cin(co[30]), .a(c_1[30]),
     .b(c_2[30]), .cout(co[31]), .sum(sum[31]), .d(s_1[31]),
     .carry(cout[31]));
mul_csa42  sc3_30_ ( .c(s_2[30]), .cin(co[29]), .a(c_1[29]),
     .b(c_2[29]), .cout(co[30]), .sum(sum[30]), .d(s_1[30]),
     .carry(cout[30]));
mul_csa42  sc3_29_ ( .c(s_2[29]), .cin(co[28]), .a(c_1[28]),
     .b(c_2[28]), .cout(co[29]), .sum(sum[29]), .d(s_1[29]),
     .carry(cout[29]));
mul_csa42  sc3_28_ ( .c(s_2[28]), .cin(co[27]), .a(c_1[27]),
     .b(c_2[27]), .cout(co[28]), .sum(sum[28]), .d(s_1[28]),
     .carry(cout[28]));
mul_csa42  sc3_27_ ( .c(s_2[27]), .cin(co[26]), .a(c_1[26]),
     .b(c_2[26]), .cout(co[27]), .sum(sum[27]), .d(s_1[27]),
     .carry(cout[27]));
mul_csa42  sc3_26_ ( .c(s_2[26]), .cin(co[25]), .a(c_1[25]),
     .b(c_2[25]), .cout(co[26]), .sum(sum[26]), .d(s_1[26]),
     .carry(cout[26]));
mul_csa42  sc3_25_ ( .c(s_2[25]), .cin(co[24]), .a(c_1[24]),
     .b(c_2[24]), .cout(co[25]), .sum(sum[25]), .d(s_1[25]),
     .carry(cout[25]));
mul_csa42  sc3_24_ ( .c(s_2[24]), .cin(co[23]), .a(c_1[23]),
     .b(c_2[23]), .cout(co[24]), .sum(sum[24]), .d(s_1[24]),
     .carry(cout[24]));
mul_csa42  sc3_23_ ( .c(s_2[23]), .cin(co[22]), .a(c_1[22]),
     .b(c_2[22]), .cout(co[23]), .sum(sum[23]), .d(s_1[23]),
     .carry(cout[23]));
mul_csa42  sc3_22_ ( .c(s_2[22]), .cin(co[21]), .a(c_1[21]),
     .b(c_2[21]), .cout(co[22]), .sum(sum[22]), .d(s_1[22]),
     .carry(cout[22]));
mul_csa42  sc3_21_ ( .c(s_2[21]), .cin(co[20]), .a(c_1[20]),
     .b(c_2[20]), .cout(co[21]), .sum(sum[21]), .d(s_1[21]),
     .carry(cout[21]));
mul_csa42  sc3_20_ ( .c(s_2[20]), .cin(co[19]), .a(c_1[19]),
     .b(c_2[19]), .cout(co[20]), .sum(sum[20]), .d(s_1[20]),
     .carry(cout[20]));
mul_csa42  sc3_19_ ( .c(s_2[19]), .cin(co[18]), .a(c_1[18]),
     .b(c_2[18]), .cout(co[19]), .sum(sum[19]), .d(s_1[19]),
     .carry(cout[19]));
mul_csa42  sc3_18_ ( .c(s_2[18]), .cin(co[17]), .a(c_1[17]),
     .b(c_2[17]), .cout(co[18]), .sum(sum[18]), .d(s_1[18]),
     .carry(cout[18]));
mul_csa42  sc3_17_ ( .c(s_2[17]), .cin(co[16]), .a(c_1[16]),
     .b(c_2[16]), .cout(co[17]), .sum(sum[17]), .d(s_1[17]),
     .carry(cout[17]));
mul_csa42  sc3_16_ ( .c(s_2[16]), .cin(co[15]), .a(c_1[15]),
     .b(c_2[15]), .cout(co[16]), .sum(sum[16]), .d(s_1[16]),
     .carry(cout[16]));
mul_csa42  sc3_15_ ( .c(s_2[15]), .cin(co[14]), .a(c_1[14]),
     .b(c_2[14]), .cout(co[15]), .sum(sum[15]), .d(s_1[15]),
     .carry(cout[15]));
mul_csa42  sc3_14_ ( .c(s_2[14]), .cin(co[13]), .a(c_1[13]),
     .b(c_2[13]), .cout(co[14]), .sum(sum[14]), .d(s_1[14]),
     .carry(cout[14]));
mul_csa42  sc3_13_ ( .c(s_2[13]), .cin(co[12]), .a(c_1[12]),
     .b(c_2[12]), .cout(co[13]), .sum(sum[13]), .d(s_1[13]),
     .carry(cout[13]));
mul_csa42  sc3_12_ ( .c(s_2[12]), .cin(co[11]), .a(c_1[11]),
     .b(c_2[11]), .cout(co[12]), .sum(sum[12]), .d(s_1[12]),
     .carry(cout[12]));
mul_csa42  sc3_11_ ( .c(s_2[11]), .cin(1'b0),
     .a(c_1[10]), .b(c_2[10]), .cout(co[11]), .sum(sum[11]),
     .d(s_1[11]), .carry(cout[11]));
mul_csa32  sc2_2_70_ ( .c(c1[63]), .b(c2[57]), .a(s2[58]),
     .cout(c_2[70]), .sum(s_2[70]));
mul_csa32  sc2_2_69_ ( .c(c1[62]), .b(c2[56]), .a(s2[57]),
     .cout(c_2[69]), .sum(s_2[69]));
mul_csa32  sc2_2_68_ ( .c(c1[61]), .b(c2[55]), .a(s2[56]),
     .cout(c_2[68]), .sum(s_2[68]));
mul_csa32  sc2_2_67_ ( .c(c1[60]), .b(c2[54]), .a(s2[55]),
     .cout(c_2[67]), .sum(s_2[67]));
mul_csa32  sc2_2_66_ ( .c(c1[59]), .b(c2[53]), .a(s2[54]),
     .cout(c_2[66]), .sum(s_2[66]));
mul_csa32  sc2_2_65_ ( .c(c1[58]), .b(c2[52]), .a(s2[53]),
     .cout(c_2[65]), .sum(s_2[65]));
mul_csa32  sc2_2_64_ ( .c(c1[57]), .b(c2[51]), .a(s2[52]),
     .cout(c_2[64]), .sum(s_2[64]));
mul_csa32  sc2_2_63_ ( .c(c1[56]), .b(c2[50]), .a(s2[51]),
     .cout(c_2[63]), .sum(s_2[63]));
mul_csa32  sc2_2_62_ ( .c(c1[55]), .b(c2[49]), .a(s2[50]),
     .cout(c_2[62]), .sum(s_2[62]));
mul_csa32  sc2_2_61_ ( .c(c1[54]), .b(c2[48]), .a(s2[49]),
     .cout(c_2[61]), .sum(s_2[61]));
mul_csa32  sc2_2_60_ ( .c(c1[53]), .b(c2[47]), .a(s2[48]),
     .cout(c_2[60]), .sum(s_2[60]));
mul_csa32  sc2_2_59_ ( .c(c1[52]), .b(c2[46]), .a(s2[47]),
     .cout(c_2[59]), .sum(s_2[59]));
mul_csa32  sc2_2_58_ ( .c(c1[51]), .b(c2[45]), .a(s2[46]),
     .cout(c_2[58]), .sum(s_2[58]));
mul_csa32  sc2_2_57_ ( .c(c1[50]), .b(c2[44]), .a(s2[45]),
     .cout(c_2[57]), .sum(s_2[57]));
mul_csa32  sc2_2_56_ ( .c(c1[49]), .b(c2[43]), .a(s2[44]),
     .cout(c_2[56]), .sum(s_2[56]));
mul_csa32  sc2_2_55_ ( .c(c1[48]), .b(c2[42]), .a(s2[43]),
     .cout(c_2[55]), .sum(s_2[55]));
mul_csa32  sc2_2_54_ ( .c(c1[47]), .b(c2[41]), .a(s2[42]),
     .cout(c_2[54]), .sum(s_2[54]));
mul_csa32  sc2_2_53_ ( .c(c1[46]), .b(c2[40]), .a(s2[41]),
     .cout(c_2[53]), .sum(s_2[53]));
mul_csa32  sc2_2_52_ ( .c(c1[45]), .b(c2[39]), .a(s2[40]),
     .cout(c_2[52]), .sum(s_2[52]));
mul_csa32  sc2_2_51_ ( .c(c1[44]), .b(c2[38]), .a(s2[39]),
     .cout(c_2[51]), .sum(s_2[51]));
mul_csa32  sc2_2_50_ ( .c(c1[43]), .b(c2[37]), .a(s2[38]),
     .cout(c_2[50]), .sum(s_2[50]));
mul_csa32  sc2_2_49_ ( .c(c1[42]), .b(c2[36]), .a(s2[37]),
     .cout(c_2[49]), .sum(s_2[49]));
mul_csa32  sc2_2_48_ ( .c(c1[41]), .b(c2[35]), .a(s2[36]),
     .cout(c_2[48]), .sum(s_2[48]));
mul_csa32  sc2_2_47_ ( .c(c1[40]), .b(c2[34]), .a(s2[35]),
     .cout(c_2[47]), .sum(s_2[47]));
mul_csa32  sc2_2_46_ ( .c(c1[39]), .b(c2[33]), .a(s2[34]),
     .cout(c_2[46]), .sum(s_2[46]));
mul_csa32  sc2_2_45_ ( .c(c1[38]), .b(c2[32]), .a(s2[33]),
     .cout(c_2[45]), .sum(s_2[45]));
mul_csa32  sc2_2_44_ ( .c(c1[37]), .b(c2[31]), .a(s2[32]),
     .cout(c_2[44]), .sum(s_2[44]));
mul_csa32  sc2_2_43_ ( .c(c1[36]), .b(c2[30]), .a(s2[31]),
     .cout(c_2[43]), .sum(s_2[43]));
mul_csa32  sc2_2_42_ ( .c(c1[35]), .b(c2[29]), .a(s2[30]),
     .cout(c_2[42]), .sum(s_2[42]));
mul_csa32  sc2_2_41_ ( .c(c1[34]), .b(c2[28]), .a(s2[29]),
     .cout(c_2[41]), .sum(s_2[41]));
mul_csa32  sc2_2_40_ ( .c(c1[33]), .b(c2[27]), .a(s2[28]),
     .cout(c_2[40]), .sum(s_2[40]));
mul_csa32  sc2_2_39_ ( .c(c1[32]), .b(c2[26]), .a(s2[27]),
     .cout(c_2[39]), .sum(s_2[39]));
mul_csa32  sc2_2_38_ ( .c(c1[31]), .b(c2[25]), .a(s2[26]),
     .cout(c_2[38]), .sum(s_2[38]));
mul_csa32  sc2_2_37_ ( .c(c1[30]), .b(c2[24]), .a(s2[25]),
     .cout(c_2[37]), .sum(s_2[37]));
mul_csa32  sc2_2_36_ ( .c(c1[29]), .b(c2[23]), .a(s2[24]),
     .cout(c_2[36]), .sum(s_2[36]));
mul_csa32  sc2_2_35_ ( .c(c1[28]), .b(c2[22]), .a(s2[23]),
     .cout(c_2[35]), .sum(s_2[35]));
mul_csa32  sc2_2_34_ ( .c(c1[27]), .b(c2[21]), .a(s2[22]),
     .cout(c_2[34]), .sum(s_2[34]));
mul_csa32  sc2_2_33_ ( .c(c1[26]), .b(c2[20]), .a(s2[21]),
     .cout(c_2[33]), .sum(s_2[33]));
mul_csa32  sc2_2_32_ ( .c(c1[25]), .b(c2[19]), .a(s2[20]),
     .cout(c_2[32]), .sum(s_2[32]));
mul_csa32  sc2_2_31_ ( .c(c1[24]), .b(c2[18]), .a(s2[19]),
     .cout(c_2[31]), .sum(s_2[31]));
mul_csa32  sc2_2_30_ ( .c(c1[23]), .b(c2[17]), .a(s2[18]),
     .cout(c_2[30]), .sum(s_2[30]));
mul_csa32  sc2_2_29_ ( .c(c1[22]), .b(c2[16]), .a(s2[17]),
     .cout(c_2[29]), .sum(s_2[29]));
mul_csa32  sc2_2_28_ ( .c(c1[21]), .b(c2[15]), .a(s2[16]),
     .cout(c_2[28]), .sum(s_2[28]));
mul_csa32  sc2_2_27_ ( .c(c1[20]), .b(c2[14]), .a(s2[15]),
     .cout(c_2[27]), .sum(s_2[27]));
mul_csa32  sc2_2_26_ ( .c(c1[19]), .b(c2[13]), .a(s2[14]),
     .cout(c_2[26]), .sum(s_2[26]));
mul_csa32  sc2_2_25_ ( .c(c1[18]), .b(c2[12]), .a(s2[13]),
     .cout(c_2[25]), .sum(s_2[25]));
mul_csa32  sc2_2_24_ ( .c(c1[17]), .b(c2[11]), .a(s2[12]),
     .cout(c_2[24]), .sum(s_2[24]));
mul_csa32  sc2_2_23_ ( .c(c1[16]), .b(c2[10]), .a(s2[11]),
     .cout(c_2[23]), .sum(s_2[23]));
mul_csa32  sc2_2_22_ ( .c(c1[15]), .b(c2[9]), .a(s2[10]),
     .cout(c_2[22]), .sum(s_2[22]));
mul_csa32  sc2_2_21_ ( .c(c1[14]), .b(c2[8]), .a(s2[9]),
     .cout(c_2[21]), .sum(s_2[21]));
mul_csa32  sc2_2_20_ ( .c(c1[13]), .b(c2[7]), .a(s2[8]),
     .cout(c_2[20]), .sum(s_2[20]));
mul_csa32  sc2_2_19_ ( .c(c1[12]), .b(c2[6]), .a(s2[7]),
     .cout(c_2[19]), .sum(s_2[19]));
mul_csa32  sc2_2_18_ ( .c(c1[11]), .b(c2[5]), .a(s2[6]),
     .cout(c_2[18]), .sum(s_2[18]));
mul_csa32  sc2_2_17_ ( .c(c1[10]), .b(c2[4]), .a(s2[5]),
     .cout(c_2[17]), .sum(s_2[17]));
mul_csa32  sc2_2_16_ ( .c(c1[9]), .b(c2[3]), .a(s2[4]),
     .cout(c_2[16]), .sum(s_2[16]));
mul_csa32  sc2_2_15_ ( .c(c1[8]), .b(c2[2]), .a(s2[3]),
     .cout(c_2[15]), .sum(s_2[15]));
mul_csa32  sc2_2_14_ ( .c(c1[7]), .b(c2[1]), .a(s2[2]),
     .cout(c_2[14]), .sum(s_2[14]));
mul_csa32  sc2_2_13_ ( .c(c1[6]), .b(s1[7]), .a(s2[1]),
     .cout(c_2[13]), .sum(s_2[13]));
mul_csa32  sc2_2_12_ ( .c(c1[5]), .b(s1[6]), .a(s2[0]),
     .cout(c_2[12]), .sum(s_2[12]));
mul_csa32  sc2_2_11_ ( .c(c1[4]), .b(s1[5]), .a(b5n[1]),
     .cout(c_2[11]), .sum(s_2[11]));
mul_csa32  sc2_2_10_ ( .c(c1[3]), .b(s1[4]), .a(b5n[0]),
     .cout(c_2[10]), .sum(s_2[10]));
mul_csa32  sc2_2_76_ ( .c(1'b1), .b(c2[63]), .a(s2[64]),
     .cout(c_2[76]), .sum(s_2[76]));
mul_csa32  sc2_2_77_ ( .c(c_2[76]), .b(c2[64]), .a(s2[65]),
     .cout(cout[77]), .sum(sum[77]));
mul_csa32  sc2_1_9_ ( .c(s1[3]), .b(c0[8]), .a(s0[9]), .cout(c_1[9]),
     .sum(s_1[9]));
mul_csa32  sc2_1_8_ ( .c(s1[2]), .b(c0[7]), .a(s0[8]), .cout(c_1[8]),
     .sum(s_1[8]));
mul_csa32  sc2_1_3_ ( .c(c_1[2]), .b(c0[2]), .a(s0[3]),
     .cout(c_1[3]), .sum(sum[3]));
mul_csa32  sc3_10_ ( .c(s_2[10]), .b(s_1[10]), .a(c_1[9]),
     .cout(cout[10]), .sum(sum[10]));
mul_csa32  sc3_9_ ( .c(c1[2]), .sum(sum[9]), .cout(cout[9]),
     .a(c_1[8]), .b(s_1[9]));
mul_csa32  sc3_8_ ( .c(c1[1]), .sum(sum[8]), .cout(cout[8]),
     .a(c_1[7]), .b(s_1[8]));
mul_csa32  sc2_2_71_ ( .c(c1[64]), .b(c2[58]), .a(s2[59]),
     .cout(c_2[71]), .sum(s_2[71]));
mul_csa32  sc2_2_75_ ( .c(c1[68]), .b(c2[62]), .a(s2[63]),
     .cout(c_2[75]), .sum(s_2[75]));
mul_csa32  sc2_2_74_ ( .c(c1[67]), .b(c2[61]), .a(s2[62]),
     .cout(c_2[74]), .sum(s_2[74]));
mul_csa32  sc2_2_73_ ( .c(c1[66]), .b(c2[60]), .a(s2[61]),
     .cout(c_2[73]), .sum(s_2[73]));
mul_csa32  sc2_2_72_ ( .c(c1[65]), .b(c2[59]), .a(s2[60]),
     .cout(c_2[72]), .sum(s_2[72]));
mul_csa32  sc2_1_69_ ( .c(s1[63]), .sum(s_1[69]), .cout(c_1[69]),
     .a(s0[69]), .b(c0[68]));
mul_csa32  sc2_1_68_ ( .c(s1[62]), .sum(s_1[68]), .cout(c_1[68]),
     .a(s0[68]), .b(c0[67]));
mul_csa32  sc2_1_67_ ( .c(s1[61]), .sum(s_1[67]), .cout(c_1[67]),
     .a(s0[67]), .b(c0[66]));
mul_csa32  sc2_1_66_ ( .c(s1[60]), .sum(s_1[66]), .cout(c_1[66]),
     .a(s0[66]), .b(c0[65]));
mul_csa32  sc2_1_65_ ( .c(s1[59]), .sum(s_1[65]), .cout(c_1[65]),
     .a(s0[65]), .b(c0[64]));
mul_csa32  sc2_1_64_ ( .c(s1[58]), .sum(s_1[64]), .cout(c_1[64]),
     .a(s0[64]), .b(c0[63]));
mul_csa32  sc2_1_63_ ( .c(s1[57]), .sum(s_1[63]), .cout(c_1[63]),
     .a(s0[63]), .b(c0[62]));
mul_csa32  sc2_1_62_ ( .c(s1[56]), .sum(s_1[62]), .cout(c_1[62]),
     .a(s0[62]), .b(c0[61]));
mul_csa32  sc2_1_61_ ( .c(s1[55]), .sum(s_1[61]), .cout(c_1[61]),
     .a(s0[61]), .b(c0[60]));
mul_csa32  sc2_1_60_ ( .c(s1[54]), .sum(s_1[60]), .cout(c_1[60]),
     .a(s0[60]), .b(c0[59]));
mul_csa32  sc2_1_59_ ( .c(s1[53]), .sum(s_1[59]), .cout(c_1[59]),
     .a(s0[59]), .b(c0[58]));
mul_csa32  sc2_1_58_ ( .c(s1[52]), .sum(s_1[58]), .cout(c_1[58]),
     .a(s0[58]), .b(c0[57]));
mul_csa32  sc2_1_57_ ( .c(s1[51]), .sum(s_1[57]), .cout(c_1[57]),
     .a(s0[57]), .b(c0[56]));
mul_csa32  sc2_1_56_ ( .c(s1[50]), .sum(s_1[56]), .cout(c_1[56]),
     .a(s0[56]), .b(c0[55]));
mul_csa32  sc2_1_55_ ( .c(s1[49]), .sum(s_1[55]), .cout(c_1[55]),
     .a(s0[55]), .b(c0[54]));
mul_csa32  sc2_1_54_ ( .c(s1[48]), .sum(s_1[54]), .cout(c_1[54]),
     .a(s0[54]), .b(c0[53]));
mul_csa32  sc2_1_53_ ( .c(s1[47]), .sum(s_1[53]), .cout(c_1[53]),
     .a(s0[53]), .b(c0[52]));
mul_csa32  sc2_1_52_ ( .c(s1[46]), .sum(s_1[52]), .cout(c_1[52]),
     .a(s0[52]), .b(c0[51]));
mul_csa32  sc2_1_51_ ( .c(s1[45]), .sum(s_1[51]), .cout(c_1[51]),
     .a(s0[51]), .b(c0[50]));
mul_csa32  sc2_1_50_ ( .c(s1[44]), .sum(s_1[50]), .cout(c_1[50]),
     .a(s0[50]), .b(c0[49]));
mul_csa32  sc2_1_49_ ( .c(s1[43]), .sum(s_1[49]), .cout(c_1[49]),
     .a(s0[49]), .b(c0[48]));
mul_csa32  sc2_1_48_ ( .c(s1[42]), .sum(s_1[48]), .cout(c_1[48]),
     .a(s0[48]), .b(c0[47]));
mul_csa32  sc2_1_47_ ( .c(s1[41]), .sum(s_1[47]), .cout(c_1[47]),
     .a(s0[47]), .b(c0[46]));
mul_csa32  sc2_1_46_ ( .c(s1[40]), .sum(s_1[46]), .cout(c_1[46]),
     .a(s0[46]), .b(c0[45]));
mul_csa32  sc2_1_45_ ( .c(s1[39]), .sum(s_1[45]), .cout(c_1[45]),
     .a(s0[45]), .b(c0[44]));
mul_csa32  sc2_1_44_ ( .c(s1[38]), .sum(s_1[44]), .cout(c_1[44]),
     .a(s0[44]), .b(c0[43]));
mul_csa32  sc2_1_43_ ( .c(s1[37]), .sum(s_1[43]), .cout(c_1[43]),
     .a(s0[43]), .b(c0[42]));
mul_csa32  sc2_1_42_ ( .c(s1[36]), .sum(s_1[42]), .cout(c_1[42]),
     .a(s0[42]), .b(c0[41]));
mul_csa32  sc2_1_41_ ( .c(s1[35]), .sum(s_1[41]), .cout(c_1[41]),
     .a(s0[41]), .b(c0[40]));
mul_csa32  sc2_1_40_ ( .c(s1[34]), .sum(s_1[40]), .cout(c_1[40]),
     .a(s0[40]), .b(c0[39]));
mul_csa32  sc2_1_39_ ( .c(s1[33]), .sum(s_1[39]), .cout(c_1[39]),
     .a(s0[39]), .b(c0[38]));
mul_csa32  sc2_1_38_ ( .c(s1[32]), .sum(s_1[38]), .cout(c_1[38]),
     .a(s0[38]), .b(c0[37]));
mul_csa32  sc2_1_37_ ( .c(s1[31]), .sum(s_1[37]), .cout(c_1[37]),
     .a(s0[37]), .b(c0[36]));
mul_csa32  sc2_1_36_ ( .c(s1[30]), .sum(s_1[36]), .cout(c_1[36]),
     .a(s0[36]), .b(c0[35]));
mul_csa32  sc2_1_35_ ( .c(s1[29]), .sum(s_1[35]), .cout(c_1[35]),
     .a(s0[35]), .b(c0[34]));
mul_csa32  sc2_1_34_ ( .c(s1[28]), .sum(s_1[34]), .cout(c_1[34]),
     .a(s0[34]), .b(c0[33]));
mul_csa32  sc2_1_33_ ( .c(s1[27]), .sum(s_1[33]), .cout(c_1[33]),
     .a(s0[33]), .b(c0[32]));
mul_csa32  sc2_1_32_ ( .c(s1[26]), .sum(s_1[32]), .cout(c_1[32]),
     .a(s0[32]), .b(c0[31]));
mul_csa32  sc2_1_31_ ( .c(s1[25]), .sum(s_1[31]), .cout(c_1[31]),
     .a(s0[31]), .b(c0[30]));
mul_csa32  sc2_1_30_ ( .c(s1[24]), .sum(s_1[30]), .cout(c_1[30]),
     .a(s0[30]), .b(c0[29]));
mul_csa32  sc2_1_29_ ( .c(s1[23]), .sum(s_1[29]), .cout(c_1[29]),
     .a(s0[29]), .b(c0[28]));
mul_csa32  sc2_1_28_ ( .c(s1[22]), .sum(s_1[28]), .cout(c_1[28]),
     .a(s0[28]), .b(c0[27]));
mul_csa32  sc2_1_27_ ( .c(s1[21]), .sum(s_1[27]), .cout(c_1[27]),
     .a(s0[27]), .b(c0[26]));
mul_csa32  sc2_1_26_ ( .c(s1[20]), .sum(s_1[26]), .cout(c_1[26]),
     .a(s0[26]), .b(c0[25]));
mul_csa32  sc2_1_25_ ( .c(s1[19]), .sum(s_1[25]), .cout(c_1[25]),
     .a(s0[25]), .b(c0[24]));
mul_csa32  sc2_1_24_ ( .c(s1[18]), .sum(s_1[24]), .cout(c_1[24]),
     .a(s0[24]), .b(c0[23]));
mul_csa32  sc2_1_23_ ( .c(s1[17]), .sum(s_1[23]), .cout(c_1[23]),
     .a(s0[23]), .b(c0[22]));
mul_csa32  sc2_1_22_ ( .c(s1[16]), .sum(s_1[22]), .cout(c_1[22]),
     .a(s0[22]), .b(c0[21]));
mul_csa32  sc2_1_21_ ( .c(s1[15]), .sum(s_1[21]), .cout(c_1[21]),
     .a(s0[21]), .b(c0[20]));
mul_csa32  sc2_1_20_ ( .c(s1[14]), .sum(s_1[20]), .cout(c_1[20]),
     .a(s0[20]), .b(c0[19]));
mul_csa32  sc2_1_19_ ( .c(s1[13]), .sum(s_1[19]), .cout(c_1[19]),
     .a(s0[19]), .b(c0[18]));
mul_csa32  sc2_1_18_ ( .c(s1[12]), .sum(s_1[18]), .cout(c_1[18]),
     .a(s0[18]), .b(c0[17]));
mul_csa32  sc2_1_17_ ( .c(s1[11]), .sum(s_1[17]), .cout(c_1[17]),
     .a(s0[17]), .b(c0[16]));
mul_csa32  sc2_1_16_ ( .c(s1[10]), .sum(s_1[16]), .cout(c_1[16]),
     .a(s0[16]), .b(c0[15]));
mul_csa32  sc2_1_15_ ( .c(s1[9]), .sum(s_1[15]), .cout(c_1[15]),
     .a(s0[15]), .b(c0[14]));
mul_csa32  sc2_1_14_ ( .c(s1[8]), .sum(s_1[14]), .cout(c_1[14]),
     .a(s0[14]), .b(c0[13]));
mul_csa32  sc2_1_7_ ( .c(s1[1]), .b(c0[6]), .a(s0[7]), .cout(c_1[7]),
     .sum(s_1[7]));
mul_csa32  sc2_1_6_ ( .c(s1[0]), .b(c0[5]), .a(s0[6]), .cout(c_1[6]),
     .sum(s_1[6]));
mul_csa32  sc2_1_5_ ( .c(b2n[1]), .b(c0[4]), .a(s0[5]),
     .cout(c_1[5]), .sum(s_1[5]));
mul_csa32  sc2_1_4_ ( .c(b2n[0]), .b(c0[3]), .a(s0[4]),
     .cout(c_1[4]), .sum(s_1[4]));
mul_ha sc2_1_10_ ( .sum(s_1[10]), .cout(c_1[10]), .a(s0[10]),
     .b(c0[9]));
mul_ha sc3_7_ ( .sum(sum[7]), .cout(cout[7]), .a(c_1[6]),
     .b(s_1[7]));
mul_ha sc3_6_ ( .sum(sum[6]), .cout(cout[6]), .a(c_1[5]),
     .b(s_1[6]));
mul_ha sc3_5_ ( .sum(sum[5]), .cout(cout[5]), .a(c_1[4]),
     .b(s_1[5]));
mul_ha sc3_4_ ( .sum(sum[4]), .cout(cout[4]), .a(c_1[3]),
     .b(s_1[4]));
mul_ha sc2_2_81_ ( .sum(sum[81]), .cout(cout[81]), .a(s2[69]),
     .b(c2[68]));
mul_ha sc2_2_80_ ( .sum(sum[80]), .cout(cout[80]), .a(s2[68]),
     .b(c2[67]));
mul_ha sc2_2_79_ ( .sum(sum[79]), .cout(cout[79]), .a(s2[67]),
     .b(c2[66]));
mul_ha sc2_2_78_ ( .sum(sum[78]), .cout(cout[78]), .a(s2[66]),
     .b(c2[65]));
mul_ha sc2_1_70_ ( .sum(s_1[70]), .cout(c_1[70]),
     .a(1'b1), .b(s1[64]));
mul_ha sc2_1_2_ ( .sum(sum[2]), .cout(c_1[2]), .a(s0[2]), .b(c0[1]));
mul_ha sc2_1_13_ ( .sum(s_1[13]), .cout(c_1[13]), .a(s0[13]),
     .b(c0[12]));
mul_ha sc2_1_12_ ( .sum(s_1[12]), .cout(c_1[12]), .a(s0[12]),
     .b(c0[11]));
mul_ha sc2_1_11_ ( .sum(s_1[11]), .cout(c_1[11]), .a(s0[11]),
     .b(c0[10]));
mul_ppgenrow3 I2 ( .head(1'b0), .bot(bot), .b2(b8[2:0]),
     .b1(b7[2:0]), .b0(b6[2:0]), .a(a[63:0]), .sum(s2[69:0]),
     .cout(c2[68:1]));
mul_ppgenrow3 I1 ( .head(1'b0), .bot(1'b1),
     .b2(b5[2:0]), .b1(b4[2:0]), .b0(b3[2:0]), .a(a[63:0]),
     .sum(s1[69:0]), .cout(c1[68:1]));
mul_ppgenrow3 I0 ( .head(head), .bot(1'b1), .b2(b2[2:0]),
     .b1(b1[2:0]), .b0(b0[2:0]), .a(a[63:0]), .sum({s0[69:2],
     sum[1:0]}), .cout(c0[68:1]));
endmodule 
module mul_array2 ( pcout, pcoutx2, psum, psumx2, a0c, a0s, a1c, a1s,
     areg, bot, pc, ps, x2 );
output  pcoutx2, psumx2;
input  bot, x2;
output [98:0]  psum;
output [98:0]  pcout;
input [81:4]  a1c;
input [98:30]  pc;
input [98:31]  ps;
input [81:0]  a0s;
input [96:0]  areg;
input [81:0]  a1s;
input [81:4]  a0c;
wire  [81:15]  s3;
wire  [81:15]  c3;
wire  [96:0]  ain;
wire  [67:20]  co;
wire  [82:0]  s1;
wire  [96:0]  c2;
wire  [82:0]  c1;
wire  [96:0]  s2;
wire	      ainx2, s1x2, c1x2;
mul_mux2 sh_82_ ( .d1(areg[83]), .z(ain[82]), .d0(areg[82]), .s(x2));
mul_mux2 sh_68_ ( .d1(areg[69]), .z(ain[68]), .d0(areg[68]), .s(x2));
mul_mux2 sh_67_ ( .d1(areg[68]), .z(ain[67]), .d0(areg[67]), .s(x2));
mul_mux2 sh_66_ ( .d1(areg[67]), .z(ain[66]), .d0(areg[66]), .s(x2));
mul_mux2 sh_65_ ( .d1(areg[66]), .z(ain[65]), .d0(areg[65]), .s(x2));
mul_mux2 sh_64_ ( .d1(areg[65]), .z(ain[64]), .d0(areg[64]), .s(x2));
mul_mux2 sh_63_ ( .d1(areg[64]), .z(ain[63]), .d0(areg[63]), .s(x2));
mul_mux2 sh_62_ ( .d1(areg[63]), .z(ain[62]), .d0(areg[62]), .s(x2));
mul_mux2 sh_61_ ( .d1(areg[62]), .z(ain[61]), .d0(areg[61]), .s(x2));
mul_mux2 sh_60_ ( .d1(areg[61]), .z(ain[60]), .d0(areg[60]), .s(x2));
mul_mux2 sh_59_ ( .d1(areg[60]), .z(ain[59]), .d0(areg[59]), .s(x2));
mul_mux2 sh_58_ ( .d1(areg[59]), .z(ain[58]), .d0(areg[58]), .s(x2));
mul_mux2 sh_57_ ( .d1(areg[58]), .z(ain[57]), .d0(areg[57]), .s(x2));
mul_mux2 sh_56_ ( .d1(areg[57]), .z(ain[56]), .d0(areg[56]), .s(x2));
mul_mux2 sh_55_ ( .d1(areg[56]), .z(ain[55]), .d0(areg[55]), .s(x2));
mul_mux2 sh_54_ ( .d1(areg[55]), .z(ain[54]), .d0(areg[54]), .s(x2));
mul_mux2 sh_53_ ( .d1(areg[54]), .z(ain[53]), .d0(areg[53]), .s(x2));
mul_mux2 sh_52_ ( .d1(areg[53]), .z(ain[52]), .d0(areg[52]), .s(x2));
mul_mux2 sh_51_ ( .d1(areg[52]), .z(ain[51]), .d0(areg[51]), .s(x2));
mul_mux2 sh_50_ ( .d1(areg[51]), .z(ain[50]), .d0(areg[50]), .s(x2));
mul_mux2 sh_49_ ( .d1(areg[50]), .z(ain[49]), .d0(areg[49]), .s(x2));
mul_mux2 sh_48_ ( .d1(areg[49]), .z(ain[48]), .d0(areg[48]), .s(x2));
mul_mux2 sh_47_ ( .d1(areg[48]), .z(ain[47]), .d0(areg[47]), .s(x2));
mul_mux2 sh_46_ ( .d1(areg[47]), .z(ain[46]), .d0(areg[46]), .s(x2));
mul_mux2 sh_45_ ( .d1(areg[46]), .z(ain[45]), .d0(areg[45]), .s(x2));
mul_mux2 sh_44_ ( .d1(areg[45]), .z(ain[44]), .d0(areg[44]), .s(x2));
mul_mux2 sh_43_ ( .d1(areg[44]), .z(ain[43]), .d0(areg[43]), .s(x2));
mul_mux2 sh_42_ ( .d1(areg[43]), .z(ain[42]), .d0(areg[42]), .s(x2));
mul_mux2 sh_41_ ( .d1(areg[42]), .z(ain[41]), .d0(areg[41]), .s(x2));
mul_mux2 sh_40_ ( .d1(areg[41]), .z(ain[40]), .d0(areg[40]), .s(x2));
mul_mux2 sh_39_ ( .d1(areg[40]), .z(ain[39]), .d0(areg[39]), .s(x2));
mul_mux2 sh_38_ ( .d1(areg[39]), .z(ain[38]), .d0(areg[38]), .s(x2));
mul_mux2 sh_37_ ( .d1(areg[38]), .z(ain[37]), .d0(areg[37]), .s(x2));
mul_mux2 sh_36_ ( .d1(areg[37]), .z(ain[36]), .d0(areg[36]), .s(x2));
mul_mux2 sh_35_ ( .d1(areg[36]), .z(ain[35]), .d0(areg[35]), .s(x2));
mul_mux2 sh_34_ ( .d1(areg[35]), .z(ain[34]), .d0(areg[34]), .s(x2));
mul_mux2 sh_33_ ( .d1(areg[34]), .z(ain[33]), .d0(areg[33]), .s(x2));
mul_mux2 sh_32_ ( .d1(areg[33]), .z(ain[32]), .d0(areg[32]), .s(x2));
mul_mux2 sh_31_ ( .d1(areg[32]), .z(ain[31]), .d0(areg[31]), .s(x2));
mul_mux2 sh_30_ ( .d1(areg[31]), .z(ain[30]), .d0(areg[30]), .s(x2));
mul_mux2 sh_29_ ( .d1(areg[30]), .z(ain[29]), .d0(areg[29]), .s(x2));
mul_mux2 sh_28_ ( .d1(areg[29]), .z(ain[28]), .d0(areg[28]), .s(x2));
mul_mux2 sh_27_ ( .d1(areg[28]), .z(ain[27]), .d0(areg[27]), .s(x2));
mul_mux2 sh_26_ ( .d1(areg[27]), .z(ain[26]), .d0(areg[26]), .s(x2));
mul_mux2 sh_25_ ( .d1(areg[26]), .z(ain[25]), .d0(areg[25]), .s(x2));
mul_mux2 sh_24_ ( .d1(areg[25]), .z(ain[24]), .d0(areg[24]), .s(x2));
mul_mux2 sh_23_ ( .d1(areg[24]), .z(ain[23]), .d0(areg[23]), .s(x2));
mul_mux2 sh_22_ ( .d1(areg[23]), .z(ain[22]), .d0(areg[22]), .s(x2));
mul_mux2 sh_21_ ( .d1(areg[22]), .z(ain[21]), .d0(areg[21]), .s(x2));
mul_mux2 sh_20_ ( .d1(areg[21]), .z(ain[20]), .d0(areg[20]), .s(x2));
mul_mux2 sh_96_ ( .d1(1'b0), .z(ain[96]), .d0(areg[96]),
     .s(x2));
mul_mux2 sh_95_ ( .d1(areg[96]), .z(ain[95]), .d0(areg[95]), .s(x2));
mul_mux2 sh_94_ ( .d1(areg[95]), .z(ain[94]), .d0(areg[94]), .s(x2));
mul_mux2 sh_93_ ( .d1(areg[94]), .z(ain[93]), .d0(areg[93]), .s(x2));
mul_mux2 sh_92_ ( .d1(areg[93]), .z(ain[92]), .d0(areg[92]), .s(x2));
mul_mux2 sh_91_ ( .d1(areg[92]), .z(ain[91]), .d0(areg[91]), .s(x2));
mul_mux2 sh_90_ ( .d1(areg[91]), .z(ain[90]), .d0(areg[90]), .s(x2));
mul_mux2 sh_89_ ( .d1(areg[90]), .z(ain[89]), .d0(areg[89]), .s(x2));
mul_mux2 sh_88_ ( .d1(areg[89]), .z(ain[88]), .d0(areg[88]), .s(x2));
mul_mux2 sh_87_ ( .d1(areg[88]), .z(ain[87]), .d0(areg[87]), .s(x2));
mul_mux2 sh_86_ ( .d1(areg[87]), .z(ain[86]), .d0(areg[86]), .s(x2));
mul_mux2 sh_85_ ( .d1(areg[86]), .z(ain[85]), .d0(areg[85]), .s(x2));
mul_mux2 sh_84_ ( .d1(areg[85]), .z(ain[84]), .d0(areg[84]), .s(x2));
mul_mux2 sh_0_ ( .d1(areg[1]), .z(ain[0]), .d0(areg[0]), .s(x2));
mul_mux2 sh_81_ ( .d1(areg[82]), .z(ain[81]), .d0(areg[81]), .s(x2));
mul_mux2 sh_80_ ( .d1(areg[81]), .z(ain[80]), .d0(areg[80]), .s(x2));
mul_mux2 sh_79_ ( .d1(areg[80]), .z(ain[79]), .d0(areg[79]), .s(x2));
mul_mux2 sh_78_ ( .d1(areg[79]), .z(ain[78]), .d0(areg[78]), .s(x2));
mul_mux2 sh_77_ ( .d1(areg[78]), .z(ain[77]), .d0(areg[77]), .s(x2));
mul_mux2 sh_76_ ( .d1(areg[77]), .z(ain[76]), .d0(areg[76]), .s(x2));
mul_mux2 sh_75_ ( .d1(areg[76]), .z(ain[75]), .d0(areg[75]), .s(x2));
mul_mux2 sh_74_ ( .d1(areg[75]), .z(ain[74]), .d0(areg[74]), .s(x2));
mul_mux2 sh_73_ ( .d1(areg[74]), .z(ain[73]), .d0(areg[73]), .s(x2));
mul_mux2 sh_72_ ( .d1(areg[73]), .z(ain[72]), .d0(areg[72]), .s(x2));
mul_mux2 sh_71_ ( .d1(areg[72]), .z(ain[71]), .d0(areg[71]), .s(x2));
mul_mux2 sh_70_ ( .d1(areg[71]), .z(ain[70]), .d0(areg[70]), .s(x2));
mul_mux2 sh_69_ ( .d1(areg[70]), .z(ain[69]), .d0(areg[69]), .s(x2));
mul_mux2 sh_19_ ( .d1(areg[20]), .z(ain[19]), .d0(areg[19]), .s(x2));
mul_mux2 sh_18_ ( .d1(areg[19]), .z(ain[18]), .d0(areg[18]), .s(x2));
mul_mux2 sh_17_ ( .d1(areg[18]), .z(ain[17]), .d0(areg[17]), .s(x2));
mul_mux2 sh_16_ ( .d1(areg[17]), .z(ain[16]), .d0(areg[16]), .s(x2));
mul_mux2 sh_15_ ( .d1(areg[16]), .z(ain[15]), .d0(areg[15]), .s(x2));
mul_mux2 sh_4_ ( .d1(areg[5]), .z(ain[4]), .d0(areg[4]), .s(x2));
mul_mux2 sh_3_ ( .d1(areg[4]), .z(ain[3]), .d0(areg[3]), .s(x2));
mul_mux2 sh_2_ ( .d1(areg[3]), .z(ain[2]), .d0(areg[2]), .s(x2));
mul_mux2 sh_1_ ( .d1(areg[2]), .z(ain[1]), .d0(areg[1]), .s(x2));
mul_mux2 shx2 ( .d1(areg[0]), .z(ainx2), .d0(1'b0),
     .s(x2));
mul_mux2 sh_83_ ( .d1(areg[84]), .z(ain[83]), .d0(areg[83]), .s(x2));
mul_mux2 sh_14_ ( .d1(areg[15]), .z(ain[14]), .d0(areg[14]), .s(x2));
mul_mux2 sh_13_ ( .d1(areg[14]), .z(ain[13]), .d0(areg[13]), .s(x2));
mul_mux2 sh_12_ ( .d1(areg[13]), .z(ain[12]), .d0(areg[12]), .s(x2));
mul_mux2 sh_11_ ( .d1(areg[12]), .z(ain[11]), .d0(areg[11]), .s(x2));
mul_mux2 sh_10_ ( .d1(areg[11]), .z(ain[10]), .d0(areg[10]), .s(x2));
mul_mux2 sh_9_ ( .d1(areg[10]), .z(ain[9]), .d0(areg[9]), .s(x2));
mul_mux2 sh_8_ ( .d1(areg[9]), .z(ain[8]), .d0(areg[8]), .s(x2));
mul_mux2 sh_7_ ( .d1(areg[8]), .z(ain[7]), .d0(areg[7]), .s(x2));
mul_mux2 sh_6_ ( .d1(areg[7]), .z(ain[6]), .d0(areg[6]), .s(x2));
mul_mux2 sh_5_ ( .d1(areg[6]), .z(ain[5]), .d0(areg[5]), .s(x2));
mul_csa42  sc3_68_ ( .cin(co[67]), .d(1'b0),
     .carry(c3[68]), .c(c2[67]), .b(s2[68]), .a(1'b0),
     .cout(), .sum(s3[68]));
mul_csa42  sc3_67_ ( .cin(co[66]), .d(1'b0),
     .carry(c3[67]), .c(c2[66]), .b(s2[67]), .a(s1[67]), .cout(co[67]),
     .sum(s3[67]));
mul_csa42  sc3_66_ ( .cin(co[65]), .d(c1[65]), .carry(c3[66]),
     .c(c2[65]), .b(s2[66]), .a(s1[66]), .cout(co[66]), .sum(s3[66]));
mul_csa42  sc3_65_ ( .cin(co[64]), .d(c1[64]), .carry(c3[65]),
     .c(c2[64]), .b(s2[65]), .a(s1[65]), .cout(co[65]), .sum(s3[65]));
mul_csa42  sc3_64_ ( .cin(co[63]), .d(c1[63]), .carry(c3[64]),
     .c(c2[63]), .b(s2[64]), .a(s1[64]), .cout(co[64]), .sum(s3[64]));
mul_csa42  sc3_63_ ( .cin(co[62]), .d(c1[62]), .carry(c3[63]),
     .c(c2[62]), .b(s2[63]), .a(s1[63]), .cout(co[63]), .sum(s3[63]));
mul_csa42  sc3_62_ ( .cin(co[61]), .d(c1[61]), .carry(c3[62]),
     .c(c2[61]), .b(s2[62]), .a(s1[62]), .cout(co[62]), .sum(s3[62]));
mul_csa42  sc3_61_ ( .cin(co[60]), .d(c1[60]), .carry(c3[61]),
     .c(c2[60]), .b(s2[61]), .a(s1[61]), .cout(co[61]), .sum(s3[61]));
mul_csa42  sc3_60_ ( .cin(co[59]), .d(c1[59]), .carry(c3[60]),
     .c(c2[59]), .b(s2[60]), .a(s1[60]), .cout(co[60]), .sum(s3[60]));
mul_csa42  sc3_59_ ( .cin(co[58]), .d(c1[58]), .carry(c3[59]),
     .c(c2[58]), .b(s2[59]), .a(s1[59]), .cout(co[59]), .sum(s3[59]));
mul_csa42  sc3_58_ ( .cin(co[57]), .d(c1[57]), .carry(c3[58]),
     .c(c2[57]), .b(s2[58]), .a(s1[58]), .cout(co[58]), .sum(s3[58]));
mul_csa42  sc3_57_ ( .cin(co[56]), .d(c1[56]), .carry(c3[57]),
     .c(c2[56]), .b(s2[57]), .a(s1[57]), .cout(co[57]), .sum(s3[57]));
mul_csa42  sc3_56_ ( .cin(co[55]), .d(c1[55]), .carry(c3[56]),
     .c(c2[55]), .b(s2[56]), .a(s1[56]), .cout(co[56]), .sum(s3[56]));
mul_csa42  sc3_55_ ( .cin(co[54]), .d(c1[54]), .carry(c3[55]),
     .c(c2[54]), .b(s2[55]), .a(s1[55]), .cout(co[55]), .sum(s3[55]));
mul_csa42  sc3_54_ ( .cin(co[53]), .d(c1[53]), .carry(c3[54]),
     .c(c2[53]), .b(s2[54]), .a(s1[54]), .cout(co[54]), .sum(s3[54]));
mul_csa42  sc3_53_ ( .cin(co[52]), .d(c1[52]), .carry(c3[53]),
     .c(c2[52]), .b(s2[53]), .a(s1[53]), .cout(co[53]), .sum(s3[53]));
mul_csa42  sc3_52_ ( .cin(co[51]), .d(c1[51]), .carry(c3[52]),
     .c(c2[51]), .b(s2[52]), .a(s1[52]), .cout(co[52]), .sum(s3[52]));
mul_csa42  sc3_51_ ( .cin(co[50]), .d(c1[50]), .carry(c3[51]),
     .c(c2[50]), .b(s2[51]), .a(s1[51]), .cout(co[51]), .sum(s3[51]));
mul_csa42  sc3_50_ ( .cin(co[49]), .d(c1[49]), .carry(c3[50]),
     .c(c2[49]), .b(s2[50]), .a(s1[50]), .cout(co[50]), .sum(s3[50]));
mul_csa42  sc3_49_ ( .cin(co[48]), .d(c1[48]), .carry(c3[49]),
     .c(c2[48]), .b(s2[49]), .a(s1[49]), .cout(co[49]), .sum(s3[49]));
mul_csa42  sc3_48_ ( .cin(co[47]), .d(c1[47]), .carry(c3[48]),
     .c(c2[47]), .b(s2[48]), .a(s1[48]), .cout(co[48]), .sum(s3[48]));
mul_csa42  sc3_47_ ( .cin(co[46]), .d(c1[46]), .carry(c3[47]),
     .c(c2[46]), .b(s2[47]), .a(s1[47]), .cout(co[47]), .sum(s3[47]));
mul_csa42  sc3_46_ ( .cin(co[45]), .d(c1[45]), .carry(c3[46]),
     .c(c2[45]), .b(s2[46]), .a(s1[46]), .cout(co[46]), .sum(s3[46]));
mul_csa42  sc3_45_ ( .cin(co[44]), .d(c1[44]), .carry(c3[45]),
     .c(c2[44]), .b(s2[45]), .a(s1[45]), .cout(co[45]), .sum(s3[45]));
mul_csa42  sc3_44_ ( .cin(co[43]), .d(c1[43]), .carry(c3[44]),
     .c(c2[43]), .b(s2[44]), .a(s1[44]), .cout(co[44]), .sum(s3[44]));
mul_csa42  sc3_43_ ( .cin(co[42]), .d(c1[42]), .carry(c3[43]),
     .c(c2[42]), .b(s2[43]), .a(s1[43]), .cout(co[43]), .sum(s3[43]));
mul_csa42  sc3_42_ ( .cin(co[41]), .d(c1[41]), .carry(c3[42]),
     .c(c2[41]), .b(s2[42]), .a(s1[42]), .cout(co[42]), .sum(s3[42]));
mul_csa42  sc3_41_ ( .cin(co[40]), .d(c1[40]), .carry(c3[41]),
     .c(c2[40]), .b(s2[41]), .a(s1[41]), .cout(co[41]), .sum(s3[41]));
mul_csa42  sc3_40_ ( .cin(co[39]), .d(c1[39]), .carry(c3[40]),
     .c(c2[39]), .b(s2[40]), .a(s1[40]), .cout(co[40]), .sum(s3[40]));
mul_csa42  sc3_39_ ( .cin(co[38]), .d(c1[38]), .carry(c3[39]),
     .c(c2[38]), .b(s2[39]), .a(s1[39]), .cout(co[39]), .sum(s3[39]));
mul_csa42  sc3_38_ ( .cin(co[37]), .d(c1[37]), .carry(c3[38]),
     .c(c2[37]), .b(s2[38]), .a(s1[38]), .cout(co[38]), .sum(s3[38]));
mul_csa42  sc3_37_ ( .cin(co[36]), .d(c1[36]), .carry(c3[37]),
     .c(c2[36]), .b(s2[37]), .a(s1[37]), .cout(co[37]), .sum(s3[37]));
mul_csa42  sc3_36_ ( .cin(co[35]), .d(c1[35]), .carry(c3[36]),
     .c(c2[35]), .b(s2[36]), .a(s1[36]), .cout(co[36]), .sum(s3[36]));
mul_csa42  sc3_35_ ( .cin(co[34]), .d(c1[34]), .carry(c3[35]),
     .c(c2[34]), .b(s2[35]), .a(s1[35]), .cout(co[35]), .sum(s3[35]));
mul_csa42  sc3_34_ ( .cin(co[33]), .d(c1[33]), .carry(c3[34]),
     .c(c2[33]), .b(s2[34]), .a(s1[34]), .cout(co[34]), .sum(s3[34]));
mul_csa42  sc3_33_ ( .cin(co[32]), .d(c1[32]), .carry(c3[33]),
     .c(c2[32]), .b(s2[33]), .a(s1[33]), .cout(co[33]), .sum(s3[33]));
mul_csa42  sc3_32_ ( .cin(co[31]), .d(c1[31]), .carry(c3[32]),
     .c(c2[31]), .b(s2[32]), .a(s1[32]), .cout(co[32]), .sum(s3[32]));
mul_csa42  sc3_31_ ( .cin(co[30]), .d(c1[30]), .carry(c3[31]),
     .c(c2[30]), .b(s2[31]), .a(s1[31]), .cout(co[31]), .sum(s3[31]));
mul_csa42  sc3_30_ ( .cin(co[29]), .d(c1[29]), .carry(c3[30]),
     .c(c2[29]), .b(s2[30]), .a(s1[30]), .cout(co[30]), .sum(s3[30]));
mul_csa42  sc3_29_ ( .cin(co[28]), .d(c1[28]), .carry(c3[29]),
     .c(c2[28]), .b(s2[29]), .a(s1[29]), .cout(co[29]), .sum(s3[29]));
mul_csa42  sc3_28_ ( .cin(co[27]), .d(c1[27]), .carry(c3[28]),
     .c(c2[27]), .b(s2[28]), .a(s1[28]), .cout(co[28]), .sum(s3[28]));
mul_csa42  sc3_27_ ( .cin(co[26]), .d(c1[26]), .carry(c3[27]),
     .c(c2[26]), .b(s2[27]), .a(s1[27]), .cout(co[27]), .sum(s3[27]));
mul_csa42  sc3_26_ ( .cin(co[25]), .d(c1[25]), .carry(c3[26]),
     .c(c2[25]), .b(s2[26]), .a(s1[26]), .cout(co[26]), .sum(s3[26]));
mul_csa42  sc3_25_ ( .cin(co[24]), .d(c1[24]), .carry(c3[25]),
     .c(c2[24]), .b(s2[25]), .a(s1[25]), .cout(co[25]), .sum(s3[25]));
mul_csa42  sc3_24_ ( .cin(co[23]), .d(c1[23]), .carry(c3[24]),
     .c(c2[23]), .b(s2[24]), .a(s1[24]), .cout(co[24]), .sum(s3[24]));
mul_csa42  sc3_23_ ( .cin(co[22]), .d(c1[22]), .carry(c3[23]),
     .c(c2[22]), .b(s2[23]), .a(s1[23]), .cout(co[23]), .sum(s3[23]));
mul_csa42  sc3_22_ ( .cin(co[21]), .d(c1[21]), .carry(c3[22]),
     .c(c2[21]), .b(s2[22]), .a(s1[22]), .cout(co[22]), .sum(s3[22]));
mul_csa42  sc3_21_ ( .cin(co[20]), .d(c1[20]), .carry(c3[21]),
     .c(c2[20]), .b(s2[21]), .a(s1[21]), .cout(co[21]), .sum(s3[21]));
mul_csa42  sc3_20_ ( .cin(1'b0), .d(c1[19]),
     .carry(c3[20]), .c(c2[19]), .b(s2[20]), .a(s1[20]), .cout(co[20]),
     .sum(s3[20]));
mul_csa32  sc4_82_ ( .c(c3[81]), .b(s2[82]), .a(ain[82]),
     .cout(pcout[82]), .sum(psum[82]));
mul_csa32  sc4_68_ ( .c(c3[67]), .b(s3[68]), .a(ain[68]),
     .cout(pcout[68]), .sum(psum[68]));
mul_csa32  sc4_67_ ( .c(c3[66]), .b(s3[67]), .a(ain[67]),
     .cout(pcout[67]), .sum(psum[67]));
mul_csa32  sc4_66_ ( .c(c3[65]), .b(s3[66]), .a(ain[66]),
     .cout(pcout[66]), .sum(psum[66]));
mul_csa32  sc4_65_ ( .c(c3[64]), .b(s3[65]), .a(ain[65]),
     .cout(pcout[65]), .sum(psum[65]));
mul_csa32  sc4_64_ ( .c(c3[63]), .b(s3[64]), .a(ain[64]),
     .cout(pcout[64]), .sum(psum[64]));
mul_csa32  sc4_63_ ( .c(c3[62]), .b(s3[63]), .a(ain[63]),
     .cout(pcout[63]), .sum(psum[63]));
mul_csa32  sc4_62_ ( .c(c3[61]), .b(s3[62]), .a(ain[62]),
     .cout(pcout[62]), .sum(psum[62]));
mul_csa32  sc4_61_ ( .c(c3[60]), .b(s3[61]), .a(ain[61]),
     .cout(pcout[61]), .sum(psum[61]));
mul_csa32  sc4_60_ ( .c(c3[59]), .b(s3[60]), .a(ain[60]),
     .cout(pcout[60]), .sum(psum[60]));
mul_csa32  sc4_59_ ( .c(c3[58]), .b(s3[59]), .a(ain[59]),
     .cout(pcout[59]), .sum(psum[59]));
mul_csa32  sc4_58_ ( .c(c3[57]), .b(s3[58]), .a(ain[58]),
     .cout(pcout[58]), .sum(psum[58]));
mul_csa32  sc4_57_ ( .c(c3[56]), .b(s3[57]), .a(ain[57]),
     .cout(pcout[57]), .sum(psum[57]));
mul_csa32  sc4_56_ ( .c(c3[55]), .b(s3[56]), .a(ain[56]),
     .cout(pcout[56]), .sum(psum[56]));
mul_csa32  sc4_55_ ( .c(c3[54]), .b(s3[55]), .a(ain[55]),
     .cout(pcout[55]), .sum(psum[55]));
mul_csa32  sc4_54_ ( .c(c3[53]), .b(s3[54]), .a(ain[54]),
     .cout(pcout[54]), .sum(psum[54]));
mul_csa32  sc4_53_ ( .c(c3[52]), .b(s3[53]), .a(ain[53]),
     .cout(pcout[53]), .sum(psum[53]));
mul_csa32  sc4_52_ ( .c(c3[51]), .b(s3[52]), .a(ain[52]),
     .cout(pcout[52]), .sum(psum[52]));
mul_csa32  sc4_51_ ( .c(c3[50]), .b(s3[51]), .a(ain[51]),
     .cout(pcout[51]), .sum(psum[51]));
mul_csa32  sc4_50_ ( .c(c3[49]), .b(s3[50]), .a(ain[50]),
     .cout(pcout[50]), .sum(psum[50]));
mul_csa32  sc4_49_ ( .c(c3[48]), .b(s3[49]), .a(ain[49]),
     .cout(pcout[49]), .sum(psum[49]));
mul_csa32  sc4_48_ ( .c(c3[47]), .b(s3[48]), .a(ain[48]),
     .cout(pcout[48]), .sum(psum[48]));
mul_csa32  sc4_47_ ( .c(c3[46]), .b(s3[47]), .a(ain[47]),
     .cout(pcout[47]), .sum(psum[47]));
mul_csa32  sc4_46_ ( .c(c3[45]), .b(s3[46]), .a(ain[46]),
     .cout(pcout[46]), .sum(psum[46]));
mul_csa32  sc4_45_ ( .c(c3[44]), .b(s3[45]), .a(ain[45]),
     .cout(pcout[45]), .sum(psum[45]));
mul_csa32  sc4_44_ ( .c(c3[43]), .b(s3[44]), .a(ain[44]),
     .cout(pcout[44]), .sum(psum[44]));
mul_csa32  sc4_43_ ( .c(c3[42]), .b(s3[43]), .a(ain[43]),
     .cout(pcout[43]), .sum(psum[43]));
mul_csa32  sc4_42_ ( .c(c3[41]), .b(s3[42]), .a(ain[42]),
     .cout(pcout[42]), .sum(psum[42]));
mul_csa32  sc4_41_ ( .c(c3[40]), .b(s3[41]), .a(ain[41]),
     .cout(pcout[41]), .sum(psum[41]));
mul_csa32  sc4_40_ ( .c(c3[39]), .b(s3[40]), .a(ain[40]),
     .cout(pcout[40]), .sum(psum[40]));
mul_csa32  sc4_39_ ( .c(c3[38]), .b(s3[39]), .a(ain[39]),
     .cout(pcout[39]), .sum(psum[39]));
mul_csa32  sc4_38_ ( .c(c3[37]), .b(s3[38]), .a(ain[38]),
     .cout(pcout[38]), .sum(psum[38]));
mul_csa32  sc4_37_ ( .c(c3[36]), .b(s3[37]), .a(ain[37]),
     .cout(pcout[37]), .sum(psum[37]));
mul_csa32  sc4_36_ ( .c(c3[35]), .b(s3[36]), .a(ain[36]),
     .cout(pcout[36]), .sum(psum[36]));
mul_csa32  sc4_35_ ( .c(c3[34]), .b(s3[35]), .a(ain[35]),
     .cout(pcout[35]), .sum(psum[35]));
mul_csa32  sc4_34_ ( .c(c3[33]), .b(s3[34]), .a(ain[34]),
     .cout(pcout[34]), .sum(psum[34]));
mul_csa32  sc4_33_ ( .c(c3[32]), .b(s3[33]), .a(ain[33]),
     .cout(pcout[33]), .sum(psum[33]));
mul_csa32  sc4_32_ ( .c(c3[31]), .b(s3[32]), .a(ain[32]),
     .cout(pcout[32]), .sum(psum[32]));
mul_csa32  sc4_31_ ( .c(c3[30]), .b(s3[31]), .a(ain[31]),
     .cout(pcout[31]), .sum(psum[31]));
mul_csa32  sc4_30_ ( .c(c3[29]), .b(s3[30]), .a(ain[30]),
     .cout(pcout[30]), .sum(psum[30]));
mul_csa32  sc4_29_ ( .c(c3[28]), .b(s3[29]), .a(ain[29]),
     .cout(pcout[29]), .sum(psum[29]));
mul_csa32  sc4_28_ ( .c(c3[27]), .b(s3[28]), .a(ain[28]),
     .cout(pcout[28]), .sum(psum[28]));
mul_csa32  sc4_27_ ( .c(c3[26]), .b(s3[27]), .a(ain[27]),
     .cout(pcout[27]), .sum(psum[27]));
mul_csa32  sc4_26_ ( .c(c3[25]), .b(s3[26]), .a(ain[26]),
     .cout(pcout[26]), .sum(psum[26]));
mul_csa32  sc4_25_ ( .c(c3[24]), .b(s3[25]), .a(ain[25]),
     .cout(pcout[25]), .sum(psum[25]));
mul_csa32  sc4_24_ ( .c(c3[23]), .b(s3[24]), .a(ain[24]),
     .cout(pcout[24]), .sum(psum[24]));
mul_csa32  sc4_23_ ( .c(c3[22]), .b(s3[23]), .a(ain[23]),
     .cout(pcout[23]), .sum(psum[23]));
mul_csa32  sc4_22_ ( .c(c3[21]), .b(s3[22]), .a(ain[22]),
     .cout(pcout[22]), .sum(psum[22]));
mul_csa32  sc4_21_ ( .c(c3[20]), .b(s3[21]), .a(ain[21]),
     .cout(pcout[21]), .sum(psum[21]));
mul_csa32  sc4_20_ ( .c(c3[19]), .b(s3[20]), .a(ain[20]),
     .cout(pcout[20]), .sum(psum[20]));
mul_csa32  sc4_96_ ( .c(c2[95]), .b(s2[96]), .a(ain[96]),
     .cout(pcout[96]), .sum(psum[96]));
mul_csa32  sc4_95_ ( .c(c2[94]), .b(s2[95]), .a(ain[95]),
     .cout(pcout[95]), .sum(psum[95]));
mul_csa32  sc4_94_ ( .c(c2[93]), .b(s2[94]), .a(ain[94]),
     .cout(pcout[94]), .sum(psum[94]));
mul_csa32  sc4_93_ ( .c(c2[92]), .b(s2[93]), .a(ain[93]),
     .cout(pcout[93]), .sum(psum[93]));
mul_csa32  sc4_92_ ( .c(c2[91]), .b(s2[92]), .a(ain[92]),
     .cout(pcout[92]), .sum(psum[92]));
mul_csa32  sc4_91_ ( .c(c2[90]), .b(s2[91]), .a(ain[91]),
     .cout(pcout[91]), .sum(psum[91]));
mul_csa32  sc4_90_ ( .c(c2[89]), .b(s2[90]), .a(ain[90]),
     .cout(pcout[90]), .sum(psum[90]));
mul_csa32  sc4_89_ ( .c(c2[88]), .b(s2[89]), .a(ain[89]),
     .cout(pcout[89]), .sum(psum[89]));
mul_csa32  sc4_88_ ( .c(c2[87]), .b(s2[88]), .a(ain[88]),
     .cout(pcout[88]), .sum(psum[88]));
mul_csa32  sc4_87_ ( .c(c2[86]), .b(s2[87]), .a(ain[87]),
     .cout(pcout[87]), .sum(psum[87]));
mul_csa32  sc4_86_ ( .c(c2[85]), .b(s2[86]), .a(ain[86]),
     .cout(pcout[86]), .sum(psum[86]));
mul_csa32  sc4_85_ ( .c(c2[84]), .b(s2[85]), .a(ain[85]),
     .cout(pcout[85]), .sum(psum[85]));
mul_csa32  sc4_84_ ( .c(c2[83]), .b(s2[84]), .a(ain[84]),
     .cout(pcout[84]), .sum(psum[84]));
mul_csa32  sc4_81_ ( .c(c3[80]), .b(s3[81]), .a(ain[81]),
     .cout(pcout[81]), .sum(psum[81]));
mul_csa32  sc4_80_ ( .c(c3[79]), .b(s3[80]), .a(ain[80]),
     .cout(pcout[80]), .sum(psum[80]));
mul_csa32  sc4_79_ ( .c(c3[78]), .b(s3[79]), .a(ain[79]),
     .cout(pcout[79]), .sum(psum[79]));
mul_csa32  sc4_78_ ( .c(c3[77]), .b(s3[78]), .a(ain[78]),
     .cout(pcout[78]), .sum(psum[78]));
mul_csa32  sc4_77_ ( .c(c3[76]), .b(s3[77]), .a(ain[77]),
     .cout(pcout[77]), .sum(psum[77]));
mul_csa32  sc4_76_ ( .c(c3[75]), .b(s3[76]), .a(ain[76]),
     .cout(pcout[76]), .sum(psum[76]));
mul_csa32  sc4_75_ ( .c(c3[74]), .b(s3[75]), .a(ain[75]),
     .cout(pcout[75]), .sum(psum[75]));
mul_csa32  sc4_74_ ( .c(c3[73]), .b(s3[74]), .a(ain[74]),
     .cout(pcout[74]), .sum(psum[74]));
mul_csa32  sc4_73_ ( .c(c3[72]), .b(s3[73]), .a(ain[73]),
     .cout(pcout[73]), .sum(psum[73]));
mul_csa32  sc4_72_ ( .c(c3[71]), .b(s3[72]), .a(ain[72]),
     .cout(pcout[72]), .sum(psum[72]));
mul_csa32  sc4_71_ ( .c(c3[70]), .b(s3[71]), .a(ain[71]),
     .cout(pcout[71]), .sum(psum[71]));
mul_csa32  sc4_70_ ( .c(c3[69]), .b(s3[70]), .a(ain[70]),
     .cout(pcout[70]), .sum(psum[70]));
mul_csa32  sc4_69_ ( .c(c3[68]), .b(s3[69]), .a(ain[69]),
     .cout(pcout[69]), .sum(psum[69]));
mul_csa32  acc_4_ ( .c(c2[3]), .sum(psum[4]), .cout(pcout[4]),
     .a(ain[4]), .b(s2[4]));
mul_csa32  acc_3_ ( .c(c2[2]), .sum(psum[3]), .cout(pcout[3]),
     .a(ain[3]), .b(s2[3]));
mul_csa32  acc_2_ ( .c(c2[1]), .sum(psum[2]), .cout(pcout[2]),
     .a(ain[2]), .b(s2[2]));
mul_csa32  acc_1_ ( .c(c2[0]), .sum(psum[1]), .cout(pcout[1]),
     .a(ain[1]), .b(s2[1]));
mul_csa32  sc3_97_ ( .c(c2[96]), .sum(psum[97]), .cout(pcout[97]),
     .a(a1s[81]), .b(a1c[80]));
mul_csa32  sc1_19_ ( .c(a1s[3]), .b(pc[50]), .a(ps[51]),
     .cout(c1[19]), .sum(s1[19]));
mul_csa32  sc1_18_ ( .c(a1s[2]), .b(pc[49]), .a(ps[50]),
     .cout(c1[18]), .sum(s1[18]));
mul_csa32  sc1_17_ ( .c(a1s[1]), .b(pc[48]), .a(ps[49]),
     .cout(c1[17]), .sum(s1[17]));
mul_csa32  sc1_16_ ( .c(a1s[0]), .b(pc[47]), .a(ps[48]),
     .cout(c1[16]), .sum(s1[16]));
mul_csa32  sc1_15_ ( .c(1'b0), .b(pc[46]), .a(ps[47]),
     .cout(c1[15]), .sum(s1[15]));
mul_csa32  sc4_83_ ( .c(c2[82]), .b(s2[83]), .a(ain[83]),
     .cout(pcout[83]), .sum(psum[83]));
mul_csa32  sc2_83_ ( .c(c1[82]), .b(a1c[66]), .a(a1s[67]),
     .cout(c2[83]), .sum(s2[83]));
mul_csa32  sc2_19_ ( .c(a0c[18]), .b(a0s[19]), .a(s1[19]),
     .cout(c2[19]), .sum(s2[19]));
mul_csa32  sc2_18_ ( .c(a0c[17]), .b(a0s[18]), .a(s1[18]),
     .cout(c2[18]), .sum(s2[18]));
mul_csa32  sc2_17_ ( .c(a0c[16]), .b(a0s[17]), .a(s1[17]),
     .cout(c2[17]), .sum(s2[17]));
mul_csa32  sc2_16_ ( .c(a0c[15]), .b(a0s[16]), .a(s1[16]),
     .cout(c2[16]), .sum(s2[16]));
mul_csa32  sc2_15_ ( .c(a0c[14]), .b(a0s[15]), .a(s1[15]),
     .cout(c2[15]), .sum(s2[15]));
mul_csa32  sc1_81_ ( .c(a0s[81]), .b(a1c[64]), .a(a1s[65]),
     .cout(c1[81]), .sum(s1[81]));
mul_csa32  sc1_80_ ( .c(a0s[80]), .b(a1c[63]), .a(a1s[64]),
     .cout(c1[80]), .sum(s1[80]));
mul_csa32  sc1_79_ ( .c(a0s[79]), .b(a1c[62]), .a(a1s[63]),
     .cout(c1[79]), .sum(s1[79]));
mul_csa32  sc1_78_ ( .c(a0s[78]), .b(a1c[61]), .a(a1s[62]),
     .cout(c1[78]), .sum(s1[78]));
mul_csa32  sc1_77_ ( .c(a0s[77]), .b(a1c[60]), .a(a1s[61]),
     .cout(c1[77]), .sum(s1[77]));
mul_csa32  sc1_76_ ( .c(a0s[76]), .b(a1c[59]), .a(a1s[60]),
     .cout(c1[76]), .sum(s1[76]));
mul_csa32  sc1_75_ ( .c(a0s[75]), .b(a1c[58]), .a(a1s[59]),
     .cout(c1[75]), .sum(s1[75]));
mul_csa32  sc1_74_ ( .c(a0s[74]), .b(a1c[57]), .a(a1s[58]),
     .cout(c1[74]), .sum(s1[74]));
mul_csa32  sc1_73_ ( .c(a0s[73]), .b(a1c[56]), .a(a1s[57]),
     .cout(c1[73]), .sum(s1[73]));
mul_csa32  sc1_72_ ( .c(a0s[72]), .b(a1c[55]), .a(a1s[56]),
     .cout(c1[72]), .sum(s1[72]));
mul_csa32  sc1_71_ ( .c(a0s[71]), .b(a1c[54]), .a(a1s[55]),
     .cout(c1[71]), .sum(s1[71]));
mul_csa32  sc1_70_ ( .c(a0s[70]), .b(a1c[53]), .a(a1s[54]),
     .cout(c1[70]), .sum(s1[70]));
mul_csa32  sc1_69_ ( .c(a0s[69]), .b(a1c[52]), .a(a1s[53]),
     .cout(c1[69]), .sum(s1[69]));
mul_csa32  sc1_68_ ( .c(a0s[68]), .b(a1c[51]), .a(a1s[52]),
     .cout(c1[68]), .sum(s1[68]));
mul_csa32  sc3_19_ ( .c(c2[18]), .b(c1[18]), .a(s2[19]),
     .cout(c3[19]), .sum(s3[19]));
mul_csa32  sc3_18_ ( .c(c2[17]), .b(c1[17]), .a(s2[18]),
     .cout(c3[18]), .sum(s3[18]));
mul_csa32  sc3_17_ ( .c(c2[16]), .b(c1[16]), .a(s2[17]),
     .cout(c3[17]), .sum(s3[17]));
mul_csa32  sc3_16_ ( .c(c2[15]), .b(c1[15]), .a(s2[16]),
     .cout(c3[16]), .sum(s3[16]));
mul_csa32  sc3_15_ ( .c(c2[14]), .b(c1[14]), .a(s2[15]),
     .cout(c3[15]), .sum(s3[15]));
mul_csa32  sc1_82_ ( .c(a0c[81]), .b(a1c[65]), .a(a1s[66]),
     .cout(c1[82]), .sum(s1[82]));
mul_csa32  acc_14_ ( .c(c2[13]), .sum(psum[14]), .cout(pcout[14]),
     .a(ain[14]), .b(s2[14]));
mul_csa32  acc_13_ ( .c(c2[12]), .sum(psum[13]), .cout(pcout[13]),
     .a(ain[13]), .b(s2[13]));
mul_csa32  acc_12_ ( .c(c2[11]), .sum(psum[12]), .cout(pcout[12]),
     .a(ain[12]), .b(s2[12]));
mul_csa32  acc_11_ ( .c(c2[10]), .sum(psum[11]), .cout(pcout[11]),
     .a(ain[11]), .b(s2[11]));
mul_csa32  acc_10_ ( .c(c2[9]), .sum(psum[10]), .cout(pcout[10]),
     .a(ain[10]), .b(s2[10]));
mul_csa32  acc_9_ ( .c(c2[8]), .sum(psum[9]), .cout(pcout[9]),
     .a(ain[9]), .b(s2[9]));
mul_csa32  acc_8_ ( .c(c2[7]), .sum(psum[8]), .cout(pcout[8]),
     .a(ain[8]), .b(s2[8]));
mul_csa32  acc_7_ ( .c(c2[6]), .sum(psum[7]), .cout(pcout[7]),
     .a(ain[7]), .b(s2[7]));
mul_csa32  acc_6_ ( .c(c2[5]), .sum(psum[6]), .cout(pcout[6]),
     .a(ain[6]), .b(s2[6]));
mul_csa32  acc_5_ ( .c(c2[4]), .sum(psum[5]), .cout(pcout[5]),
     .a(ain[5]), .b(s2[5]));
mul_csa32  sc2_67_ ( .c(a0c[66]), .b(c1[66]), .a(a0s[67]),
     .cout(c2[67]), .sum(s2[67]));
mul_csa32  sc1_14_ ( .c(a0s[14]), .b(pc[45]), .a(ps[46]),
     .cout(c1[14]), .sum(s1[14]));
mul_csa32  sc1_13_ ( .c(a0s[13]), .b(pc[44]), .a(ps[45]),
     .cout(c1[13]), .sum(s1[13]));
mul_csa32  sc1_12_ ( .c(a0s[12]), .b(pc[43]), .a(ps[44]),
     .cout(c1[12]), .sum(s1[12]));
mul_csa32  sc1_11_ ( .c(a0s[11]), .b(pc[42]), .a(ps[43]),
     .cout(c1[11]), .sum(s1[11]));
mul_csa32  sc1_10_ ( .c(a0s[10]), .b(pc[41]), .a(ps[42]),
     .cout(c1[10]), .sum(s1[10]));
mul_csa32  sc1_9_ ( .c(a0s[9]), .b(pc[40]), .a(ps[41]), .cout(c1[9]),
     .sum(s1[9]));
mul_csa32  sc1_8_ ( .c(a0s[8]), .b(pc[39]), .a(ps[40]), .cout(c1[8]),
     .sum(s1[8]));
mul_csa32  sc1_7_ ( .c(a0s[7]), .b(pc[38]), .a(ps[39]), .cout(c1[7]),
     .sum(s1[7]));
mul_csa32  sc1_6_ ( .c(a0s[6]), .b(pc[37]), .a(ps[38]), .cout(c1[6]),
     .sum(s1[6]));
mul_csa32  sc1_5_ ( .c(a0s[5]), .b(pc[36]), .a(ps[37]), .cout(c1[5]),
     .sum(s1[5]));
mul_csa32  sc2_14_ ( .c(a0c[13]), .b(c1[13]), .a(s1[14]),
     .cout(c2[14]), .sum(s2[14]));
mul_csa32  sc2_13_ ( .c(a0c[12]), .b(c1[12]), .a(s1[13]),
     .cout(c2[13]), .sum(s2[13]));
mul_csa32  sc2_12_ ( .c(a0c[11]), .b(c1[11]), .a(s1[12]),
     .cout(c2[12]), .sum(s2[12]));
mul_csa32  sc2_11_ ( .c(a0c[10]), .b(c1[10]), .a(s1[11]),
     .cout(c2[11]), .sum(s2[11]));
mul_csa32  sc2_10_ ( .c(a0c[9]), .b(c1[9]), .a(s1[10]),
     .cout(c2[10]), .sum(s2[10]));
mul_csa32  sc2_9_ ( .c(a0c[8]), .b(c1[8]), .a(s1[9]), .cout(c2[9]),
     .sum(s2[9]));
mul_csa32  sc2_8_ ( .c(a0c[7]), .b(c1[7]), .a(s1[8]), .cout(c2[8]),
     .sum(s2[8]));
mul_csa32  sc2_7_ ( .c(a0c[6]), .b(c1[6]), .a(s1[7]), .cout(c2[7]),
     .sum(s2[7]));
mul_csa32  sc2_6_ ( .c(a0c[5]), .b(c1[5]), .a(s1[6]), .cout(c2[6]),
     .sum(s2[6]));
mul_csa32  sc2_5_ ( .c(a0c[4]), .b(c1[4]), .a(s1[5]), .cout(c2[5]),
     .sum(s2[5]));
mul_csa32  sc2_82_ ( .c(c2[81]), .b(c1[81]), .a(s1[82]),
     .cout(c2[82]), .sum(s2[82]));
mul_csa32  sc1_4_ ( .c(a0s[4]), .b(pc[35]), .a(ps[36]), .cout(c1[4]),
     .sum(s1[4]));
mul_csa32  sc1_3_ ( .c(a0s[3]), .b(pc[34]), .a(ps[35]), .cout(c1[3]),
     .sum(s1[3]));
mul_csa32  sc1_2_ ( .c(a0s[2]), .b(pc[33]), .a(ps[34]), .cout(c1[2]),
     .sum(s1[2]));
mul_csa32  sc1_1_ ( .c(a0s[1]), .b(pc[32]), .a(ps[33]), .cout(c1[1]),
     .sum(s1[1]));
mul_csa32  sc2_66_ ( .c(a0c[65]), .b(a0s[66]), .a(a1c[49]),
     .cout(c2[66]), .sum(s2[66]));
mul_csa32  sc2_65_ ( .c(a0c[64]), .b(a0s[65]), .a(a1c[48]),
     .cout(c2[65]), .sum(s2[65]));
mul_csa32  sc2_64_ ( .c(a0c[63]), .b(a0s[64]), .a(a1c[47]),
     .cout(c2[64]), .sum(s2[64]));
mul_csa32  sc2_63_ ( .c(a0c[62]), .b(a0s[63]), .a(a1c[46]),
     .cout(c2[63]), .sum(s2[63]));
mul_csa32  sc2_62_ ( .c(a0c[61]), .b(a0s[62]), .a(a1c[45]),
     .cout(c2[62]), .sum(s2[62]));
mul_csa32  sc2_61_ ( .c(a0c[60]), .b(a0s[61]), .a(a1c[44]),
     .cout(c2[61]), .sum(s2[61]));
mul_csa32  sc2_60_ ( .c(a0c[59]), .b(a0s[60]), .a(a1c[43]),
     .cout(c2[60]), .sum(s2[60]));
mul_csa32  sc2_59_ ( .c(a0c[58]), .b(a0s[59]), .a(a1c[42]),
     .cout(c2[59]), .sum(s2[59]));
mul_csa32  sc2_58_ ( .c(a0c[57]), .b(a0s[58]), .a(a1c[41]),
     .cout(c2[58]), .sum(s2[58]));
mul_csa32  sc2_57_ ( .c(a0c[56]), .b(a0s[57]), .a(a1c[40]),
     .cout(c2[57]), .sum(s2[57]));
mul_csa32  sc2_56_ ( .c(a0c[55]), .b(a0s[56]), .a(a1c[39]),
     .cout(c2[56]), .sum(s2[56]));
mul_csa32  sc2_55_ ( .c(a0c[54]), .b(a0s[55]), .a(a1c[38]),
     .cout(c2[55]), .sum(s2[55]));
mul_csa32  sc2_54_ ( .c(a0c[53]), .b(a0s[54]), .a(a1c[37]),
     .cout(c2[54]), .sum(s2[54]));
mul_csa32  sc2_53_ ( .c(a0c[52]), .b(a0s[53]), .a(a1c[36]),
     .cout(c2[53]), .sum(s2[53]));
mul_csa32  sc2_52_ ( .c(a0c[51]), .b(a0s[52]), .a(a1c[35]),
     .cout(c2[52]), .sum(s2[52]));
mul_csa32  sc2_51_ ( .c(a0c[50]), .b(a0s[51]), .a(a1c[34]),
     .cout(c2[51]), .sum(s2[51]));
mul_csa32  sc2_50_ ( .c(a0c[49]), .b(a0s[50]), .a(a1c[33]),
     .cout(c2[50]), .sum(s2[50]));
mul_csa32  sc2_49_ ( .c(a0c[48]), .b(a0s[49]), .a(a1c[32]),
     .cout(c2[49]), .sum(s2[49]));
mul_csa32  sc2_48_ ( .c(a0c[47]), .b(a0s[48]), .a(a1c[31]),
     .cout(c2[48]), .sum(s2[48]));
mul_csa32  sc2_47_ ( .c(a0c[46]), .b(a0s[47]), .a(a1c[30]),
     .cout(c2[47]), .sum(s2[47]));
mul_csa32  sc2_46_ ( .c(a0c[45]), .b(a0s[46]), .a(a1c[29]),
     .cout(c2[46]), .sum(s2[46]));
mul_csa32  sc2_45_ ( .c(a0c[44]), .b(a0s[45]), .a(a1c[28]),
     .cout(c2[45]), .sum(s2[45]));
mul_csa32  sc2_44_ ( .c(a0c[43]), .b(a0s[44]), .a(a1c[27]),
     .cout(c2[44]), .sum(s2[44]));
mul_csa32  sc2_43_ ( .c(a0c[42]), .b(a0s[43]), .a(a1c[26]),
     .cout(c2[43]), .sum(s2[43]));
mul_csa32  sc2_42_ ( .c(a0c[41]), .b(a0s[42]), .a(a1c[25]),
     .cout(c2[42]), .sum(s2[42]));
mul_csa32  sc2_41_ ( .c(a0c[40]), .b(a0s[41]), .a(a1c[24]),
     .cout(c2[41]), .sum(s2[41]));
mul_csa32  sc2_40_ ( .c(a0c[39]), .b(a0s[40]), .a(a1c[23]),
     .cout(c2[40]), .sum(s2[40]));
mul_csa32  sc2_39_ ( .c(a0c[38]), .b(a0s[39]), .a(a1c[22]),
     .cout(c2[39]), .sum(s2[39]));
mul_csa32  sc2_38_ ( .c(a0c[37]), .b(a0s[38]), .a(a1c[21]),
     .cout(c2[38]), .sum(s2[38]));
mul_csa32  sc2_37_ ( .c(a0c[36]), .b(a0s[37]), .a(a1c[20]),
     .cout(c2[37]), .sum(s2[37]));
mul_csa32  sc2_36_ ( .c(a0c[35]), .b(a0s[36]), .a(a1c[19]),
     .cout(c2[36]), .sum(s2[36]));
mul_csa32  sc2_35_ ( .c(a0c[34]), .b(a0s[35]), .a(a1c[18]),
     .cout(c2[35]), .sum(s2[35]));
mul_csa32  sc2_34_ ( .c(a0c[33]), .b(a0s[34]), .a(a1c[17]),
     .cout(c2[34]), .sum(s2[34]));
mul_csa32  sc2_33_ ( .c(a0c[32]), .b(a0s[33]), .a(a1c[16]),
     .cout(c2[33]), .sum(s2[33]));
mul_csa32  sc2_32_ ( .c(a0c[31]), .b(a0s[32]), .a(a1c[15]),
     .cout(c2[32]), .sum(s2[32]));
mul_csa32  sc2_31_ ( .c(a0c[30]), .b(a0s[31]), .a(a1c[14]),
     .cout(c2[31]), .sum(s2[31]));
mul_csa32  sc2_30_ ( .c(a0c[29]), .b(a0s[30]), .a(a1c[13]),
     .cout(c2[30]), .sum(s2[30]));
mul_csa32  sc2_29_ ( .c(a0c[28]), .b(a0s[29]), .a(a1c[12]),
     .cout(c2[29]), .sum(s2[29]));
mul_csa32  sc2_28_ ( .c(a0c[27]), .b(a0s[28]), .a(a1c[11]),
     .cout(c2[28]), .sum(s2[28]));
mul_csa32  sc2_27_ ( .c(a0c[26]), .b(a0s[27]), .a(a1c[10]),
     .cout(c2[27]), .sum(s2[27]));
mul_csa32  sc2_26_ ( .c(a0c[25]), .b(a0s[26]), .a(a1c[9]),
     .cout(c2[26]), .sum(s2[26]));
mul_csa32  sc2_25_ ( .c(a0c[24]), .b(a0s[25]), .a(a1c[8]),
     .cout(c2[25]), .sum(s2[25]));
mul_csa32  sc2_24_ ( .c(a0c[23]), .b(a0s[24]), .a(a1c[7]),
     .cout(c2[24]), .sum(s2[24]));
mul_csa32  sc2_23_ ( .c(a0c[22]), .b(a0s[23]), .a(a1c[6]),
     .cout(c2[23]), .sum(s2[23]));
mul_csa32  sc2_22_ ( .c(a0c[21]), .b(a0s[22]), .a(a1c[5]),
     .cout(c2[22]), .sum(s2[22]));
mul_csa32  sc2_21_ ( .c(a0c[20]), .b(a0s[21]), .a(a1c[4]),
     .cout(c2[21]), .sum(s2[21]));
mul_csa32  sc2_20_ ( .c(a0c[19]), .b(a0s[20]), .a(1'b0),
     .cout(c2[20]), .sum(s2[20]));
mul_csa32  sc1_66_ ( .c(a1s[50]), .b(pc[97]), .a(ps[98]),
     .cout(c1[66]), .sum(s1[66]));
mul_csa32  sc1_65_ ( .c(a1s[49]), .b(pc[96]), .a(ps[97]),
     .cout(c1[65]), .sum(s1[65]));
mul_csa32  sc1_64_ ( .c(a1s[48]), .b(pc[95]), .a(ps[96]),
     .cout(c1[64]), .sum(s1[64]));
mul_csa32  sc1_63_ ( .c(a1s[47]), .b(pc[94]), .a(ps[95]),
     .cout(c1[63]), .sum(s1[63]));
mul_csa32  sc1_62_ ( .c(a1s[46]), .b(pc[93]), .a(ps[94]),
     .cout(c1[62]), .sum(s1[62]));
mul_csa32  sc1_61_ ( .c(a1s[45]), .b(pc[92]), .a(ps[93]),
     .cout(c1[61]), .sum(s1[61]));
mul_csa32  sc1_60_ ( .c(a1s[44]), .b(pc[91]), .a(ps[92]),
     .cout(c1[60]), .sum(s1[60]));
mul_csa32  sc1_59_ ( .c(a1s[43]), .b(pc[90]), .a(ps[91]),
     .cout(c1[59]), .sum(s1[59]));
mul_csa32  sc1_58_ ( .c(a1s[42]), .b(pc[89]), .a(ps[90]),
     .cout(c1[58]), .sum(s1[58]));
mul_csa32  sc1_57_ ( .c(a1s[41]), .b(pc[88]), .a(ps[89]),
     .cout(c1[57]), .sum(s1[57]));
mul_csa32  sc1_56_ ( .c(a1s[40]), .b(pc[87]), .a(ps[88]),
     .cout(c1[56]), .sum(s1[56]));
mul_csa32  sc1_55_ ( .c(a1s[39]), .b(pc[86]), .a(ps[87]),
     .cout(c1[55]), .sum(s1[55]));
mul_csa32  sc1_54_ ( .c(a1s[38]), .b(pc[85]), .a(ps[86]),
     .cout(c1[54]), .sum(s1[54]));
mul_csa32  sc1_53_ ( .c(a1s[37]), .b(pc[84]), .a(ps[85]),
     .cout(c1[53]), .sum(s1[53]));
mul_csa32  sc1_52_ ( .c(a1s[36]), .b(pc[83]), .a(ps[84]),
     .cout(c1[52]), .sum(s1[52]));
mul_csa32  sc1_51_ ( .c(a1s[35]), .b(pc[82]), .a(ps[83]),
     .cout(c1[51]), .sum(s1[51]));
mul_csa32  sc1_50_ ( .c(a1s[34]), .b(pc[81]), .a(ps[82]),
     .cout(c1[50]), .sum(s1[50]));
mul_csa32  sc1_49_ ( .c(a1s[33]), .b(pc[80]), .a(ps[81]),
     .cout(c1[49]), .sum(s1[49]));
mul_csa32  sc1_48_ ( .c(a1s[32]), .b(pc[79]), .a(ps[80]),
     .cout(c1[48]), .sum(s1[48]));
mul_csa32  sc1_47_ ( .c(a1s[31]), .b(pc[78]), .a(ps[79]),
     .cout(c1[47]), .sum(s1[47]));
mul_csa32  sc1_46_ ( .c(a1s[30]), .b(pc[77]), .a(ps[78]),
     .cout(c1[46]), .sum(s1[46]));
mul_csa32  sc1_45_ ( .c(a1s[29]), .b(pc[76]), .a(ps[77]),
     .cout(c1[45]), .sum(s1[45]));
mul_csa32  sc1_44_ ( .c(a1s[28]), .b(pc[75]), .a(ps[76]),
     .cout(c1[44]), .sum(s1[44]));
mul_csa32  sc1_43_ ( .c(a1s[27]), .b(pc[74]), .a(ps[75]),
     .cout(c1[43]), .sum(s1[43]));
mul_csa32  sc1_42_ ( .c(a1s[26]), .b(pc[73]), .a(ps[74]),
     .cout(c1[42]), .sum(s1[42]));
mul_csa32  sc1_41_ ( .c(a1s[25]), .b(pc[72]), .a(ps[73]),
     .cout(c1[41]), .sum(s1[41]));
mul_csa32  sc1_40_ ( .c(a1s[24]), .b(pc[71]), .a(ps[72]),
     .cout(c1[40]), .sum(s1[40]));
mul_csa32  sc1_39_ ( .c(a1s[23]), .b(pc[70]), .a(ps[71]),
     .cout(c1[39]), .sum(s1[39]));
mul_csa32  sc1_38_ ( .c(a1s[22]), .b(pc[69]), .a(ps[70]),
     .cout(c1[38]), .sum(s1[38]));
mul_csa32  sc1_37_ ( .c(a1s[21]), .b(pc[68]), .a(ps[69]),
     .cout(c1[37]), .sum(s1[37]));
mul_csa32  sc1_36_ ( .c(a1s[20]), .b(pc[67]), .a(ps[68]),
     .cout(c1[36]), .sum(s1[36]));
mul_csa32  sc1_35_ ( .c(a1s[19]), .b(pc[66]), .a(ps[67]),
     .cout(c1[35]), .sum(s1[35]));
mul_csa32  sc1_34_ ( .c(a1s[18]), .b(pc[65]), .a(ps[66]),
     .cout(c1[34]), .sum(s1[34]));
mul_csa32  sc1_33_ ( .c(a1s[17]), .b(pc[64]), .a(ps[65]),
     .cout(c1[33]), .sum(s1[33]));
mul_csa32  sc1_32_ ( .c(a1s[16]), .b(pc[63]), .a(ps[64]),
     .cout(c1[32]), .sum(s1[32]));
mul_csa32  sc1_31_ ( .c(a1s[15]), .b(pc[62]), .a(ps[63]),
     .cout(c1[31]), .sum(s1[31]));
mul_csa32  sc1_30_ ( .c(a1s[14]), .b(pc[61]), .a(ps[62]),
     .cout(c1[30]), .sum(s1[30]));
mul_csa32  sc1_29_ ( .c(a1s[13]), .b(pc[60]), .a(ps[61]),
     .cout(c1[29]), .sum(s1[29]));
mul_csa32  sc1_28_ ( .c(a1s[12]), .b(pc[59]), .a(ps[60]),
     .cout(c1[28]), .sum(s1[28]));
mul_csa32  sc1_27_ ( .c(a1s[11]), .b(pc[58]), .a(ps[59]),
     .cout(c1[27]), .sum(s1[27]));
mul_csa32  sc1_26_ ( .c(a1s[10]), .b(pc[57]), .a(ps[58]),
     .cout(c1[26]), .sum(s1[26]));
mul_csa32  sc1_25_ ( .c(a1s[9]), .b(pc[56]), .a(ps[57]),
     .cout(c1[25]), .sum(s1[25]));
mul_csa32  sc1_24_ ( .c(a1s[8]), .b(pc[55]), .a(ps[56]),
     .cout(c1[24]), .sum(s1[24]));
mul_csa32  sc1_23_ ( .c(a1s[7]), .b(pc[54]), .a(ps[55]),
     .cout(c1[23]), .sum(s1[23]));
mul_csa32  sc1_22_ ( .c(a1s[6]), .b(pc[53]), .a(ps[54]),
     .cout(c1[22]), .sum(s1[22]));
mul_csa32  sc1_21_ ( .c(a1s[5]), .b(pc[52]), .a(ps[53]),
     .cout(c1[21]), .sum(s1[21]));
mul_csa32  sc1_20_ ( .c(a1s[4]), .b(pc[51]), .a(ps[52]),
     .cout(c1[20]), .sum(s1[20]));
mul_csa32  sc2_81_ ( .c(a0c[80]), .b(c1[80]), .a(s1[81]),
     .cout(c2[81]), .sum(s2[81]));
mul_csa32  sc2_80_ ( .c(a0c[79]), .b(c1[79]), .a(s1[80]),
     .cout(c2[80]), .sum(s2[80]));
mul_csa32  sc2_79_ ( .c(a0c[78]), .b(c1[78]), .a(s1[79]),
     .cout(c2[79]), .sum(s2[79]));
mul_csa32  sc2_78_ ( .c(a0c[77]), .b(c1[77]), .a(s1[78]),
     .cout(c2[78]), .sum(s2[78]));
mul_csa32  sc2_77_ ( .c(a0c[76]), .b(c1[76]), .a(s1[77]),
     .cout(c2[77]), .sum(s2[77]));
mul_csa32  sc2_76_ ( .c(a0c[75]), .b(c1[75]), .a(s1[76]),
     .cout(c2[76]), .sum(s2[76]));
mul_csa32  sc2_75_ ( .c(a0c[74]), .b(c1[74]), .a(s1[75]),
     .cout(c2[75]), .sum(s2[75]));
mul_csa32  sc2_74_ ( .c(a0c[73]), .b(c1[73]), .a(s1[74]),
     .cout(c2[74]), .sum(s2[74]));
mul_csa32  sc2_73_ ( .c(a0c[72]), .b(c1[72]), .a(s1[73]),
     .cout(c2[73]), .sum(s2[73]));
mul_csa32  sc2_72_ ( .c(a0c[71]), .b(c1[71]), .a(s1[72]),
     .cout(c2[72]), .sum(s2[72]));
mul_csa32  sc2_71_ ( .c(a0c[70]), .b(c1[70]), .a(s1[71]),
     .cout(c2[71]), .sum(s2[71]));
mul_csa32  sc2_70_ ( .c(a0c[69]), .b(c1[69]), .a(s1[70]),
     .cout(c2[70]), .sum(s2[70]));
mul_csa32  sc2_69_ ( .c(a0c[68]), .b(c1[68]), .a(s1[69]),
     .cout(c2[69]), .sum(s2[69]));
mul_csa32  sc2_68_ ( .c(a0c[67]), .b(c1[67]), .a(s1[68]),
     .cout(c2[68]), .sum(s2[68]));
mul_csa32  acc_19_ ( .c(c3[18]), .b(s3[19]), .a(ain[19]),
     .cout(pcout[19]), .sum(psum[19]));
mul_csa32  acc_18_ ( .c(c3[17]), .b(s3[18]), .a(ain[18]),
     .cout(pcout[18]), .sum(psum[18]));
mul_csa32  acc_17_ ( .c(c3[16]), .b(s3[17]), .a(ain[17]),
     .cout(pcout[17]), .sum(psum[17]));
mul_csa32  acc_16_ ( .c(c3[15]), .b(s3[16]), .a(ain[16]),
     .cout(pcout[16]), .sum(psum[16]));
mul_csa32  acc_15_ ( .c(1'b0), .b(s3[15]), .a(ain[15]),
     .cout(pcout[15]), .sum(psum[15]));
mul_csa32  sc1_0_ ( .c(a0s[0]), .sum(s1[0]), .cout(c1[0]),
     .a(ps[32]), .b(pc[31]));
mul_csa32  sc1_67_ ( .c(a1c[50]), .b(pc[98]), .a(a1s[51]),
     .cout(c1[67]), .sum(s1[67]));
mul_ha acc_0_ ( .sum(psum[0]), .cout(pcout[0]), .a(ain[0]),
     .b(s2[0]));
mul_ha sc3_98_ ( .sum(psum[98]), .cout(pcout[98]), .a(bot),
     .b(a1c[81]));
mul_ha sc2_96_ ( .b(a1c[79]), .a(a1s[80]), .cout(c2[96]),
     .sum(s2[96]));
mul_ha sc2_95_ ( .b(a1c[78]), .a(a1s[79]), .cout(c2[95]),
     .sum(s2[95]));
mul_ha sc2_94_ ( .b(a1c[77]), .a(a1s[78]), .cout(c2[94]),
     .sum(s2[94]));
mul_ha sc2_93_ ( .b(a1c[76]), .a(a1s[77]), .cout(c2[93]),
     .sum(s2[93]));
mul_ha sc2_92_ ( .b(a1c[75]), .a(a1s[76]), .cout(c2[92]),
     .sum(s2[92]));
mul_ha sc2_91_ ( .b(a1c[74]), .a(a1s[75]), .cout(c2[91]),
     .sum(s2[91]));
mul_ha sc2_90_ ( .b(a1c[73]), .a(a1s[74]), .cout(c2[90]),
     .sum(s2[90]));
mul_ha sc2_89_ ( .b(a1c[72]), .a(a1s[73]), .cout(c2[89]),
     .sum(s2[89]));
mul_ha sc2_88_ ( .b(a1c[71]), .a(a1s[72]), .cout(c2[88]),
     .sum(s2[88]));
mul_ha sc2_87_ ( .b(a1c[70]), .a(a1s[71]), .cout(c2[87]),
     .sum(s2[87]));
mul_ha sc2_86_ ( .b(a1c[69]), .a(a1s[70]), .cout(c2[86]),
     .sum(s2[86]));
mul_ha sc2_85_ ( .b(a1c[68]), .a(a1s[69]), .cout(c2[85]),
     .sum(s2[85]));
mul_ha sc2_84_ ( .b(a1c[67]), .a(a1s[68]), .cout(c2[84]),
     .sum(s2[84]));
mul_ha sc3_81_ ( .b(c2[80]), .a(s2[81]), .cout(c3[81]),
     .sum(s3[81]));
mul_ha sc3_80_ ( .b(c2[79]), .a(s2[80]), .cout(c3[80]),
     .sum(s3[80]));
mul_ha sc3_79_ ( .b(c2[78]), .a(s2[79]), .cout(c3[79]),
     .sum(s3[79]));
mul_ha sc3_78_ ( .b(c2[77]), .a(s2[78]), .cout(c3[78]),
     .sum(s3[78]));
mul_ha sc3_77_ ( .b(c2[76]), .a(s2[77]), .cout(c3[77]),
     .sum(s3[77]));
mul_ha sc3_76_ ( .b(c2[75]), .a(s2[76]), .cout(c3[76]),
     .sum(s3[76]));
mul_ha sc3_75_ ( .b(c2[74]), .a(s2[75]), .cout(c3[75]),
     .sum(s3[75]));
mul_ha sc3_74_ ( .b(c2[73]), .a(s2[74]), .cout(c3[74]),
     .sum(s3[74]));
mul_ha sc3_73_ ( .b(c2[72]), .a(s2[73]), .cout(c3[73]),
     .sum(s3[73]));
mul_ha sc3_72_ ( .b(c2[71]), .a(s2[72]), .cout(c3[72]),
     .sum(s3[72]));
mul_ha sc3_71_ ( .b(c2[70]), .a(s2[71]), .cout(c3[71]),
     .sum(s3[71]));
mul_ha sc3_70_ ( .b(c2[69]), .a(s2[70]), .cout(c3[70]),
     .sum(s3[70]));
mul_ha sc3_69_ ( .b(c2[68]), .a(s2[69]), .cout(c3[69]),
     .sum(s3[69]));
mul_ha accx2 ( .sum(psumx2), .cout(pcoutx2), .a(ainx2), .b(s1x2));
mul_ha sc2_4_ ( .sum(s2[4]), .cout(c2[4]), .a(s1[4]), .b(c1[3]));
mul_ha sc2_3_ ( .sum(s2[3]), .cout(c2[3]), .a(s1[3]), .b(c1[2]));
mul_ha sc2_2_ ( .sum(s2[2]), .cout(c2[2]), .a(s1[2]), .b(c1[1]));
mul_ha sc2_1_ ( .sum(s2[1]), .cout(c2[1]), .a(s1[1]), .b(c1[0]));
mul_ha sc2_0_ ( .sum(s2[0]), .cout(c2[0]), .a(s1[0]), .b(c1x2));
mul_ha sc1x2 ( .sum(s1x2), .cout(c1x2), .a(ps[31]), .b(pc[30]));
endmodule 
module mul_csa32 (sum, cout, a, b, c);
output sum, cout;
input a, b, c;
wire x, y0, y1, y2;
assign x = a ^ b;
assign sum = c ^ x;
assign y0 = a & b ;
assign y1 = a & c ;
assign y2 = b & c ;
assign cout = y0 | y1 | y2 ;
endmodule 
module mul_csa42 (sum, carry, cout, a, b, c, d, cin);
output sum, carry, cout;
input a, b, c, d, cin;
wire x, y, z;
assign x = a ^ b;
assign y = c ^ d;
assign z = x ^ y;
assign sum = z ^ cin ;
assign carry = (b & ~z) | (cin & z);
assign cout = (d & ~y) | (a & y);
endmodule 
module mul_ha ( cout, sum, a, b );
output  cout, sum;
input  a, b;
assign sum = a ^ b;
assign cout = a & b ;
endmodule 
module mul_negen ( n0, n1, b );
output  n0, n1;
input [2:0]  b;
assign n0 = b[2] & b[1] & ~b[0] ;
assign n1 = b[2] & b[1] & b[0] ;
endmodule 
module mul_ppgen3lsb4 (cout, p0_l, p1_l, sum, a, b0, b1 );
output  p0_l, p1_l;
output [3:0]  sum;
output [3:1]  cout;
input [3:0]  a;
input [2:0]  b0;
input [2:0]  b1;
wire b0n, b0n_0, b0n_1, b1n_0, b1n_1;
wire p0_0, p0_1, p0_2, p0_3, p1_2, p1_3;
wire p0_l_0, p0_l_1, p0_l_2, p1_l_2;
assign b0n = b0n_1 | (b0n_0 & p0_0) ;
assign sum[0] = b0n_0 ^ p0_0 ;
mul_negen p0n ( .b(b0[2:0]), .n1(b0n_1), .n0(b0n_0));
mul_negen p1n ( .b(b1[2:0]), .n1(b1n_1), .n0(b1n_0));
mul_csa32  sc1_2_ ( .c(b1n_0), .sum(sum[2]), .cout(cout[2]),
     .a(p0_2), .b(p1_2));
mul_csa32  sc1_3_ ( .c(b1n_1), .sum(sum[3]), .cout(cout[3]),
     .a(p0_3), .b(p1_3));
mul_ha sc1_1_ ( .sum(sum[1]), .cout(cout[1]), .a(p0_1),
     .b(b0n));
mul_ppgen p0_3_ ( .pm1_l(p0_l_2), .p_l(p0_l), .b(b0[2:0]), .a(a[3]),
     .z(p0_3));
mul_ppgen p1_3_ ( .pm1_l(p1_l_2), .p_l(p1_l), .b(b1[2:0]), .a(a[1]),
     .z(p1_3));
mul_ppgen p0_2_ ( .pm1_l(p0_l_1), .p_l(p0_l_2), .b(b0[2:0]),
     .a(a[2]), .z(p0_2));
mul_ppgen p0_1_ ( .pm1_l(p0_l_0), .p_l(p0_l_1), .b(b0[2:0]),
     .a(a[1]), .z(p0_1));
mul_ppgen p0_0_ ( .pm1_l(1'b1), .p_l(p0_l_0),
     .b(b0[2:0]), .a(a[0]), .z(p0_0));
mul_ppgen p1_2_ ( .pm1_l(1'b1), .p_l(p1_l_2),
     .b(b1[2:0]), .a(a[0]), .z(p1_2));
endmodule 
module mul_ppgen3sign ( cout, sum, am1, am2, am3, am4, b0, b1, b2,
     bot, head, p0m1_l, p1m1_l, p2m1_l );
input  am1, am2, am3, am4;
input  bot, head, p0m1_l, p1m1_l, p2m1_l;
output [5:0]  sum;
output [4:0]  cout;
input [2:0]  b0;
input [2:0]  b2;
input [2:0]  b1;
wire net37, net42, net075, net088, net0117; 
wire net47, net073, net38, net0118, net078, net8, net15, net43, net48, net35;
wire p2_l_67, p2_l_66, p2_l_65, p2_l_64; 
wire p1_l_65, p1_l_64; 
assign sum[5] = bot & net075 ;
assign net0117 = head & net088 ; 
assign net37 = ~net0117 ;
assign net42 = head ^ net088 ;
mul_ppgensign p0_64_ ( .b(b0[2:0]), .z(net47), .p_l(net088),
     .pm1_l(p0m1_l));
mul_ppgensign p2_68_ ( .pm1_l(p2_l_67), .b(b2[2:0]), .z(net073),
     .p_l(net075));
mul_ppgensign p1_66_ ( .pm1_l(p1_l_65), .b(b1[2:0]), .z(net38),
     .p_l(net0118));
mul_ha sc1_68_ ( .b(net073), .a(1'b1), .cout(cout[4]),
     .sum(sum[4]));
mul_ppgen p2_67_ ( .pm1_l(p2_l_66), .b(b2[2:0]), .a(am1), .z(net078),
     .p_l(p2_l_67));
mul_ppgen p2_66_ ( .pm1_l(p2_l_65), .b(b2[2:0]), .a(am2), .z(net8),
     .p_l(p2_l_66));
mul_ppgen p2_65_ ( .pm1_l(p2_l_64), .p_l(p2_l_65), .b(b2[2:0]),
     .a(am3), .z(net15));
mul_ppgen p1_65_ ( .pm1_l(p1_l_64), .p_l(p1_l_65), .b(b1[2:0]),
     .a(am1), .z(net43));
mul_ppgen p1_64_ ( .pm1_l(p1m1_l), .p_l(p1_l_64), .b(b1[2:0]),
     .a(am2), .z(net48));
mul_ppgen p2_64_ ( .pm1_l(p2m1_l), .p_l(p2_l_64), .b(b2[2:0]),
     .a(am4), .z(net35));
mul_csa32  sc1_67_ ( .c(net078), .b(net0117), .a(net0118),
     .cout(cout[3]), .sum(sum[3]));
mul_csa32  sc1_66_ ( .c(net8), .b(net37), .a(net38), .cout(cout[2]),
     .sum(sum[2]));
mul_csa32  sc1_65_ ( .c(net15), .b(net42), .a(net43), .cout(cout[1]),
     .sum(sum[1]));
mul_csa32  sc1_64_ ( .c(net35), .b(net47), .a(net48), .cout(cout[0]),
     .sum(sum[0]));
endmodule 
module mul_ppgen3 ( cout, p0_l, p1_l, p2_l, sum, am2, am4,
     a, b0, b1, b2, p0m1_l, p1m1_l, p2m1_l );
output  cout, p0_l, p1_l, p2_l, sum;
input  am2, am4;
input  a, p0m1_l, p1m1_l, p2m1_l;
input [2:0]  b0;
input [2:0]  b2;
input [2:0]  b1;
wire net046, net32, net043;
mul_csa32  sc1 ( .a(net046), .b(net32), .cout(cout), .sum(sum),
     .c(net043));
mul_ppgen p2 ( .pm1_l(p2m1_l), .p_l(p2_l), .b(b2[2:0]), .a(am4),
     .z(net043));
mul_ppgen p1 ( .pm1_l(p1m1_l), .p_l(p1_l), .b(b1[2:0]), .a(am2),
     .z(net046));
mul_ppgen p0 ( .pm1_l(p0m1_l), .p_l(p0_l), .b(b0[2:0]), .a(a),
     .z(net32));
endmodule 
module mul_ppgenrow3 ( cout, sum, a, b0, b1, b2, bot, head );
output [68:1]  cout;
output [69:0]  sum;
input [63:0]  a;
input [2:0]  b2;
input [2:0]  b0;
input [2:0]  b1;
input  bot, head;
wire  [63:4]  p2_l;
wire  [63:3]  p1_l;
wire  [63:3]  p0_l;
mul_ppgen3sign I2 ( .am4(a[60]), .am3(a[61]), .am2(a[62]),
     .am1(a[63]), .p2m1_l(p2_l[63]), .p1m1_l(p1_l[63]),
     .p0m1_l(p0_l[63]), .b2(b2[2:0]), .head(head), .bot(bot),
     .sum(sum[69:64]), .cout(cout[68:64]), .b1(b1[2:0]), .b0(b0[2:0]));
mul_ppgen3 I1_63_ ( .p2_l(p2_l[63]), .b2(b2[2:0]),
     .am2(a[61]), .a(a[63]), .p2m1_l(p2_l[62]),
     .p1m1_l(p1_l[62]), .p0m1_l(p0_l[62]), .am4(a[59]), .sum(sum[63]),
     .cout(cout[63]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[63]),
     .p0_l(p0_l[63]));
mul_ppgen3 I1_62_ ( .p2_l(p2_l[62]), .b2(b2[2:0]), 
     .am2(a[60]), .a(a[62]), .p2m1_l(p2_l[61]),
     .p1m1_l(p1_l[61]), .p0m1_l(p0_l[61]), .am4(a[58]), .sum(sum[62]),
     .cout(cout[62]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[62]),
     .p0_l(p0_l[62]));
mul_ppgen3 I1_61_ ( .p2_l(p2_l[61]), .b2(b2[2:0]), 
     .am2(a[59]), .a(a[61]), .p2m1_l(p2_l[60]),
     .p1m1_l(p1_l[60]), .p0m1_l(p0_l[60]), .am4(a[57]), .sum(sum[61]),
     .cout(cout[61]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[61]),
     .p0_l(p0_l[61]));
mul_ppgen3 I1_60_ ( .p2_l(p2_l[60]), .b2(b2[2:0]), 
     .am2(a[58]), .a(a[60]), .p2m1_l(p2_l[59]),
     .p1m1_l(p1_l[59]), .p0m1_l(p0_l[59]), .am4(a[56]), .sum(sum[60]),
     .cout(cout[60]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[60]),
     .p0_l(p0_l[60]));
mul_ppgen3 I1_59_ ( .p2_l(p2_l[59]), .b2(b2[2:0]), 
     .am2(a[57]), .a(a[59]), .p2m1_l(p2_l[58]),
     .p1m1_l(p1_l[58]), .p0m1_l(p0_l[58]), .am4(a[55]), .sum(sum[59]),
     .cout(cout[59]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[59]),
     .p0_l(p0_l[59]));
mul_ppgen3 I1_58_ ( .p2_l(p2_l[58]), .b2(b2[2:0]), 
     .am2(a[56]), .a(a[58]), .p2m1_l(p2_l[57]),
     .p1m1_l(p1_l[57]), .p0m1_l(p0_l[57]), .am4(a[54]), .sum(sum[58]),
     .cout(cout[58]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[58]),
     .p0_l(p0_l[58]));
mul_ppgen3 I1_57_ ( .p2_l(p2_l[57]), .b2(b2[2:0]), 
     .am2(a[55]), .a(a[57]), .p2m1_l(p2_l[56]),
     .p1m1_l(p1_l[56]), .p0m1_l(p0_l[56]), .am4(a[53]), .sum(sum[57]),
     .cout(cout[57]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[57]),
     .p0_l(p0_l[57]));
mul_ppgen3 I1_56_ ( .p2_l(p2_l[56]), .b2(b2[2:0]), 
     .am2(a[54]), .a(a[56]), .p2m1_l(p2_l[55]),
     .p1m1_l(p1_l[55]), .p0m1_l(p0_l[55]), .am4(a[52]), .sum(sum[56]),
     .cout(cout[56]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[56]),
     .p0_l(p0_l[56]));
mul_ppgen3 I1_55_ ( .p2_l(p2_l[55]), .b2(b2[2:0]), 
     .am2(a[53]), .a(a[55]), .p2m1_l(p2_l[54]),
     .p1m1_l(p1_l[54]), .p0m1_l(p0_l[54]), .am4(a[51]), .sum(sum[55]),
     .cout(cout[55]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[55]),
     .p0_l(p0_l[55]));
mul_ppgen3 I1_54_ ( .p2_l(p2_l[54]), .b2(b2[2:0]), 
     .am2(a[52]), .a(a[54]), .p2m1_l(p2_l[53]),
     .p1m1_l(p1_l[53]), .p0m1_l(p0_l[53]), .am4(a[50]), .sum(sum[54]),
     .cout(cout[54]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[54]),
     .p0_l(p0_l[54]));
mul_ppgen3 I1_53_ ( .p2_l(p2_l[53]), .b2(b2[2:0]), 
     .am2(a[51]), .a(a[53]), .p2m1_l(p2_l[52]),
     .p1m1_l(p1_l[52]), .p0m1_l(p0_l[52]), .am4(a[49]), .sum(sum[53]),
     .cout(cout[53]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[53]),
     .p0_l(p0_l[53]));
mul_ppgen3 I1_52_ ( .p2_l(p2_l[52]), .b2(b2[2:0]), 
     .am2(a[50]), .a(a[52]), .p2m1_l(p2_l[51]),
     .p1m1_l(p1_l[51]), .p0m1_l(p0_l[51]), .am4(a[48]), .sum(sum[52]),
     .cout(cout[52]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[52]),
     .p0_l(p0_l[52]));
mul_ppgen3 I1_51_ ( .p2_l(p2_l[51]), .b2(b2[2:0]), 
     .am2(a[49]), .a(a[51]), .p2m1_l(p2_l[50]),
     .p1m1_l(p1_l[50]), .p0m1_l(p0_l[50]), .am4(a[47]), .sum(sum[51]),
     .cout(cout[51]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[51]),
     .p0_l(p0_l[51]));
mul_ppgen3 I1_50_ ( .p2_l(p2_l[50]), .b2(b2[2:0]), 
     .am2(a[48]), .a(a[50]), .p2m1_l(p2_l[49]),
     .p1m1_l(p1_l[49]), .p0m1_l(p0_l[49]), .am4(a[46]), .sum(sum[50]),
     .cout(cout[50]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[50]),
     .p0_l(p0_l[50]));
mul_ppgen3 I1_49_ ( .p2_l(p2_l[49]), .b2(b2[2:0]), 
     .am2(a[47]), .a(a[49]), .p2m1_l(p2_l[48]),
     .p1m1_l(p1_l[48]), .p0m1_l(p0_l[48]), .am4(a[45]), .sum(sum[49]),
     .cout(cout[49]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[49]),
     .p0_l(p0_l[49]));
mul_ppgen3 I1_48_ ( .p2_l(p2_l[48]), .b2(b2[2:0]), 
     .am2(a[46]), .a(a[48]), .p2m1_l(p2_l[47]),
     .p1m1_l(p1_l[47]), .p0m1_l(p0_l[47]), .am4(a[44]), .sum(sum[48]),
     .cout(cout[48]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[48]),
     .p0_l(p0_l[48]));
mul_ppgen3 I1_47_ ( .p2_l(p2_l[47]), .b2(b2[2:0]), 
     .am2(a[45]), .a(a[47]), .p2m1_l(p2_l[46]),
     .p1m1_l(p1_l[46]), .p0m1_l(p0_l[46]), .am4(a[43]), .sum(sum[47]),
     .cout(cout[47]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[47]),
     .p0_l(p0_l[47]));
mul_ppgen3 I1_46_ ( .p2_l(p2_l[46]), .b2(b2[2:0]), 
     .am2(a[44]), .a(a[46]), .p2m1_l(p2_l[45]),
     .p1m1_l(p1_l[45]), .p0m1_l(p0_l[45]), .am4(a[42]), .sum(sum[46]),
     .cout(cout[46]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[46]),
     .p0_l(p0_l[46]));
mul_ppgen3 I1_45_ ( .p2_l(p2_l[45]), .b2(b2[2:0]), 
     .am2(a[43]), .a(a[45]), .p2m1_l(p2_l[44]),
     .p1m1_l(p1_l[44]), .p0m1_l(p0_l[44]), .am4(a[41]), .sum(sum[45]),
     .cout(cout[45]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[45]),
     .p0_l(p0_l[45]));
mul_ppgen3 I1_44_ ( .p2_l(p2_l[44]), .b2(b2[2:0]), 
     .am2(a[42]), .a(a[44]), .p2m1_l(p2_l[43]),
     .p1m1_l(p1_l[43]), .p0m1_l(p0_l[43]), .am4(a[40]), .sum(sum[44]),
     .cout(cout[44]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[44]),
     .p0_l(p0_l[44]));
mul_ppgen3 I1_43_ ( .p2_l(p2_l[43]), .b2(b2[2:0]), 
     .am2(a[41]), .a(a[43]), .p2m1_l(p2_l[42]),
     .p1m1_l(p1_l[42]), .p0m1_l(p0_l[42]), .am4(a[39]), .sum(sum[43]),
     .cout(cout[43]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[43]),
     .p0_l(p0_l[43]));
mul_ppgen3 I1_42_ ( .p2_l(p2_l[42]), .b2(b2[2:0]), 
     .am2(a[40]), .a(a[42]), .p2m1_l(p2_l[41]),
     .p1m1_l(p1_l[41]), .p0m1_l(p0_l[41]), .am4(a[38]), .sum(sum[42]),
     .cout(cout[42]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[42]),
     .p0_l(p0_l[42]));
mul_ppgen3 I1_41_ ( .p2_l(p2_l[41]), .b2(b2[2:0]), 
     .am2(a[39]), .a(a[41]), .p2m1_l(p2_l[40]),
     .p1m1_l(p1_l[40]), .p0m1_l(p0_l[40]), .am4(a[37]), .sum(sum[41]),
     .cout(cout[41]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[41]),
     .p0_l(p0_l[41]));
mul_ppgen3 I1_40_ ( .p2_l(p2_l[40]), .b2(b2[2:0]), 
     .am2(a[38]), .a(a[40]), .p2m1_l(p2_l[39]),
     .p1m1_l(p1_l[39]), .p0m1_l(p0_l[39]), .am4(a[36]), .sum(sum[40]),
     .cout(cout[40]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[40]),
     .p0_l(p0_l[40]));
mul_ppgen3 I1_39_ ( .p2_l(p2_l[39]), .b2(b2[2:0]), 
     .am2(a[37]), .a(a[39]), .p2m1_l(p2_l[38]),
     .p1m1_l(p1_l[38]), .p0m1_l(p0_l[38]), .am4(a[35]), .sum(sum[39]),
     .cout(cout[39]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[39]),
     .p0_l(p0_l[39]));
mul_ppgen3 I1_38_ ( .p2_l(p2_l[38]), .b2(b2[2:0]), 
     .am2(a[36]), .a(a[38]), .p2m1_l(p2_l[37]),
     .p1m1_l(p1_l[37]), .p0m1_l(p0_l[37]), .am4(a[34]), .sum(sum[38]),
     .cout(cout[38]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[38]),
     .p0_l(p0_l[38]));
mul_ppgen3 I1_37_ ( .p2_l(p2_l[37]), .b2(b2[2:0]), 
     .am2(a[35]), .a(a[37]), .p2m1_l(p2_l[36]),
     .p1m1_l(p1_l[36]), .p0m1_l(p0_l[36]), .am4(a[33]), .sum(sum[37]),
     .cout(cout[37]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[37]),
     .p0_l(p0_l[37]));
mul_ppgen3 I1_36_ ( .p2_l(p2_l[36]), .b2(b2[2:0]), 
     .am2(a[34]), .a(a[36]), .p2m1_l(p2_l[35]),
     .p1m1_l(p1_l[35]), .p0m1_l(p0_l[35]), .am4(a[32]), .sum(sum[36]),
     .cout(cout[36]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[36]),
     .p0_l(p0_l[36]));
mul_ppgen3 I1_35_ ( .p2_l(p2_l[35]), .b2(b2[2:0]), 
     .am2(a[33]), .a(a[35]), .p2m1_l(p2_l[34]),
     .p1m1_l(p1_l[34]), .p0m1_l(p0_l[34]), .am4(a[31]), .sum(sum[35]),
     .cout(cout[35]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[35]),
     .p0_l(p0_l[35]));
mul_ppgen3 I1_34_ ( .p2_l(p2_l[34]), .b2(b2[2:0]), 
     .am2(a[32]), .a(a[34]), .p2m1_l(p2_l[33]),
     .p1m1_l(p1_l[33]), .p0m1_l(p0_l[33]), .am4(a[30]), .sum(sum[34]),
     .cout(cout[34]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[34]),
     .p0_l(p0_l[34]));
mul_ppgen3 I1_33_ ( .p2_l(p2_l[33]), .b2(b2[2:0]), 
     .am2(a[31]), .a(a[33]), .p2m1_l(p2_l[32]),
     .p1m1_l(p1_l[32]), .p0m1_l(p0_l[32]), .am4(a[29]), .sum(sum[33]),
     .cout(cout[33]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[33]),
     .p0_l(p0_l[33]));
mul_ppgen3 I1_32_ ( .p2_l(p2_l[32]), .b2(b2[2:0]), 
     .am2(a[30]), .a(a[32]), .p2m1_l(p2_l[31]),
     .p1m1_l(p1_l[31]), .p0m1_l(p0_l[31]), .am4(a[28]), .sum(sum[32]),
     .cout(cout[32]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[32]),
     .p0_l(p0_l[32]));
mul_ppgen3 I1_31_ ( .p2_l(p2_l[31]), .b2(b2[2:0]), 
     .am2(a[29]), .a(a[31]), .p2m1_l(p2_l[30]),
     .p1m1_l(p1_l[30]), .p0m1_l(p0_l[30]), .am4(a[27]), .sum(sum[31]),
     .cout(cout[31]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[31]),
     .p0_l(p0_l[31]));
mul_ppgen3 I1_30_ ( .p2_l(p2_l[30]), .b2(b2[2:0]), 
     .am2(a[28]), .a(a[30]), .p2m1_l(p2_l[29]),
     .p1m1_l(p1_l[29]), .p0m1_l(p0_l[29]), .am4(a[26]), .sum(sum[30]),
     .cout(cout[30]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[30]),
     .p0_l(p0_l[30]));
mul_ppgen3 I1_29_ ( .p2_l(p2_l[29]), .b2(b2[2:0]), 
     .am2(a[27]), .a(a[29]), .p2m1_l(p2_l[28]),
     .p1m1_l(p1_l[28]), .p0m1_l(p0_l[28]), .am4(a[25]), .sum(sum[29]),
     .cout(cout[29]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[29]),
     .p0_l(p0_l[29]));
mul_ppgen3 I1_28_ ( .p2_l(p2_l[28]), .b2(b2[2:0]), 
     .am2(a[26]), .a(a[28]), .p2m1_l(p2_l[27]),
     .p1m1_l(p1_l[27]), .p0m1_l(p0_l[27]), .am4(a[24]), .sum(sum[28]),
     .cout(cout[28]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[28]),
     .p0_l(p0_l[28]));
mul_ppgen3 I1_27_ ( .p2_l(p2_l[27]), .b2(b2[2:0]), 
     .am2(a[25]), .a(a[27]), .p2m1_l(p2_l[26]),
     .p1m1_l(p1_l[26]), .p0m1_l(p0_l[26]), .am4(a[23]), .sum(sum[27]),
     .cout(cout[27]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[27]),
     .p0_l(p0_l[27]));
mul_ppgen3 I1_26_ ( .p2_l(p2_l[26]), .b2(b2[2:0]), 
     .am2(a[24]), .a(a[26]), .p2m1_l(p2_l[25]),
     .p1m1_l(p1_l[25]), .p0m1_l(p0_l[25]), .am4(a[22]), .sum(sum[26]),
     .cout(cout[26]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[26]),
     .p0_l(p0_l[26]));
mul_ppgen3 I1_25_ ( .p2_l(p2_l[25]), .b2(b2[2:0]), 
     .am2(a[23]), .a(a[25]), .p2m1_l(p2_l[24]),
     .p1m1_l(p1_l[24]), .p0m1_l(p0_l[24]), .am4(a[21]), .sum(sum[25]),
     .cout(cout[25]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[25]),
     .p0_l(p0_l[25]));
mul_ppgen3 I1_24_ ( .p2_l(p2_l[24]), .b2(b2[2:0]), 
     .am2(a[22]), .a(a[24]), .p2m1_l(p2_l[23]),
     .p1m1_l(p1_l[23]), .p0m1_l(p0_l[23]), .am4(a[20]), .sum(sum[24]),
     .cout(cout[24]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[24]),
     .p0_l(p0_l[24]));
mul_ppgen3 I1_23_ ( .p2_l(p2_l[23]), .b2(b2[2:0]), 
     .am2(a[21]), .a(a[23]), .p2m1_l(p2_l[22]),
     .p1m1_l(p1_l[22]), .p0m1_l(p0_l[22]), .am4(a[19]), .sum(sum[23]),
     .cout(cout[23]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[23]),
     .p0_l(p0_l[23]));
mul_ppgen3 I1_22_ ( .p2_l(p2_l[22]), .b2(b2[2:0]), 
     .am2(a[20]), .a(a[22]), .p2m1_l(p2_l[21]),
     .p1m1_l(p1_l[21]), .p0m1_l(p0_l[21]), .am4(a[18]), .sum(sum[22]),
     .cout(cout[22]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[22]),
     .p0_l(p0_l[22]));
mul_ppgen3 I1_21_ ( .p2_l(p2_l[21]), .b2(b2[2:0]), 
     .am2(a[19]), .a(a[21]), .p2m1_l(p2_l[20]),
     .p1m1_l(p1_l[20]), .p0m1_l(p0_l[20]), .am4(a[17]), .sum(sum[21]),
     .cout(cout[21]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[21]),
     .p0_l(p0_l[21]));
mul_ppgen3 I1_20_ ( .p2_l(p2_l[20]), .b2(b2[2:0]), 
     .am2(a[18]), .a(a[20]), .p2m1_l(p2_l[19]),
     .p1m1_l(p1_l[19]), .p0m1_l(p0_l[19]), .am4(a[16]), .sum(sum[20]),
     .cout(cout[20]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[20]),
     .p0_l(p0_l[20]));
mul_ppgen3 I1_19_ ( .p2_l(p2_l[19]), .b2(b2[2:0]), 
     .am2(a[17]), .a(a[19]), .p2m1_l(p2_l[18]),
     .p1m1_l(p1_l[18]), .p0m1_l(p0_l[18]), .am4(a[15]), .sum(sum[19]),
     .cout(cout[19]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[19]),
     .p0_l(p0_l[19]));
mul_ppgen3 I1_18_ ( .p2_l(p2_l[18]), .b2(b2[2:0]), 
     .am2(a[16]), .a(a[18]), .p2m1_l(p2_l[17]),
     .p1m1_l(p1_l[17]), .p0m1_l(p0_l[17]), .am4(a[14]), .sum(sum[18]),
     .cout(cout[18]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[18]),
     .p0_l(p0_l[18]));
mul_ppgen3 I1_17_ ( .p2_l(p2_l[17]), .b2(b2[2:0]), 
     .am2(a[15]), .a(a[17]), .p2m1_l(p2_l[16]),
     .p1m1_l(p1_l[16]), .p0m1_l(p0_l[16]), .am4(a[13]), .sum(sum[17]),
     .cout(cout[17]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[17]),
     .p0_l(p0_l[17]));
mul_ppgen3 I1_16_ ( .p2_l(p2_l[16]), .b2(b2[2:0]), 
     .am2(a[14]), .a(a[16]), .p2m1_l(p2_l[15]),
     .p1m1_l(p1_l[15]), .p0m1_l(p0_l[15]), .am4(a[12]), .sum(sum[16]),
     .cout(cout[16]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[16]),
     .p0_l(p0_l[16]));
mul_ppgen3 I1_15_ ( .p2_l(p2_l[15]), .b2(b2[2:0]), 
     .am2(a[13]), .a(a[15]), .p2m1_l(p2_l[14]),
     .p1m1_l(p1_l[14]), .p0m1_l(p0_l[14]), .am4(a[11]), .sum(sum[15]),
     .cout(cout[15]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[15]),
     .p0_l(p0_l[15]));
mul_ppgen3 I1_14_ ( .p2_l(p2_l[14]), .b2(b2[2:0]), 
     .am2(a[12]), .a(a[14]), .p2m1_l(p2_l[13]),
     .p1m1_l(p1_l[13]), .p0m1_l(p0_l[13]), .am4(a[10]), .sum(sum[14]),
     .cout(cout[14]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[14]),
     .p0_l(p0_l[14]));
mul_ppgen3 I1_13_ ( .p2_l(p2_l[13]), .b2(b2[2:0]), 
     .am2(a[11]), .a(a[13]), .p2m1_l(p2_l[12]),
     .p1m1_l(p1_l[12]), .p0m1_l(p0_l[12]), .am4(a[9]), .sum(sum[13]),
     .cout(cout[13]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[13]),
     .p0_l(p0_l[13]));
mul_ppgen3 I1_12_ ( .p2_l(p2_l[12]), .b2(b2[2:0]), 
     .am2(a[10]), .a(a[12]), .p2m1_l(p2_l[11]),
     .p1m1_l(p1_l[11]), .p0m1_l(p0_l[11]), .am4(a[8]), .sum(sum[12]),
     .cout(cout[12]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[12]),
     .p0_l(p0_l[12]));
mul_ppgen3 I1_11_ ( .p2_l(p2_l[11]), .b2(b2[2:0]), 
     .am2(a[9]), .a(a[11]), .p2m1_l(p2_l[10]),
     .p1m1_l(p1_l[10]), .p0m1_l(p0_l[10]), .am4(a[7]), .sum(sum[11]),
     .cout(cout[11]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[11]),
     .p0_l(p0_l[11]));
mul_ppgen3 I1_10_ ( .p2_l(p2_l[10]), .b2(b2[2:0]), 
     .am2(a[8]), .a(a[10]), .p2m1_l(p2_l[9]),
     .p1m1_l(p1_l[9]), .p0m1_l(p0_l[9]), .am4(a[6]), .sum(sum[10]),
     .cout(cout[10]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[10]),
     .p0_l(p0_l[10]));
mul_ppgen3 I1_9_ ( .p2_l(p2_l[9]), .b2(b2[2:0]), 
     .am2(a[7]), .a(a[9]), .p2m1_l(p2_l[8]),
     .p1m1_l(p1_l[8]), .p0m1_l(p0_l[8]), .am4(a[5]), .sum(sum[9]),
     .cout(cout[9]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[9]),
     .p0_l(p0_l[9]));
mul_ppgen3 I1_8_ ( .p2_l(p2_l[8]), .b2(b2[2:0]), 
     .am2(a[6]), .a(a[8]), .p2m1_l(p2_l[7]),
     .p1m1_l(p1_l[7]), .p0m1_l(p0_l[7]), .am4(a[4]), .sum(sum[8]),
     .cout(cout[8]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[8]),
     .p0_l(p0_l[8]));
mul_ppgen3 I1_7_ ( .p2_l(p2_l[7]), .b2(b2[2:0]), 
     .am2(a[5]), .a(a[7]), .p2m1_l(p2_l[6]),
     .p1m1_l(p1_l[6]), .p0m1_l(p0_l[6]), .am4(a[3]), .sum(sum[7]),
     .cout(cout[7]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[7]),
     .p0_l(p0_l[7]));
mul_ppgen3 I1_6_ ( .p2_l(p2_l[6]), .b2(b2[2:0]), 
     .am2(a[4]), .a(a[6]), .p2m1_l(p2_l[5]),
     .p1m1_l(p1_l[5]), .p0m1_l(p0_l[5]), .am4(a[2]), .sum(sum[6]),
     .cout(cout[6]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[6]),
     .p0_l(p0_l[6]));
mul_ppgen3 I1_5_ ( .p2_l(p2_l[5]), .b2(b2[2:0]), 
     .am2(a[3]), .a(a[5]), .p2m1_l(p2_l[4]),
     .p1m1_l(p1_l[4]), .p0m1_l(p0_l[4]), .am4(a[1]), .sum(sum[5]),
     .cout(cout[5]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[5]),
     .p0_l(p0_l[5]));
mul_ppgen3 I1_4_ ( .p2_l(p2_l[4]), .b2(b2[2:0]), 
     .am2(a[2]), .a(a[4]), .p2m1_l(1'b1),
     .p1m1_l(p1_l[3]), .p0m1_l(p0_l[3]), .am4(a[0]), .sum(sum[4]),
     .cout(cout[4]), .b1(b1[2:0]), .b0(b0[2:0]), .p1_l(p1_l[4]),
     .p0_l(p0_l[4]));
mul_ppgen3lsb4 I0 ( .cout(cout[3:1]), .a(a[3:0]), .sum(sum[3:0]),
     .p1_l(p1_l[3]), .p0_l(p0_l[3]), .b1(b1[2:0]), .b0(b0[2:0]));
endmodule 
module mul_ppgensign ( p_l, z, b, pm1_l );
output  p_l, z;
input  pm1_l;
input [2:0]  b;
assign p_l = ~(b[1] & b[2]);
assign z = b[0] ? ~pm1_l : ~p_l ;
endmodule 
module mul_ppgen ( p_l, z, a, b, pm1_l );
output  p_l, z;
input  a, pm1_l;
input [2:0]  b;
assign p_l = ~((a ^ b[2]) & b[1]) ;
assign z = b[0] ? ~pm1_l : ~p_l ;
endmodule 
module mul_mux2 ( z, d0, d1, s );
output  z;
input  d0, d1, s;
assign z = s ? d1 : d0 ;
endmodule 
module mul_booth(
	head,
        b_in,
        b0, b1, b2, b3, b4, b5, b6, b7,
	b8, b9, b10, b11, b12, b13, b14, b15, b16,
	clk, se, si, so, mul_step, tm_l
	);
input		head;		
input   [63:0] 	b_in;
input		clk, se, si, mul_step, tm_l;
output  [2:0]  	b0, b1, b2, b3, b4, b5, b6, b7, b8, b9, b10, b11, b12, b13, b14, b15;
output 		b16;
output 		so;
wire  [63:31] 	b;
wire [2:0] 	b0_in0, b1_in0,  b2_in0,  b3_in0,  b4_in0,  b5_in0,  b6_in0,  b7_in0 ;
wire [2:0] 	b8_in0, b9_in0, b10_in0, b11_in0, b12_in0, b13_in0, b14_in0, b15_in0 ;
wire [2:0] 	b0_in1, b1_in1,  b2_in1,  b3_in1,  b4_in1,  b5_in1,  b6_in1,  b7_in1 ;
wire [2:0] 	b8_in1, b9_in1, b10_in1, b11_in1, b12_in1, b13_in1, b14_in1, b15_in1 ;
wire 	   	b16_in1;
wire [2:0] 	b0_outmx, b1_outmx, b2_outmx, b3_outmx, b4_outmx, b5_outmx, b6_outmx;
wire [2:0] 	b7_outmx, b8_outmx, b9_outmx, b10_outmx, b11_outmx, b12_outmx, b13_outmx;
wire [2:0] 	b14_outmx, b15_outmx;
wire 	   	b16_outmx;
wire		clk_enb0, clk_enb1;
  mul_bodec 		encode0_a(
				.x  (1'b0),
				.b  (b_in[15:0]),
				.b0 (b0_in0),
				.b1 (b1_in0),
				.b2 (b2_in0),
				.b3 (b3_in0),
				.b4 (b4_in0),
				.b5 (b5_in0),
				.b6 (b6_in0),
				.b7 (b7_in0)
				);
				
				
  mul_bodec		encode0_b(
				.x  (b_in[15]),
				.b  (b_in[31:16]),
				.b0 (b8_in0),
				.b1 (b9_in0),
				.b2 (b10_in0),
				.b3 (b11_in0),
				.b4 (b12_in0),
				.b5 (b13_in0),
				.b6 (b14_in0),
				.b7 (b15_in0)
				);
				
				
  
  clken_buf     ckbuf_0(.clk(clk_enb0), .rclk(clk), .enb_l(~mul_step), .tmb_l(tm_l));
  clken_buf     ckbuf_1(.clk(clk_enb1), .rclk(clk), .enb_l(~(head & mul_step)), .tmb_l(tm_l));
  dff_s 			hld_dff0(.din(b_in[31]), .clk(clk_enb1), .q(b[31]),
                        	.se(se), .si(), .so());
  dff_s #(32) 		hld_dff(.din(b_in[63:32]), .clk(clk_enb1), .q(b[63:32]),
				.se(se), .si(), .so());
  mul_bodec     	encode1_a(
                        	.x  (b[31]),
                        	.b  (b[47:32]),
                        	.b0 (b0_in1),
                        	.b1 (b1_in1),
                        	.b2 (b2_in1),
                        	.b3 (b3_in1),
                        	.b4 (b4_in1),
                        	.b5 (b5_in1),
                        	.b6 (b6_in1),
                        	.b7 (b7_in1)
                        	);
                        	
                        	
  mul_bodec     	encode1_b(
                        	.x  (b[47]),
                        	.b  (b[63:48]),
                        	.b0 (b8_in1),
                        	.b1 (b9_in1),
                        	.b2 (b10_in1),
                        	.b3 (b11_in1),
                        	.b4 (b12_in1),
                        	.b5 (b13_in1),
                        	.b6 (b14_in1),
                        	.b7 (b15_in1)
                        	);
				assign b16_in1 = b[63] ;
  dp_mux2es #(3)    out_mux0(.dout(b0_outmx[2:0]),
                        .in0(b0_in0[2:0]),
                        .in1(b0_in1[2:0]),
                        .sel(~head));
  dp_mux2es #(3)    out_mux1(.dout(b1_outmx[2:0]),
                        .in0(b1_in0[2:0]),
                        .in1(b1_in1[2:0]),
                        .sel(~head));
  dp_mux2es #(3)    out_mux2(.dout(b2_outmx[2:0]),
                        .in0(b2_in0[2:0]),
                        .in1(b2_in1[2:0]),
                        .sel(~head));
  dp_mux2es #(3)    out_mux3(.dout(b3_outmx[2:0]),
                        .in0(b3_in0[2:0]),
                        .in1(b3_in1[2:0]),
                        .sel(~head));
  dp_mux2es #(3)    out_mux4(.dout(b4_outmx[2:0]),
                        .in0(b4_in0[2:0]),
                        .in1(b4_in1[2:0]),
                        .sel(~head));
  dp_mux2es #(3)    out_mux5(.dout(b5_outmx[2:0]),
                        .in0(b5_in0[2:0]),
                        .in1(b5_in1[2:0]),
                        .sel(~head));
  dp_mux2es #(3)    out_mux6(.dout(b6_outmx[2:0]),
                        .in0(b6_in0[2:0]),
                        .in1(b6_in1[2:0]),
                        .sel(~head));
  dp_mux2es #(3)    out_mux7(.dout(b7_outmx[2:0]),
                        .in0(b7_in0[2:0]),
                        .in1(b7_in1[2:0]),
                        .sel(~head));
  dp_mux2es #(3)    out_mux8(.dout(b8_outmx[2:0]),
                        .in0(b8_in0[2:0]),
                        .in1(b8_in1[2:0]),
                        .sel(~head));
  dp_mux2es #(3)    out_mux9(.dout(b9_outmx[2:0]),
                        .in0(b9_in0[2:0]),
                        .in1(b9_in1[2:0]),
                        .sel(~head));
  dp_mux2es #(3)    out_mux10(.dout(b10_outmx[2:0]),
                        .in0(b10_in0[2:0]),
                        .in1(b10_in1[2:0]),
                        .sel(~head));
  dp_mux2es #(3)    out_mux11(.dout(b11_outmx[2:0]),
                        .in0(b11_in0[2:0]),
                        .in1(b11_in1[2:0]),
                        .sel(~head));
  dp_mux2es #(3)    out_mux12(.dout(b12_outmx[2:0]),
                        .in0(b12_in0[2:0]),
                        .in1(b12_in1[2:0]),
                        .sel(~head));
  dp_mux2es #(3)    out_mux13(.dout(b13_outmx[2:0]),
                        .in0(b13_in0[2:0]),
                        .in1(b13_in1[2:0]),
                        .sel(~head));
  dp_mux2es #(3)    out_mux14(.dout(b14_outmx[2:0]),
                        .in0(b14_in0[2:0]),
                        .in1(b14_in1[2:0]),
                        .sel(~head));
  dp_mux2es #(3)    out_mux15(.dout(b15_outmx[2:0]),
                        .in0(b15_in0[2:0]),
                        .in1(b15_in1[2:0]),
                        .sel(~head));
  dp_mux2es         out_mux16(.dout(b16_outmx),
                        .in0(1'b0),
                        .in1(b16_in1),
                        .sel(~head));
  dff_s #(3)    out_dff0 (.din(b0_outmx[2:0]), .clk(clk_enb0), .q(b0[2:0]),
			.se(se), .si(), .so());
  dff_s #(3)    out_dff1 (.din(b1_outmx[2:0]), .clk(clk_enb0), .q(b1[2:0]),
			.se(se), .si(), .so());
  dff_s #(3)    out_dff2 (.din(b2_outmx[2:0]), .clk(clk_enb0), .q(b2[2:0]),
			.se(se), .si(), .so());
  dff_s #(3)    out_dff3 (.din(b3_outmx[2:0]), .clk(clk_enb0), .q(b3[2:0]),
			.se(se), .si(), .so());
  dff_s #(3)    out_dff4 (.din(b4_outmx[2:0]), .clk(clk_enb0), .q(b4[2:0]),
			.se(se), .si(), .so());
  dff_s #(3)    out_dff5 (.din(b5_outmx[2:0]), .clk(clk_enb0), .q(b5[2:0]),
			.se(se), .si(), .so());
  dff_s #(3)    out_dff6 (.din(b6_outmx[2:0]), .clk(clk_enb0), .q(b6[2:0]),
			.se(se), .si(), .so());
  dff_s #(3)    out_dff7 (.din(b7_outmx[2:0]), .clk(clk_enb0), .q(b7[2:0]),
			.se(se), .si(), .so());
  dff_s #(3)    out_dff8 (.din(b8_outmx[2:0]), .clk(clk_enb0), .q(b8[2:0]),
			.se(se), .si(), .so());
  dff_s #(3)    out_dff9 (.din(b9_outmx[2:0]), .clk(clk_enb0), .q(b9[2:0]),
			.se(se), .si(), .so());
  dff_s #(3)    out_dff10 (.din(b10_outmx[2:0]), .clk(clk_enb0), .q(b10[2:0]),
			.se(se), .si(), .so());
  dff_s #(3)    out_dff11 (.din(b11_outmx[2:0]), .clk(clk_enb0), .q(b11[2:0]),
			.se(se), .si(), .so());
  dff_s #(3)    out_dff12 (.din(b12_outmx[2:0]), .clk(clk_enb0), .q(b12[2:0]),
			.se(se), .si(), .so());
  dff_s #(3)    out_dff13 (.din(b13_outmx[2:0]), .clk(clk_enb0), .q(b13[2:0]),
			.se(se), .si(), .so());
  dff_s #(3)    out_dff14 (.din(b14_outmx[2:0]), .clk(clk_enb0), .q(b14[2:0]),
			.se(se), .si(), .so());
  dff_s #(3)    out_dff15 (.din(b15_outmx[2:0]), .clk(clk_enb0), .q(b15[2:0]),
			.se(se), .si(), .so());
  dff_s 	      out_dff16 (.din(b16_outmx), .clk(clk_enb0), .q(b16),
			.se(se), .si(), .so());
endmodule 
module mul_bodec (x, b,  
        b0, b1, b2, b3, b4, b5, b6, b7);
input	x;
input   [15:0] 	b;
output  [2:0] 	b0, b1, b2, b3, b4, b5, b6, b7; 
assign b0[2] = b[1];
assign b0[1] = ~((b[1] & b[0] & x) | (~b[1] & ~b[0] & ~x)) ;
assign b0[0] = (~b[1] & b[0] & x) | (b[1] & ~b[0] & ~x) ;
assign b1[2] = b[3]; 
assign b1[1] = ~((b[3] & b[2] & b[1]) | (~b[3] & ~b[2] & ~b[1])) ;
assign b1[0] = (~b[3] & b[2] & b[1]) | (b[3] & ~b[2] & ~b[1]) ;
assign b2[2] = b[5]; 
assign b2[1] = ~((b[5] & b[4] & b[3]) | (~b[5] & ~b[4] & ~b[3])) ;
assign b2[0] = (~b[5] & b[4] & b[3]) | (b[5] & ~b[4] & ~b[3]) ;
assign b3[2] = b[7] ;
assign b3[1] = ~((b[7] & b[6] & b[5]) | (~b[7] & ~b[6] & ~b[5])) ;
assign b3[0] = (~b[7] & b[6] & b[5]) | (b[7] & ~b[6] & ~b[5]) ;
assign b4[2] = b[9] ;
assign b4[1] = ~((b[9] & b[8] & b[7]) | (~b[9] & ~b[8] & ~b[7])) ;
assign b4[0] = (~b[9] & b[8] & b[7]) | (b[9] & ~b[8] & ~b[7]) ;
assign b5[2] = b[11] ;
assign b5[1] = ~((b[11] & b[10] & b[9]) | (~b[11] & ~b[10] & ~b[9])) ;
assign b5[0] = (~b[11] & b[10] & b[9]) | (b[11] & ~b[10] & ~b[9]) ;
assign b6[2] = b[13] ;
assign b6[1] = ~((b[13] & b[12] & b[11]) | (~b[13] & ~b[12] & ~b[11])) ;
assign b6[0] = (~b[13] & b[12] & b[11]) | (b[13] & ~b[12] & ~b[11]) ;
assign b7[2] = b[15] ;
assign b7[1] = ~((b[15] & b[14] & b[13]) | (~b[15] & ~b[14] & ~b[13])) ;
assign b7[0] = (~b[15] & b[14] & b[13]) | (b[15] & ~b[14] & ~b[13]) ;
endmodule 
                 
 
module dff_s (din, clk, q, se, si, so);
parameter SIZE = 1;
input	[SIZE-1:0]	din ;	
input			clk ;	
output	[SIZE-1:0]	q ;	
input			se ;	
input	[SIZE-1:0]	si ;	
output	[SIZE-1:0]	so ;	
reg 	[SIZE-1:0]	q ;
always @ (posedge clk)
  q[SIZE-1:0]  <= din[SIZE-1:0] ;
endmodule 
module dff_sscan (din, clk, q, se, si, so);
parameter SIZE = 1;
input	[SIZE-1:0]	din ;	
input			clk ;	
output	[SIZE-1:0]	q ;	
input			se ;	
input	[SIZE-1:0]	si ;	
output	[SIZE-1:0]	so ;	
reg 	[SIZE-1:0]	q ;
always @ (posedge clk)
  q[SIZE-1:0]  <= din[SIZE-1:0] ;
assign so={SIZE{1'b0}};
endmodule 
module dff_ns (din, clk, q);
parameter SIZE = 1;
input	[SIZE-1:0]	din ;	
input			clk ;	
output	[SIZE-1:0]	q ;	
reg 	[SIZE-1:0]	q ;
always @ (posedge clk)
	q[SIZE-1:0]  <= din[SIZE-1:0] ;
endmodule 
module dffr_s (din, clk, rst, q, se, si, so);
parameter SIZE = 1;
input	[SIZE-1:0]	din ;	
input			clk ;	
input			rst ;	
output	[SIZE-1:0]	q ;	
input			se ;	
input	[SIZE-1:0]	si ;	
output	[SIZE-1:0]	so ;	
reg 	[SIZE-1:0]	q ;
always @ (posedge clk)
	q[SIZE-1:0]  <= ((rst) ? {SIZE{1'b0}}  : din[SIZE-1:0] );
endmodule 
module dffrl_s (din, clk, rst_l, q, se, si, so);
parameter SIZE = 1;
input	[SIZE-1:0]	din ;	
input			clk ;	
input			rst_l ;	
output	[SIZE-1:0]	q ;	
input			se ;	
input	[SIZE-1:0]	si ;	
output	[SIZE-1:0]	so ;	
reg 	[SIZE-1:0]	q ;
always @ (posedge clk)
	q[SIZE-1:0]  <= rst_l ? din[SIZE-1:0] : {SIZE{1'b0}};
endmodule 
module dffr_ns (din, clk, rst, q);
parameter SIZE = 1;
input	[SIZE-1:0]	din ;	
input			clk ;	
input			rst ;	
output	[SIZE-1:0]	q ;	
reg 	[SIZE-1:0]	q ;
always @ (posedge clk)
  q[SIZE-1:0] <= rst ? {SIZE{1'b0}} : din[SIZE-1:0];
   
endmodule 
module dffrl_ns (din, clk, rst_l, q);
parameter SIZE = 1;
input	[SIZE-1:0]	din ;	
input			clk ;	
input			rst_l ;	
output	[SIZE-1:0]	q ;	
reg 	[SIZE-1:0]	q ;
always @ (posedge clk)
  q[SIZE-1:0] <= rst_l ? din[SIZE-1:0] : {SIZE{1'b0}};
endmodule 
module dffe_s (din, en, clk, q, se, si, so);
parameter SIZE = 1;
input	[SIZE-1:0]	din ;	
input			en ;	
input			clk ;	
output	[SIZE-1:0]	q ;	
input			se ;	
input	[SIZE-1:0]	si ;	
output	[SIZE-1:0]	so ;	
reg 	[SIZE-1:0]	q ;
always @ (posedge clk)
	q[SIZE-1:0]  <= ((en) ? din[SIZE-1:0] : q[SIZE-1:0]) ;
endmodule 
module dffe_ns (din, en, clk, q);
parameter SIZE = 1;
input	[SIZE-1:0]	din ;	
input			en ;	
input			clk ;	
output	[SIZE-1:0]	q ;	
reg 	[SIZE-1:0]	q ;
always @ (posedge clk)
  q[SIZE-1:0] <= en ? din[SIZE-1:0] : q[SIZE-1:0];
endmodule 
module dffre_s (din, rst, en, clk, q, se, si, so);
parameter SIZE = 1;
input	[SIZE-1:0]	din ;	
input			en ;	
input			rst ;	
input			clk ;	
output	[SIZE-1:0]	q ;	
input			se ;	
input	[SIZE-1:0]	si ;	
output	[SIZE-1:0]	so ;	
reg 	[SIZE-1:0]	q ;
always @ (posedge clk)
	q[SIZE-1:0]  <= (rst ? {SIZE{1'b0}} : ((en) ? din[SIZE-1:0] : q[SIZE-1:0])) ;
endmodule 
module dffrle_s (din, rst_l, en, clk, q, se, si, so);
parameter SIZE = 1;
input	[SIZE-1:0]	din ;	
input			en ;	
input			rst_l ;	
input			clk ;	
output	[SIZE-1:0]	q ;	
input			se ;	
input	[SIZE-1:0]	si ;	
output	[SIZE-1:0]	so ;	
reg 	[SIZE-1:0]	q ;
always @ (posedge clk)
	 q[SIZE-1:0]  <= (rst_l ? ((en) ? din[SIZE-1:0] : q[SIZE-1:0]) : {SIZE{1'b0}}) ;
endmodule 
module dffre_ns (din, rst, en, clk, q);
parameter SIZE = 1;
input	[SIZE-1:0]	din ;	
input			en ;	
input			rst ;	
input			clk ;	
output	[SIZE-1:0]	q ;	
reg 	[SIZE-1:0]	q ;
always @ (posedge clk)
  q[SIZE-1:0] <= rst ? {SIZE{1'b0}} : ((en) ? din[SIZE-1:0] : q[SIZE-1:0]);
endmodule 
module dffrle_ns (din, rst_l, en, clk, q);
parameter SIZE = 1;
input	[SIZE-1:0]	din ;	
input			en ;	
input			rst_l ;	
input			clk ;	
output	[SIZE-1:0]	q ;	
reg 	[SIZE-1:0]	q ;
always @ (posedge clk)
  q[SIZE-1:0] <= rst_l ? ((en) ? din[SIZE-1:0] : q[SIZE-1:0]) : {SIZE{1'b0}} ;
endmodule 
module dffr_async (din, clk, rst, q, se, si, so);
parameter SIZE = 1;
input   [SIZE-1:0]      din ;   
input                   clk ;   
input                   rst ;   
output  [SIZE-1:0]      q ;     
input                   se ;    
input   [SIZE-1:0]      si ;    
output  [SIZE-1:0]      so ;    
reg     [SIZE-1:0]      q ;
always @ (posedge clk or posedge rst)
	q[SIZE-1:0]  <= rst ? {SIZE{1'b0}} : din[SIZE-1:0];
endmodule 
module dffrl_async (din, clk, rst_l, q, se, si, so);
parameter SIZE = 1;
input   [SIZE-1:0]      din ;   
input                   clk ;   
input                   rst_l ;   
output  [SIZE-1:0]      q ;     
input                   se ;    
input   [SIZE-1:0]      si ;    
output  [SIZE-1:0]      so ;    
reg     [SIZE-1:0]      q ;
always @ (posedge clk or negedge rst_l)
 
   q[SIZE-1:0]  <= (!rst_l) ? {SIZE{1'b0}} : din[SIZE-1:0];
 
 
endmodule 
module dffrl_async_ns (din, clk, rst_l, q);
parameter SIZE = 1;
input   [SIZE-1:0]      din ;   
input                   clk ;   
input                   rst_l ;   
output  [SIZE-1:0]      q ;     
 reg [SIZE-1:0] q;   
always @ (posedge clk or negedge rst_l) begin
 
    q[SIZE-1:0] <= ~rst_l ?  {SIZE{1'b0}} : ({SIZE{rst_l}} & din[SIZE-1:0]);
 
 
end
endmodule 
module mux2ds (dout, in0, in1, sel0, sel1) ;
parameter SIZE = 1;
output 	[SIZE-1:0] 	dout;
input	[SIZE-1:0]	in0;
input	[SIZE-1:0]	in1;
input			sel0;
input			sel1;
reg	[SIZE-1:0]	dout ;
wire [1:0] sel = {sel1, sel0}; 
   
always @ (sel0 or sel1 or in0 or in1)
	case ({sel1,sel0}) 
		2'b01 :	dout = in0 ;
		2'b10 : dout = in1 ;
		2'b11 : dout = {SIZE{1'bx}} ;
		2'b00 : dout = {SIZE{1'bx}} ;
			
			
			
			
			
			
			
			
			
			
			
		default : dout = {SIZE{1'bx}};
	endcase
endmodule 
module mux3ds (dout, in0, in1, in2, sel0, sel1, sel2) ;
parameter SIZE = 1;
output 	[SIZE-1:0] 	dout;
input	[SIZE-1:0]	in0;
input	[SIZE-1:0]	in1;
input	[SIZE-1:0]	in2;
input			sel0;
input			sel1;
input			sel2;
reg	[SIZE-1:0]	dout ;
wire [2:0] sel = {sel2,sel1,sel0}; 
   
always @ (sel0 or sel1 or sel2 or in0 or in1 or in2)
	case ({sel2,sel1,sel0}) 
		3'b001 : dout = in0 ;
		3'b010 : dout = in1 ;
		3'b100 : dout = in2 ;
		3'b000 : dout = {SIZE{1'bx}} ;
		3'b011 : dout = {SIZE{1'bx}} ;
		3'b101 : dout = {SIZE{1'bx}} ;
		3'b110 : dout = {SIZE{1'bx}} ;
		3'b111 : dout = {SIZE{1'bx}} ;
		default : dout = {SIZE{1'bx}};
			
	endcase
endmodule 
module mux4ds (dout, in0, in1, in2, in3, sel0, sel1, sel2, sel3) ;
parameter SIZE = 1;
output 	[SIZE-1:0] 	dout;
input	[SIZE-1:0]	in0;
input	[SIZE-1:0]	in1;
input	[SIZE-1:0]	in2;
input	[SIZE-1:0]	in3;
input			sel0;
input			sel1;
input			sel2;
input			sel3;
reg	[SIZE-1:0]	dout ;
   
wire [3:0] sel = {sel3,sel2,sel1,sel0}; 
   
always @ (sel0 or sel1 or sel2 or sel3 or in0 or in1 or in2 or in3)
	case ({sel3,sel2,sel1,sel0}) 
		4'b0001 : dout = in0 ;
		4'b0010 : dout = in1 ;
		4'b0100 : dout = in2 ;
		4'b1000 : dout = in3 ;
		4'b0000 : dout = {SIZE{1'bx}} ;
		4'b0011 : dout = {SIZE{1'bx}} ;
		4'b0101 : dout = {SIZE{1'bx}} ;
		4'b0110 : dout = {SIZE{1'bx}} ;
		4'b0111 : dout = {SIZE{1'bx}} ;
		4'b1001 : dout = {SIZE{1'bx}} ;
		4'b1010 : dout = {SIZE{1'bx}} ;
		4'b1011 : dout = {SIZE{1'bx}} ;
		4'b1100 : dout = {SIZE{1'bx}} ;
		4'b1101 : dout = {SIZE{1'bx}} ;
		4'b1110 : dout = {SIZE{1'bx}} ;
		4'b1111 : dout = {SIZE{1'bx}} ;
		default : dout = {SIZE{1'bx}};
			
	endcase
endmodule 
module sink (in);
parameter SIZE = 1;
input [SIZE-1:0] in;
   
   
   wire    a;
   assign		a = | in;
endmodule 
module source (out) ;
parameter SIZE = 1;
output  [SIZE-1:0] out;
assign  out = {SIZE{1'b0}};
endmodule 
module clken_buf (clk, rclk, enb_l, tmb_l);
output clk;
input  rclk, enb_l, tmb_l;
reg    clken;
  always @ (rclk or enb_l or tmb_l)
    if (!rclk)  
      clken = !enb_l | !tmb_l;
  assign clk = clken & rclk;
endmodule
module dffsl_ns (din, clk, set_l, q);
parameter SIZE = 1;
input   [SIZE-1:0]      din ;   
input                   clk ;   
input                   set_l ; 
output  [SIZE-1:0]      q ;     
reg     [SIZE-1:0]      q ;
always @ (posedge clk)
  q[SIZE-1:0] <= set_l ? din[SIZE-1:0] : {SIZE{1'b1}};
endmodule 
module dffsl_async_ns (din, clk, set_l, q);
parameter SIZE = 1;
input   [SIZE-1:0]      din ;   
input                   clk ;   
input                   set_l ; 
output  [SIZE-1:0]      q ;     
reg     [SIZE-1:0]      q ;
always @ (posedge clk or negedge set_l) begin
   q[SIZE-1:0] <= ~set_l ? {SIZE{1'b1}} : ({SIZE{~set_l}} | din[SIZE-1:0]);
end
endmodule 
module dffr_ns_r1 (din, clk, rst, q);
parameter SIZE = 1;
input   [SIZE-1:0]      din ;   
input                   clk ;   
input                   rst ;   
output  [SIZE-1:0]      q ;     
reg     [SIZE-1:0]      q ;
always @ (posedge clk)
  q[SIZE-1:0] <= rst ? {SIZE{1'b1}} : din[SIZE-1:0];
endmodule 
module dffr_async_ns (din, clk, rst, q);
parameter SIZE = 1;
input   [SIZE-1:0]      din ;   
input                   clk ;   
input                   rst;   
output  [SIZE-1:0]      q ;     
reg     [SIZE-1:0]      q ;
always @ (posedge clk or posedge rst)
  q[SIZE-1:0] <= rst ? {SIZE{1'b0}} : din[SIZE-1:0];
endmodule 
module dffr_async_ns_r1 (din, clk, rst, q);
parameter SIZE = 1;
input   [SIZE-1:0]      din ;   
input                   clk ;   
input                   rst;   
output  [SIZE-1:0]      q ;     
reg     [SIZE-1:0]      q ;
always @ (posedge clk or posedge rst)
  q[SIZE-1:0] <= rst ? {SIZE{1'b1}} : din[SIZE-1:0];
endmodule 
module dffr_async_ns_cl_r1 (din, clkl, rst, q);
parameter SIZE = 1;
input   [SIZE-1:0]      din ;   
input                   clkl ;  
input                   rst ;   
output  [SIZE-1:0]      q ;     
reg     [SIZE-1:0]      q ;
always @ (negedge clkl or posedge rst)
  q[SIZE-1:0] <= rst ? {SIZE{1'b1}} : din[SIZE-1:0];
endmodule 
module dp_mux2es (dout, in0, in1, sel) ;
parameter SIZE = 1;
output 	[SIZE-1:0] 	dout;
input	[SIZE-1:0]	in0;
input	[SIZE-1:0]	in1;
input			sel;
reg	[SIZE-1:0]	dout ;
always @ (sel or in0 or in1)
 begin
	   case (sel)
	     1'b1: dout = in1 ; 
	     1'b0: dout = in0;
	     default: 
         begin
            if (in0 == in1) begin
               dout = in0;
            end
            else
              dout = {SIZE{1'bx}};
         end
	   endcase 
 end
endmodule 
module dp_mux4ds (dout, in0, in1, in2, in3, 
		     sel0_l, sel1_l, sel2_l, sel3_l) ;
parameter SIZE = 1;
output 	[SIZE-1:0] 	dout;
input	[SIZE-1:0]	in0;
input	[SIZE-1:0]	in1;
input	[SIZE-1:0]	in2;
input	[SIZE-1:0]	in3;
input			sel0_l;
input			sel1_l;
input			sel2_l;
input			sel3_l;
reg	[SIZE-1:0]	dout ;
wire [3:0] sel = {sel3_l,sel2_l,sel1_l,sel0_l}; 
   
always @ (sel0_l or sel1_l or sel2_l or sel3_l or in0 or in1 or in2 or in3)
	case ({sel3_l,sel2_l,sel1_l,sel0_l})
		4'b1110 : dout = in0 ;
		4'b1101 : dout = in1 ;
		4'b1011 : dout = in2 ;
		4'b0111 : dout = in3 ;
		4'b1111 : dout = {SIZE{1'bx}} ;
		default : dout = {SIZE{1'bx}} ;
	endcase
endmodule 
module dp_mux5ds (dout, in0, in1, in2, in3,  in4,
		     sel0_l, sel1_l, sel2_l, sel3_l, sel4_l) ;
parameter SIZE = 1;
output 	[SIZE-1:0] 	dout;
input	[SIZE-1:0]	in0;
input	[SIZE-1:0]	in1;
input	[SIZE-1:0]	in2;
input	[SIZE-1:0]	in3;
input	[SIZE-1:0]	in4;
input			sel0_l;
input			sel1_l;
input			sel2_l;
input			sel3_l;
input			sel4_l;
reg	[SIZE-1:0]	dout ;
   
wire [4:0] sel = {sel4_l,sel3_l,sel2_l,sel1_l,sel0_l}; 
always @ (sel0_l or sel1_l or sel2_l or sel3_l or sel4_l or
		in0 or in1 or in2 or in3 or in4)
	case ({sel4_l,sel3_l,sel2_l,sel1_l,sel0_l})
		5'b11110 : dout = in0 ;
		5'b11101 : dout = in1 ;
		5'b11011 : dout = in2 ;
		5'b10111 : dout = in3 ;
		5'b01111 : dout = in4 ;
		5'b11111 : dout = {SIZE{1'bx}} ;
		default : dout = {SIZE{1'bx}} ;
	endcase
endmodule 
module dp_mux8ds (dout, in0, in1, in2, in3, 
			in4, in5, in6, in7,
		     sel0_l, sel1_l, sel2_l, sel3_l,
		     sel4_l, sel5_l, sel6_l, sel7_l) ;
parameter SIZE = 1;
output 	[SIZE-1:0] 	dout;
input	[SIZE-1:0]	in0;
input	[SIZE-1:0]	in1;
input	[SIZE-1:0]	in2;
input	[SIZE-1:0]	in3;
input	[SIZE-1:0]	in4;
input	[SIZE-1:0]	in5;
input	[SIZE-1:0]	in6;
input	[SIZE-1:0]	in7;
input			sel0_l;
input			sel1_l;
input			sel2_l;
input			sel3_l;
input			sel4_l;
input			sel5_l;
input			sel6_l;
input			sel7_l;
reg	[SIZE-1:0]	dout ;
wire [7:0] sel = {sel7_l,sel6_l,sel5_l,sel4_l,
                  sel3_l,sel2_l,sel1_l,sel0_l}; 
always @ (sel0_l or sel1_l or sel2_l or sel3_l or in0 or in1 or in2 or in3 or
	  sel4_l or sel5_l or sel6_l or sel7_l or in4 or in5 or in6 or in7)
	case ({sel7_l,sel6_l,sel5_l,sel4_l,sel3_l,sel2_l,sel1_l,sel0_l})
		8'b11111110 : dout = in0 ;
		8'b11111101 : dout = in1 ;
		8'b11111011 : dout = in2 ;
		8'b11110111 : dout = in3 ;
		8'b11101111 : dout = in4 ;
		8'b11011111 : dout = in5 ;
		8'b10111111 : dout = in6 ;
		8'b01111111 : dout = in7 ;
		8'b11111111 : dout = {SIZE{1'bx}} ;
		default : dout = {SIZE{1'bx}} ;
	endcase
endmodule 
module dp_mux3ds (dout, in0, in1, in2, 
		     sel0_l, sel1_l, sel2_l);
parameter SIZE = 1;
output 	[SIZE-1:0] 	dout;
input	[SIZE-1:0]	in0;
input	[SIZE-1:0]	in1;
input	[SIZE-1:0]	in2;
input			sel0_l;
input			sel1_l;
input			sel2_l;
reg	[SIZE-1:0]	dout ;
wire [2:0] sel = {sel2_l,sel1_l,sel0_l}; 
   
always @ (sel0_l or sel1_l or sel2_l or in0 or in1 or in2)
	case ({sel2_l,sel1_l,sel0_l})
		3'b110 : dout = in0 ;
		3'b101 : dout = in1 ;
		3'b011 : dout = in2 ;
	        default : dout = {SIZE{1'bx}} ;
	endcase
endmodule 
module dp_mux2ds (dout, in0, in1,
             sel0_l, sel1_l);
parameter SIZE = 1;
output  [SIZE-1:0]  dout;
input   [SIZE-1:0]  in0;
input   [SIZE-1:0]  in1;
input           sel0_l;
input           sel1_l;
reg [SIZE-1:0]  dout ;
wire [1:0] sel = {sel1_l,sel0_l}; 
always @ (sel0_l or sel1_l or in0 or in1)
    case ({sel1_l,sel0_l})
        3'b10 : dout = in0 ;
        3'b01 : dout = in1 ;
            default : dout = {SIZE{1'bx}} ;
    endcase
endmodule 
module dp_buffer(dout, in);
parameter SIZE = 1;
output 	[SIZE-1:0] 	dout;
input	[SIZE-1:0]	in;
assign dout = in;
endmodule 
module test_stub_scan (
mux_drive_disable, mem_write_disable, sehold, se, testmode_l, 
mem_bypass, so_0, so_1, so_2, 
ctu_tst_pre_grst_l, arst_l, global_shift_enable, 
ctu_tst_scan_disable, ctu_tst_scanmode, ctu_tst_macrotest, 
ctu_tst_short_chain, long_chain_so_0, short_chain_so_0, 
long_chain_so_1, short_chain_so_1, long_chain_so_2, short_chain_so_2
);
   input        ctu_tst_pre_grst_l;
   input        arst_l;                
   input        global_shift_enable;
   input        ctu_tst_scan_disable;  
   input        ctu_tst_scanmode;
   input 	ctu_tst_macrotest;
   input 	ctu_tst_short_chain;
   input 	long_chain_so_0;
   input 	short_chain_so_0;
   input 	long_chain_so_1;
   input 	short_chain_so_1;
   input 	long_chain_so_2;
   input 	short_chain_so_2;
   
   output 	mux_drive_disable;
   output 	mem_write_disable;
   output 	sehold;
   output 	se;
   output 	testmode_l;
   output 	mem_bypass;
   output 	so_0;
   output 	so_1;
   output 	so_2;
   wire         pin_based_scan;
   wire         short_chain_en;
   wire         short_chain_select;
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   assign  mux_drive_disable  = ~ctu_tst_pre_grst_l | short_chain_select | se;
   assign  mem_write_disable  = ~ctu_tst_pre_grst_l | se;
   assign  sehold             = ctu_tst_macrotest & ~se;
   assign  se                 = global_shift_enable;
   assign  testmode_l         = ~ctu_tst_scanmode;
   assign  mem_bypass         = ~ctu_tst_macrotest & ~testmode_l;
   assign  pin_based_scan     = ctu_tst_scan_disable;
   assign  short_chain_en     = ~(pin_based_scan & se);
   assign  short_chain_select = ctu_tst_short_chain & ~testmode_l & short_chain_en;
   assign  so_0               = short_chain_select ? short_chain_so_0 : long_chain_so_0;
   assign  so_1               = short_chain_select ? short_chain_so_1 : long_chain_so_1;
   assign  so_2               = short_chain_select ? short_chain_so_2 : long_chain_so_2;
   
endmodule 
module bw_u1_inv_0p6x (
    z,
    a );
    output z;
    input  a;
    assign z = ~( a );
endmodule
module bw_u1_inv_1x (
    z,
    a );
    output z;
    input  a;
    assign z = ~( a );
endmodule
module bw_u1_inv_1p4x (
    z,
    a );
    output z;
    input  a;
    assign z = ~( a );
endmodule
module bw_u1_inv_2x (
    z,
    a );
    output z;
    input  a;
    assign z = ~( a );
endmodule
module bw_u1_inv_3x (
    z,
    a );
    output z;
    input  a;
    assign z = ~( a );
endmodule
module bw_u1_inv_4x (
    z,
    a );
    output z;
    input  a;
    assign z = ~( a );
endmodule
module bw_u1_inv_5x (
    z,
    a );
    output z;
    input  a;
    assign z = ~( a );
endmodule
module bw_u1_inv_8x (
    z,
    a );
    output z;
    input  a;
    assign z = ~( a );
endmodule
module bw_u1_inv_10x (
    z,
    a );
    output z;
    input  a;
    assign z = ~( a );
endmodule
module bw_u1_inv_15x (
    z,
    a );
    output z;
    input  a;
    assign z = ~( a );
endmodule
module bw_u1_inv_20x (
    z,
    a );
    output z;
    input  a;
    assign z = ~( a );
endmodule
module bw_u1_inv_30x (
    z,
    a );
    output z;
    input  a;
    assign z = ~( a );
endmodule
module bw_u1_inv_40x (
    z,
    a );
    output z;
    input  a;
    assign z = ~( a );
endmodule
module bw_u1_invh_15x (
    z,
    a );
    output z;
    input  a;
    assign z = ~( a );
endmodule
module bw_u1_invh_25x (
    z,
    a );
    output z;
    input  a;
    assign z = ~( a );
endmodule
module bw_u1_invh_30x (
    z,
    a );
    output z;
    input  a;
    assign z = ~( a );
endmodule
module bw_u1_invh_50x (
    z,
    a );
    output z;
    input  a;
    assign z = ~( a );
endmodule
module bw_u1_invh_60x (
    z,
    a );
    output z;
    input  a;
    assign z = ~( a );
endmodule
module bw_u1_nand2_0p4x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a & b );
endmodule
module bw_u1_nand2_0p6x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a & b );
endmodule
module bw_u1_nand2_1x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a & b );
endmodule
module bw_u1_nand2_1p4x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a & b );
endmodule
module bw_u1_nand2_2x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a & b );
endmodule
module bw_u1_nand2_3x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a & b );
endmodule
module bw_u1_nand2_4x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a & b );
endmodule
module bw_u1_nand2_5x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a & b );
endmodule
module bw_u1_nand2_7x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a & b );
endmodule
module bw_u1_nand2_10x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a & b );
endmodule
module bw_u1_nand2_15x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a & b );
endmodule
module bw_u1_nand3_0p4x (
    z,
    a,
    b,
    c );
    output z;
    input  a;
    input  b;
    input  c;
    assign z = ~( a & b & c );
endmodule
module bw_u1_nand3_0p6x (
    z,
    a,
    b,
    c );
    output z;
    input  a;
    input  b;
    input  c;
    assign z = ~( a & b & c );
endmodule
module bw_u1_nand3_1x (
    z,
    a,  
    b,  
    c );
    
    output z;
    input  a;
    input  b;
    input  c;
    
    assign z = ~( a & b & c );
endmodule
module bw_u1_nand3_1p4x (
    z,
    a,  
    b,  
    c );
    
    output z;
    input  a;
    input  b;
    input  c;
    
    assign z = ~( a & b & c );
endmodule
module bw_u1_nand3_2x (
    z,
    a,  
    b,  
    c );
    
    output z;
    input  a;
    input  b;
    input  c;
    
    assign z = ~( a & b & c );
endmodule
module bw_u1_nand3_3x (
    z,
    a,  
    b,  
    c );
    
    output z;
    input  a;
    input  b;
    input  c;
    
    assign z = ~( a & b & c );
endmodule
module bw_u1_nand3_4x (
    z,
    a,  
    b,  
    c );
    
    output z;
    input  a;
    input  b;
    input  c;
    
    assign z = ~( a & b & c );
endmodule
module bw_u1_nand3_5x (
    z,
    a,  
    b,  
    c );
    
    output z;
    input  a;
    input  b;
    input  c;
    
    assign z = ~( a & b & c );
endmodule
module bw_u1_nand3_7x (
    z,
    a,  
    b,  
    c );
    
    output z;
    input  a;
    input  b;
    input  c;
    
    assign z = ~( a & b & c );
endmodule
module bw_u1_nand3_10x (
    z,
    a,  
    b,  
    c );
    
    output z;
    input  a;
    input  b;
    input  c;
    
    assign z = ~( a & b & c );
endmodule
module bw_u1_nand4_0p6x (
    z,
    a,  
    b,  
    c,  
    d );
    
    output z;
    input  a;
    input  b;
    input  c;
    input  d;
    
    assign z = ~( a & b & c & d );
endmodule
module bw_u1_nand4_1x (
    z,
    a,
    b,
    c,
    d );
    output z;
    input  a;
    input  b;
    input  c;
    input  d;
    assign z = ~( a & b & c & d );
endmodule
module bw_u1_nand4_1p4x (
    z,
    a,
    b,
    c,
    d );
    output z;
    input  a;
    input  b;
    input  c;
    input  d;
    assign z = ~( a & b & c & d );
endmodule
module bw_u1_nand4_2x (
    z,
    a,
    b,
    c,
    d );
    output z;
    input  a;
    input  b;
    input  c;
    input  d;
    assign z = ~( a & b & c & d );
endmodule
module bw_u1_nand4_3x (
    z,
    a,
    b,
    c,
    d );
    output z;
    input  a;
    input  b;
    input  c;
    input  d;
    assign z = ~( a & b & c & d );
endmodule
module bw_u1_nand4_4x (
    z,
    a,
    b,
    c,
    d );
    output z;
    input  a;
    input  b;
    input  c;
    input  d;
    assign z = ~( a & b & c & d );
endmodule
module bw_u1_nand4_6x (
    z,
    a,
    b,
    c,
    d );
    output z;
    input  a;
    input  b;
    input  c;
    input  d;
    nand( z, a, b,c,d);
endmodule
module bw_u1_nand4_8x (
    z,
    a,
    b,
    c,
    d );
    output z;
    input  a;
    input  b;
    input  c;
    input  d;
    nand( z, a, b,c,d);
endmodule
module bw_u1_nor2_0p6x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a | b );
endmodule
module bw_u1_nor2_1x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a | b );
endmodule
module bw_u1_nor2_1p4x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a | b );
endmodule
module bw_u1_nor2_2x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a | b );
endmodule
module bw_u1_nor2_3x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a | b );
endmodule
module bw_u1_nor2_4x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a | b );
endmodule
module bw_u1_nor2_6x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a | b );
endmodule
module bw_u1_nor2_8x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a | b );
endmodule
module bw_u1_nor2_12x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a | b );
endmodule
module bw_u1_nor3_0p6x (
    z,
    a,
    b,
    c );
    output z;
    input  a;
    input  b;
    input  c;
    assign z = ~( a | b | c );
endmodule
module bw_u1_nor3_1x (
    z,
    a,
    b,
    c );
    output z;
    input  a;
    input  b;
    input  c;
    assign z = ~( a | b | c );
endmodule
module bw_u1_nor3_1p4x (
    z,
    a,
    b,
    c );
    output z;
    input  a;
    input  b;
    input  c;
    assign z = ~( a | b | c );
endmodule
module bw_u1_nor3_2x (
    z,
    a,
    b,
    c );
    output z;
    input  a;
    input  b;
    input  c;
    assign z = ~( a | b | c );
endmodule
module bw_u1_nor3_3x (
    z,
    a,
    b,
    c );
    output z;
    input  a;
    input  b;
    input  c;
    assign z = ~( a | b | c );
endmodule
module bw_u1_nor3_4x (
    z,
    a,
    b,
    c );
    output z;
    input  a;
    input  b;
    input  c;
    assign z = ~( a | b | c );
endmodule
module bw_u1_nor3_6x (
    z,
    a,
    b,
    c );
    output z;
    input  a;
    input  b;
    input  c;
    assign z = ~( a | b | c );
endmodule
module bw_u1_nor3_8x (
    z,
    a,
    b,
    c );
    output z;
    input  a;
    input  b;
    input  c;
    assign z = ~( a | b | c );
endmodule
module bw_u1_aoi21_0p4x (
    z,
    b1,
    b2,
    a );
    output z;
    input  b1;
    input  b2;
    input  a;
    assign z = ~(( b1 & b2 ) | ( a ));
endmodule
module bw_u1_aoi21_1x (
    z,
    b1,
    b2,
    a );
    output z;
    input  b1;
    input  b2;
    input  a;
    assign z = ~(( b1 & b2 ) | ( a  ));
endmodule
module bw_u1_aoi21_2x (
    z,
    b1,
    b2,
    a );
    output z;
    input  b1;
    input  b2;
    input  a;
    assign z = ~(( b1 & b2 ) | ( a ));
endmodule
module bw_u1_aoi21_4x (
    z,
    b1,
    b2,
    a );
    output z;
    input  b1;
    input  b2;
    input  a;
    assign z = ~(( b1 & b2 ) | ( a ));
endmodule
module bw_u1_aoi21_8x (
    z,
    b1,
    b2,
    a );
    output z;
    input  b1;
    input  b2;
    input  a;
    assign z = ~(( b1 & b2 ) | ( a ));
endmodule
module bw_u1_aoi21_12x (
    z,
    b1,
    b2,
    a );
    output z;
    input  b1;
    input  b2;
    input  a;
    assign z = ~(( b1 & b2 ) | ( a ));
endmodule
module bw_u1_aoi22_0p4x (
    z,
    a1,
    a2,
    b1,
    b2 );
    output z;
    input  a1;
    input  a2;
    input  b1;
    input  b2;
    assign z = ~(( a1 & a2 ) | ( b1 & b2 ));
endmodule
module bw_u1_aoi22_1x (
    z,
    b1,
    b2,
    a1,
    a2 );
    output z;
    input  b1;
    input  b2;
    input  a1;
    input  a2;
    assign z = ~(( a1 & a2 ) | ( b1 & b2 ));
endmodule
module bw_u1_aoi22_2x (
    z,
    b1,
    b2,
    a1,
    a2 );
    output z;
    input  b1;
    input  b2;
    input  a1;
    input  a2;
 
    assign z = ~(( a1 & a2 ) | ( b1 & b2 ));
endmodule
module bw_u1_aoi22_4x (
    z,
    b1,
    b2,
    a1,
    a2 );
    output z;
    input  b1;
    input  b2;
    input  a1;
    input  a2;
    assign z = ~(( a1 & a2 ) | ( b1 & b2 ));
endmodule
module bw_u1_aoi22_8x (
    z,
    b1,
    b2,
    a1,
    a2 );
    output z;
    input  b1;
    input  b2;
    input  a1;
    input  a2;
    assign z = ~(( a1 & a2 ) | ( b1 & b2 ));
endmodule
module bw_u1_aoi211_0p3x (
    z,
    c1,
    c2,
    b,
    a );
    output z;
    input  c1;
    input  c2;
    input  b;
    input  a;
    assign z = ~(( c1 & c2 ) | (a)| (b));
endmodule
module bw_u1_aoi211_1x (
    z,
    c1,
    c2,
    b,
    a );
    output z;
    input  c1;
    input  c2;
    input  b;
    input  a;
    assign z = ~(( c1 & c2 ) | (a)| (b));
endmodule
module bw_u1_aoi211_2x (
    z,
    c1,
    c2,
    b, 
    a );
    output z;
    input  c1;
    input  c2;
    input  b;
    input  a;
 
    assign z = ~(( c1 & c2 ) | (a)| (b));
endmodule
module bw_u1_aoi211_4x (
    z,
    c1,
    c2,
    b, 
    a );
    output z;
    input  c1;
    input  c2;
    input  b;
    input  a;
 
    assign z = ~(( c1 & c2 ) | (a)| (b));
endmodule
module bw_u1_aoi211_8x (
    z,
    c1,
    c2,
    b, 
    a );
    output z;
    input  c1;
    input  c2;
    input  b;
    input  a;
 
    assign z = ~(( c1 & c2 ) | (a)| (b));
endmodule
module bw_u1_oai21_0p4x (
    z,
    b1,
    b2,
    a );
    output z;
    input  b1;
    input  b2;
    input  a;
    assign z = ~(( b1 | b2 ) & ( a ));
endmodule
module bw_u1_oai21_1x (
    z,
    b1,
    b2,
    a );
    output z;
    input  b1;
    input  b2;
    input  a;
    assign z = ~(( b1 | b2 ) & ( a ));
endmodule
module bw_u1_oai21_2x (
    z,
    b1,
    b2,
    a );
    output z;
    input  b1;
    input  b2;
    input  a;
    assign z = ~(( b1 | b2 ) & ( a ));
endmodule
module bw_u1_oai21_4x (
    z,
    b1,
    b2,
    a );
    output z;
    input  b1;
    input  b2;
    input  a;
    assign z = ~(( b1 | b2 ) & ( a ));
endmodule
module bw_u1_oai21_8x (
    z,
    b1,
    b2,
    a );
    output z;
    input  b1;
    input  b2;
    input  a;
    assign z = ~(( b1 | b2 ) & ( a ));
endmodule
module bw_u1_oai21_12x (
    z,
    b1,
    b2,
    a );
    output z;
    input  b1;
    input  b2;
    input  a;
    assign z = ~(( b1 | b2 ) & ( a ));
endmodule
module bw_u1_oai22_0p4x (
    z,
    a1,
    a2,
    b1,
    b2 );
    output z;
    input  a1;
    input  a2;
    input  b1;
    input  b2;
    assign z = ~(( a1 | a2 ) & ( b1 | b2 ));
endmodule
module bw_u1_oai22_1x (
    z,
    a1,
    a2,
    b1,
    b2 );
    output z;
    input  a1;
    input  a2;
    input  b1;
    input  b2;
    assign z = ~(( a1 | a2 ) & ( b1 | b2 ));
endmodule
module bw_u1_oai22_2x (
    z,
    a1,
    a2,
    b1,
    b2 );
    output z;
    input  a1;
    input  a2;
    input  b1;
    input  b2;
    assign z = ~(( a1 | a2 ) & ( b1 | b2 ));
endmodule
module bw_u1_oai22_4x (
    z,
    a1,
    a2,
    b1,
    b2 );
    output z;
    input  a1;
    input  a2;
    input  b1;
    input  b2;
    assign z = ~(( a1 | a2 ) & ( b1 | b2 ));
endmodule
module bw_u1_oai22_8x (
    z,
    a1,
    a2,
    b1,
    b2 );
    output z;
    input  a1;
    input  a2;
    input  b1;
    input  b2;
    assign z = ~(( a1 | a2 ) & ( b1 | b2 ));
endmodule
module bw_u1_oai211_0p3x (
    z,
    c1,
    c2,
    b,
    a );
    output z;
    input  c1;
    input  c2;
    input  b;
    input  a;
    assign z = ~(( c1 | c2 ) & ( a ) & (b));
endmodule
module bw_u1_oai211_1x (
    z,
    c1,
    c2,
    b,
    a );
    output z;
    input  c1;
    input  c2;
    input  b;
    input  a;
    assign z = ~(( c1 | c2 ) & ( a ) & (b));
endmodule
module bw_u1_oai211_2x (
    z,
    c1,
    c2,
    b,
    a );
    output z;
    input  c1;
    input  c2;
    input  b;
    input  a;
    assign z = ~(( c1 | c2 ) & ( a ) & (b));
endmodule
module bw_u1_oai211_4x (
    z,
    c1,
    c2,
    b,
    a );
    output z;
    input  c1;
    input  c2;
    input  b;
    input  a;
    assign z = ~(( c1 | c2 ) & ( a ) & (b));
endmodule
module bw_u1_oai211_8x (
    z,
    c1,
    c2,
    b,
    a );
    output z;
    input  c1;
    input  c2;
    input  b;
    input  a;
    assign z = ~(( c1 | c2 ) & ( a ) & (b));
endmodule
module bw_u1_aoi31_1x (
    z,
    b1,
    b2,
    b3,
    a );
    output z;
    input  b1;
    input  b2;
    input  b3;
    input  a;
    assign z = ~(( b1 & b2&b3 ) | ( a ));
endmodule
module bw_u1_aoi31_2x (
    z, 
    b1,
    b2, 
    b3, 
    a );
    
    output z; 
    input  b1;
    input  b2;
    input  b3;
    input  a;
    assign z = ~(( b1 & b2&b3 ) | ( a ));
endmodule
module bw_u1_aoi31_4x (
    z, 
    b1,
    b2, 
    b3, 
    a );
    
    output z; 
    input  b1;
    input  b2;
    input  b3;
    input  a;
    assign z = ~(( b1 & b2&b3 ) | ( a ));
endmodule
module bw_u1_aoi31_8x (
    z, 
    b1,
    b2, 
    b3, 
    a );
    
    output z; 
    input  b1;
    input  b2;
    input  b3;
    input  a;
    assign z = ~(( b1 & b2&b3 ) | ( a ));
endmodule
module bw_u1_aoi32_1x (
    z,
    b1,
    b2,
    b3,
    a1,
    a2 );
    output z;
    input  b1;
    input  b2;
    input  b3;
    input  a1;
    input  a2;
    assign z = ~(( b1 & b2&b3 ) | ( a1 & a2 ));
endmodule
module bw_u1_aoi32_2x (
    z,
    b1, 
    b2,
    b3,
    a1,
    a2 );
    output z;
    input  b1; 
    input  b2; 
    input  b3; 
    input  a1;
    input  a2;
 
    assign z = ~(( b1 & b2&b3 ) | ( a1 & a2 ));
endmodule
module bw_u1_aoi32_4x (
    z,
    b1, 
    b2,
    b3,
    a1,
    a2 );
    output z;
    input  b1; 
    input  b2; 
    input  b3; 
    input  a1;
    input  a2;
 
    assign z = ~(( b1 & b2&b3 ) | ( a1 & a2 ));
endmodule
module bw_u1_aoi32_8x (
    z,
    b1, 
    b2,
    b3,
    a1,
    a2 );
    output z;
    input  b1; 
    input  b2; 
    input  b3; 
    input  a1;
    input  a2;
 
    assign z = ~(( b1 & b2&b3 ) | ( a1 & a2 ));
endmodule
module bw_u1_aoi33_1x (
    z,
    b1,
    b2,
    b3,
    a1,
    a2,
    a3 );
    output z;
    input  b1;
    input  b2;
    input  b3;
    input  a1;
    input  a2;
    input  a3;
    assign z = ~(( b1 & b2&b3 ) | ( a1&a2&a3 ));
endmodule
module bw_u1_aoi33_2x (
       
    z, 
    b1, 
    b2,  
    b3,  
    a1,  
    a2,  
    a3 );
    
    output z;
    input  b1;
    input  b2;
    input  b3;
    input  a1;
    input  a2;
    input  a3;
    
    assign z = ~(( b1 & b2&b3 ) | ( a1&a2&a3 ));
endmodule
module bw_u1_aoi33_4x (
       
    z, 
    b1, 
    b2,  
    b3,  
    a1,  
    a2,  
    a3 );
    
    output z;
    input  b1;
    input  b2;
    input  b3;
    input  a1;
    input  a2;
    input  a3;
    
    assign z = ~(( b1 & b2&b3 ) | ( a1&a2&a3 ));
endmodule
module bw_u1_aoi33_8x (
       
    z, 
    b1, 
    b2,  
    b3,  
    a1,  
    a2,  
    a3 );
    
    output z;
    input  b1;
    input  b2;
    input  b3;
    input  a1;
    input  a2;
    input  a3;
    
    assign z = ~(( b1 & b2&b3 ) | ( a1&a2&a3 ));
endmodule
module bw_u1_aoi221_1x (
    z,
    c1,
    c2,
    b1,
    b2,
    a );
    output z;
    input  c1;
    input  c2;
    input  b1;
    input  b2;
    input  a;
    assign z = ~(( c1 & c2 ) | (b1&b2)| (a));
endmodule
module bw_u1_aoi221_2x (
    z,
    c1,
    c2,
    b1,
    b2,
    a );
    output z;
    input  c1;
    input  c2;
    input  b1;
    input  b2;
    input  a; 
    assign z = ~(( c1 & c2 ) | (b1&b2)| (a));
endmodule
module bw_u1_aoi221_4x (
    z,
    c1,
    c2,
    b1,
    b2,
    a );
    output z;
    input  c1;
    input  c2;
    input  b1;
    input  b2;
    input  a; 
    assign z = ~(( c1 & c2 ) | (b1&b2)| (a));
endmodule
module bw_u1_aoi221_8x (
    z,
    c1,
    c2,
    b1,
    b2,
    a );
    output z;
    input  c1;
    input  c2;
    input  b1;
    input  b2;
    input  a; 
    assign z = ~(( c1 & c2 ) | (b1&b2)| (a));
endmodule
module bw_u1_aoi222_1x (
    z,
    a1,
    a2,
    b1,
    b2,
    c1,
    c2 );
    output z;
    input  a1;
    input  a2;
    input  b1;
    input  b2;
    input  c1;
    input  c2;
    assign z = ~(( c1 & c2 ) | (b1&b2)| (a1& a2));
endmodule
module bw_u1_aoi222_2x (
    z,
    a1,
    a2,
    b1,
    b2,
    c1,
    c2 );
    output z;
    input  a1;
    input  a2;
    input  b1;
    input  b2;
    input  c1;
    input  c2;
    assign z = ~(( c1 & c2 ) | (b1&b2)| (a1& a2));
endmodule
module bw_u1_aoi222_4x (
    z,
    a1,
    a2,
    b1,
    b2,
    c1,
    c2 );
    output z;
    input  a1;
    input  a2;
    input  b1;
    input  b2;
    input  c1;
    input  c2;
    assign z = ~(( c1 & c2 ) | (b1&b2)| (a1& a2));
endmodule
module bw_u1_aoi311_1x (
    z,
    c1,
    c2,
    c3,
    b, 
    a );
    output z;
    input  c1;
    input  c2;
    input  c3;
    input  b;
    input  a;
    assign z = ~(( c1 & c2& c3 ) | (a)| (b));
endmodule
module bw_u1_aoi311_2x (
    z,
    c1,
    c2,
    c3,
    b, 
    a );
    output z;
    input  c1;
    input  c2;
    input  c3;
    input  b;
    input  a;
    assign z = ~(( c1 & c2& c3 ) | (a)| (b));
endmodule
module bw_u1_aoi311_4x (
    z,
    c1,
    c2,
    c3,
    b, 
    a );
    output z;
    input  c1;
    input  c2;
    input  c3;
    input  b;
    input  a;
    assign z = ~(( c1 & c2& c3 ) | (a)| (b));
endmodule
module bw_u1_aoi311_8x (
    z,
    c1,
    c2,
    c3,
    b, 
    a );
    output z;
    input  c1;
    input  c2;
    input  c3;
    input  b;
    input  a;
    assign z = ~(( c1 & c2& c3 ) | (a)| (b));
endmodule
module bw_u1_oai31_1x (
    z,
    b1,
    b2,
    b3,
    a );
    output z;
    input  b1;
    input  b2;
    input  b3;
    input  a;
    assign z = ~(( b1 | b2|b3 ) & ( a ));
endmodule
module bw_u1_oai31_2x (
    z,
    b1,
    b2,
    b3,
    a );
    output z;
    input  b1;
    input  b2;
    input  b3;
    input  a;
    assign z = ~(( b1 | b2|b3 ) & ( a ));
endmodule
module bw_u1_oai31_4x (
    z,
    b1,
    b2,
    b3,
    a );
    output z;
    input  b1;
    input  b2;
    input  b3;
    input  a;
    assign z = ~(( b1 | b2|b3 ) & ( a ));
endmodule
module bw_u1_oai31_8x (
    z,
    b1,
    b2,
    b3,
    a );
    output z;
    input  b1;
    input  b2;
    input  b3;
    input  a;
    assign z = ~(( b1 | b2|b3 ) & ( a ));
endmodule
module bw_u1_oai32_1x (
    z,
    b1,
    b2,
    b3,
    a1,
    a2 );
    output z;
    input  b1;
    input  b2;
    input  b3;
    input  a1;
    input  a2;
    assign z = ~(( b1 | b2 | b3 ) & ( a1 | a2 ));
endmodule
module bw_u1_oai32_2x (
    z,
    b1,
    b2,
    b3,
    a1,
    a2 );
    output z;
    input  b1;
    input  b2;
    input  b3;
    input  a1;
    input  a2;
    assign z = ~(( b1 | b2 | b3 ) & ( a1 | a2 ));
endmodule
module bw_u1_oai32_4x (
    z,
    b1,
    b2,
    b3,
    a1,
    a2 );
    output z;
    input  b1;
    input  b2;
    input  b3;
    input  a1;
    input  a2;
    assign z = ~(( b1 | b2 | b3 ) & ( a1 | a2 ));
endmodule
module bw_u1_oai32_8x (
    z,
    b1,
    b2,
    b3,
    a1,
    a2 );
    output z;
    input  b1;
    input  b2;
    input  b3;
    input  a1;
    input  a2;
    assign z = ~(( b1 | b2 | b3 ) & ( a1 | a2 ));
endmodule
module bw_u1_oai33_1x (
    z,
    b1,
    b2,
    b3,
    a1,
    a2,
    a3 );
    output z;
    input  b1;
    input  b2;
    input  b3;
    input  a1;
    input  a2;
    input  a3;
    assign z = ~(( b1 | b2|b3 ) & ( a1|a2|a3 ));
endmodule
module bw_u1_oai33_2x (
    z,
    b1,
    b2,
    b3,
    a1,
    a2,
    a3 );
    output z;
    input  b1;
    input  b2;
    input  b3;
    input  a1;
    input  a2;
    input  a3;
    assign z = ~(( b1 | b2|b3 ) & ( a1|a2|a3 ));
endmodule
module bw_u1_oai33_4x (
    z,
    b1,
    b2,
    b3,
    a1,
    a2,
    a3 );
    output z;
    input  b1;
    input  b2;
    input  b3;
    input  a1;
    input  a2;
    input  a3;
    assign z = ~(( b1 | b2|b3 ) & ( a1|a2|a3 ));
endmodule
module bw_u1_oai33_8x (
    z,
    b1,
    b2,
    b3,
    a1,
    a2,
    a3 );
    output z;
    input  b1;
    input  b2;
    input  b3;
    input  a1;
    input  a2;
    input  a3;
    assign z = ~(( b1 | b2|b3 ) & ( a1|a2|a3 ));
endmodule
module bw_u1_oai221_1x (
    z,
    c1,
    c2,
    b1,
    b2,
    a );
    output z;
    input  c1;
    input  c2;
    input  b1;
    input  b2;
    input  a;
    assign z = ~(( c1 | c2 ) & ( a ) & (b1|b2));
endmodule
module bw_u1_oai221_2x (
    z,
    c1,
    c2,
    b1,
    b2,
    a );
    output z;
    input  c1;
    input  c2;
    input  b1;
    input  b2;
    input  a;
    assign z = ~(( c1 | c2 ) & ( a ) & (b1|b2));
endmodule
module bw_u1_oai221_4x (
    z,
    c1,
    c2,
    b1,
    b2,
    a );
    output z;
    input  c1;
    input  c2;
    input  b1;
    input  b2;
    input  a;
    assign z = ~(( c1 | c2 ) & ( a ) & (b1|b2));
endmodule
module bw_u1_oai221_8x (
    z,
    c1,
    c2,
    b1,
    b2,
    a );
    output z;
    input  c1;
    input  c2;
    input  b1;
    input  b2;
    input  a;
    assign z = ~(( c1 | c2 ) & ( a ) & (b1|b2));
endmodule
module bw_u1_oai222_1x (
    z,
    c1,
    c2,
    b1,
    b2,
    a1,
    a2 );
    output z;
    input  c1;
    input  c2;
    input  b1;
    input  b2;
    input  a1;
    input  a2;
    assign z = ~(( c1 | c2 ) & ( a1|a2 ) & (b1|b2));
endmodule
module bw_u1_oai222_2x (
    z,
    c1,
    c2,
    b1,
    b2,
    a1,
    a2 );
    output z;
    input  c1;
    input  c2;
    input  b1;
    input  b2;
    input  a1;
    input  a2;
    assign z = ~(( c1 | c2 ) & ( a1|a2 ) & (b1|b2));
endmodule
module bw_u1_oai222_4x (
    z,
    c1,
    c2,
    b1,
    b2,
    a1,
    a2 );
    output z;
    input  c1;
    input  c2;
    input  b1;
    input  b2;
    input  a1;
    input  a2;
    assign z = ~(( c1 | c2 ) & ( a1|a2 ) & (b1|b2));
endmodule
module bw_u1_oai311_1x (
    z,
    c1,
    c2,
    c3,
    b,
    a );
    output z;
    input  c1;
    input  c2;
    input  c3;
    input  b;
    input  a;
    assign z = ~(( c1 | c2|c3 ) & ( a ) & (b));
endmodule
module bw_u1_oai311_2x (
    z,
    c1,
    c2,
    c3,
    b,
    a );
    output z;
    input  c1;
    input  c2;
    input  c3;
    input  b;
    input  a;
    assign z = ~(( c1 | c2|c3 ) & ( a ) & (b));
endmodule
module bw_u1_oai311_4x (
    z,
    c1,
    c2,
    c3,
    b,
    a );
    output z;
    input  c1;
    input  c2;
    input  c3;
    input  b;
    input  a;
    assign z = ~(( c1 | c2 | c3 ) & ( a ) & (b));
endmodule
module bw_u1_oai311_8x (
    z,
    c1,
    c2,
    c3,
    b,
    a );
    output z;
    input  c1;
    input  c2;
    input  c3;
    input  b;
    input  a;
    assign z = ~(( c1 | c2|c3 ) & ( a ) & (b));
endmodule
module bw_u1_muxi21_0p6x (z, d0, d1, s);
output z;
input  d0, d1, s;
    assign z = s ? ~d1 : ~d0;
endmodule
module bw_u1_muxi21_1x (z, d0, d1, s);
output z;
input  d0, d1, s;
    assign z = s ? ~d1 : ~d0;
endmodule
module bw_u1_muxi21_2x (z, d0, d1, s);
output z;
input  d0, d1, s;
    assign z = s ? ~d1 : ~d0;
endmodule
module bw_u1_muxi21_4x (z, d0, d1, s);
output z;
input  d0, d1, s;
    assign z = s ? ~d1 : ~d0;
endmodule
module bw_u1_muxi21_6x (z, d0, d1, s);
output z;
input  d0, d1, s;
    assign z = s ? ~d1 : ~d0;
endmodule
module bw_u1_muxi31d_4x (z, d0, d1, d2, s0, s1, s2);
output z;
input  d0, d1, d2, s0, s1, s2;
        zmuxi31d_prim i0 ( z, d0, d1, d2, s0, s1, s2 );
endmodule
module bw_u1_muxi41d_4x (z, d0, d1, d2, d3, s0, s1, s2, s3);
output z;
input  d0, d1, d2, d3, s0, s1, s2, s3;
        zmuxi41d_prim i0 ( z, d0, d1, d2, d3, s0, s1, s2, s3 );
endmodule
module bw_u1_muxi41d_6x (z, d0, d1, d2, d3, s0, s1, s2, s3);
output z;
input  d0, d1, d2, d3, s0, s1, s2, s3;
        zmuxi41d_prim i0 ( z, d0, d1, d2, d3, s0, s1, s2, s3 );
endmodule
 
module bw_u1_xor2_0p6x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ( a ^ b );
endmodule
module bw_u1_xor2_1x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ( a ^ b );
endmodule
module bw_u1_xor2_2x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ( a ^ b );
endmodule
module bw_u1_xor2_4x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ( a ^ b );
endmodule
module bw_u1_xnor2_0p6x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a ^ b );
endmodule
module bw_u1_xnor2_1x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a ^ b );
endmodule
module bw_u1_xnor2_2x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a ^ b );
endmodule
module bw_u1_xnor2_4x (
    z,
    a,
    b );
    output z;
    input  a;
    input  b;
    assign z = ~( a ^ b );
endmodule
module bw_u1_buf_1x (
    z,
    a );
    output z;
    input  a;
    assign z = ( a );
endmodule
module bw_u1_buf_5x (
    z,
    a );
    output z;
    input  a;
    assign z = ( a );
endmodule
module bw_u1_buf_10x (
    z,
    a );
    output z;
    input  a;
    assign z = ( a );
endmodule
module bw_u1_buf_15x (
    z,
    a );
    output z;
    input  a;
    assign z = ( a );
endmodule
module bw_u1_buf_20x (
    z,
    a );
    output z;
    input  a;
    assign z = ( a );
endmodule
module bw_u1_buf_30x (
    z,
    a );
    output z;
    input  a;
    assign z = ( a );
endmodule
module bw_u1_buf_40x (
    z,
    a );
    output z;
    input  a;
    assign z = ( a );
endmodule
module bw_u1_ao2222_1x (
    z,
    a1,
    a2,
    b1,
    b2,
    c1,
    c2,
    d1,
    d2 );
    output z;
    input  a1;
    input  a2;
    input  b1;
    input  b2;
    input  c1;
    input  c2;
    input  d1;
    input  d2;
    assign z = ((d1&d2) | ( c1 & c2 ) | (b1&b2)| (a1& a2));
endmodule
module bw_u1_ao2222_2x (
    z,
    a1,
    a2,
    b1,
    b2,
    c1,
    c2,
    d1,
    d2 );
    output z;
    input  a1;
    input  a2;
    input  b1;
    input  b2;
    input  c1;
    input  c2;
    input  d1;
    input  d2;
    assign z = ((d1&d2) | ( c1 & c2 ) | (b1&b2)| (a1& a2));
endmodule
module bw_u1_ao2222_4x (
    z,
    a1,
    a2,
    b1,
    b2,
    c1,
    c2,
    d1,
    d2 );
    output z;
    input  a1;
    input  a2;
    input  b1;
    input  b2;
    input  c1;
    input  c2;
    input  d1;
    input  d2;
    assign z = ((d1&d2) | ( c1 & c2 ) | (b1&b2)| (a1& a2));
endmodule
module bw_u1_soff_1x (q, so, ck, d, se, sd);
output q, so;
input  ck, d, se, sd;
        zsoff_prim i0 ( q, so, ck, d, se, sd );
endmodule
module bw_u1_soff_2x (q, so, ck, d, se, sd);
output q, so;
input  ck, d, se, sd;
        zsoff_prim i0 ( q, so, ck, d, se, sd );
endmodule
module bw_u1_soff_4x (q, so, ck, d, se, sd);
output q, so;
input  ck, d, se, sd;
        zsoff_prim i0 ( q, so, ck, d, se, sd );
endmodule
module bw_u1_soff_8x (q, so, ck, d, se, sd);
output q, so;
input  ck, d, se, sd;
        zsoff_prim i0 ( q, so, ck, d, se, sd );
endmodule
module bw_u1_soffi_4x (q_l, so, ck, d, se, sd);
output q_l, so;
input  ck, d, se, sd;
        zsoffi_prim i0 ( q_l, so, ck, d, se, sd );
endmodule
  
module bw_u1_soffi_8x (q_l, so, ck, d, se, sd);
output q_l, so;
input  ck, d, se, sd;
        zsoffi_prim i0 ( q_l, so, ck, d, se, sd );
endmodule
module bw_u1_soffm2_4x (q, so, ck, d0, d1, s, se, sd);
output q, so;
input  ck, d0, d1, s, se, sd;
        zsoffm2_prim i0 ( q, so, ck, d0, d1, s, se, sd );
endmodule
module bw_u1_soffm2_8x (q, so, ck, d0, d1, s, se, sd);
output q, so;
input  ck, d0, d1, s, se, sd;
        zsoffm2_prim i0 ( q, so, ck, d0, d1, s, se, sd );
endmodule
module bw_u1_soffr_2x (q, so, ck, d, se, sd, r_l);
output q, so;
input  ck, d, se, sd, r_l;
        zsoffr_prim i0 ( q, so, ck, d, se, sd, r_l );
endmodule
  
module bw_u1_soffr_4x (q, so, ck, d, se, sd, r_l);
output q, so;
input  ck, d, se, sd, r_l;
        zsoffr_prim i0 ( q, so, ck, d, se, sd, r_l );
endmodule
module bw_u1_soffr_8x (q, so, ck, d, se, sd, r_l);
output q, so;
input  ck, d, se, sd, r_l;
        zsoffr_prim i0 ( q, so, ck, d, se, sd, r_l );
endmodule
module bw_u1_soffasr_2x (q, so, ck, d, r_l, s_l, se, sd);
output q, so;
input  ck, d, r_l, s_l, se, sd;
        zsoffasr_prim i0 (q, so, ck, d, r_l, s_l, se, sd);
endmodule
module bw_u1_ckbuf_1p5x  (clk, rclk);
output clk;
input  rclk;
        buf (clk, rclk);
endmodule
module bw_u1_ckbuf_3x  (clk, rclk);
output clk;
input  rclk;
        buf (clk, rclk);
endmodule
module bw_u1_ckbuf_4p5x  (clk, rclk);
output clk;
input  rclk;
        buf (clk, rclk);
endmodule
module bw_u1_ckbuf_6x  (clk, rclk);
output clk;
input  rclk;
        buf (clk, rclk);
endmodule
module bw_u1_ckbuf_7x  (clk, rclk);
output clk;
input  rclk;
        buf (clk, rclk);
endmodule
module bw_u1_ckbuf_8x  (clk, rclk);
output clk;
input  rclk;
        buf (clk, rclk);
endmodule
module bw_u1_ckbuf_11x (clk, rclk);
output clk;
input  rclk;
    assign clk = ( rclk );
endmodule
module bw_u1_ckbuf_14x (clk, rclk);
output clk;
input  rclk;
    assign clk = ( rclk );
endmodule
module bw_u1_ckbuf_17x (clk, rclk);
output clk;
input  rclk;
    assign clk = ( rclk );
endmodule
module bw_u1_ckbuf_19x (clk, rclk);
output clk;
input  rclk;
    assign clk = ( rclk );
endmodule
module bw_u1_ckbuf_22x (clk, rclk);
output clk;
input  rclk;
    assign clk = ( rclk );
endmodule
module bw_u1_ckbuf_25x (clk, rclk);
output clk;
input  rclk;
    assign clk = ( rclk );
endmodule
module bw_u1_ckbuf_28x (clk, rclk);
output clk;
input  rclk;
    assign clk = ( rclk );
endmodule
module bw_u1_ckbuf_30x (clk, rclk);
output clk;
input  rclk;
    assign clk = ( rclk );
endmodule
module bw_u1_ckbuf_33x (clk, rclk);
output clk;
input  rclk;
    assign clk = ( rclk );
endmodule
module bw_u1_ckbuf_40x (clk, rclk);
output clk;
input  rclk;
    assign clk = ( rclk );
endmodule
module bw_u1_ckenbuf_6x  (clk, rclk, en_l, tm_l);
output clk;
input  rclk, en_l, tm_l;
        zckenbuf_prim i0 ( clk, rclk, en_l, tm_l );
endmodule 
module bw_u1_ckenbuf_14x (clk, rclk, en_l, tm_l);
output clk;
input  rclk, en_l, tm_l;
        zckenbuf_prim i0 ( clk, rclk, en_l, tm_l );
endmodule   
module bw_u1_zhinv_0p6x (z, a);
output z;
input  a;
        not (z, a);
endmodule
module bw_u1_zhinv_1x (z, a);
output z;
input  a;
        not (z, a);
endmodule
module bw_u1_zhinv_1p4x (z, a);
output z;
input  a;
        not (z, a);
endmodule
module bw_u1_zhinv_2x (z, a);
output z;
input  a;
        not (z, a);
endmodule
module bw_u1_zhinv_3x (z, a);
output z;
input  a;
        not (z, a);
endmodule
module bw_u1_zhinv_4x (z, a);
output z;
input  a;
        not (z, a);
endmodule
module bw_u1_zhnand2_0p4x (z, a, b);
output z;
input  a, b;
        nand (z, a, b);
endmodule
module bw_u1_zhnand2_0p6x (z, a, b);
output z;   
input  a, b;
        nand (z, a, b);
endmodule   
module bw_u1_zhnand2_1x (z, a, b);
output z;   
input  a, b;
        nand (z, a, b);
endmodule   
module bw_u1_zhnand2_1p4x (z, a, b);
output z;   
input  a, b;
        nand (z, a, b);
endmodule   
module bw_u1_zhnand2_2x (z, a, b);
output z;   
input  a, b;
        nand (z, a, b);
endmodule   
module bw_u1_zhnand2_3x (z, a, b);
output z;   
input  a, b;
        nand (z, a, b);
endmodule   
module bw_u1_zhnand3_0p6x (z, a, b, c);
output z;
input  a, b, c;
        nand (z, a, b, c);
endmodule
module bw_u1_zhnand3_1x (z, a, b, c);
output z;
input  a, b, c;
        nand (z, a, b, c);
endmodule
module bw_u1_zhnand3_2x (z, a, b, c);
output z;
input  a, b, c;
        nand (z, a, b, c);
endmodule
module bw_u1_zhnand4_0p6x (z, a, b, c, d);
output z;
input  a, b, c, d;
        nand (z, a, b, c, d);
endmodule
module bw_u1_zhnand4_1x (z, a, b, c, d);
output z;
input  a, b, c, d;
        nand (z, a, b, c, d);
endmodule
module bw_u1_zhnand4_2x (z, a, b, c, d);
output z;
input  a, b, c, d;
        nand (z, a, b, c, d);
endmodule
        
module bw_u1_zhnor2_0p6x (z, a, b);
output z;
input  a, b;
        nor (z, a, b);
endmodule
module bw_u1_zhnor2_1x (z, a, b);
output z;   
input  a, b;
        nor (z, a, b);
endmodule
module bw_u1_zhnor2_2x (z, a, b);
output z;   
input  a, b;
        nor (z, a, b);
endmodule
module bw_u1_zhnor3_0p6x (z, a, b, c);
output z;
input  a, b, c;
        nor (z, a, b, c);
endmodule
module bw_u1_zhaoi21_0p4x (z,b1,b2,a);
    output z;   
    input  b1;
    input  b2;
    input  a;
    assign z = ~(( b1 & b2 ) | ( a ));
    
endmodule
module bw_u1_zhaoi21_1x (z, a, b1, b2);
    output z;
    input  b1;
    input  b2;
    input  a;
    assign z = ~(( b1 & b2 ) | ( a ));
endmodule
module bw_u1_zhoai21_1x (z,b1,b2,a );
    
    output z;
    input  b1;
    input  b2;  
    input  a;
  
    assign z = ~(( b1 | b2 ) & ( a ));
      
endmodule
module bw_u1_zhoai211_0p3x (z, a, b, c1, c2);
    output z; 
    input  c1;  
    input  c2;
    input  b;
    input  a;
      
    assign z = ~(( c1 | c2 ) & ( a ) & (b));
       
endmodule
module bw_u1_zhoai211_1x (z, a, b, c1, c2);
output z;
input  a, b, c1, c2;
    assign z = ~(( c1 | c2 ) & ( a ) & (b));
       
endmodule
module bw_u1_scanlg_2x (so, sd, ck, se);
output so;
input sd, ck, se;
reg so_l;
    assign so = ~so_l;
    always @ ( ck or sd or se )
       if (~ck) so_l <= ~(sd & se) ;
endmodule
module bw_u1_scanl_2x (so, sd, ck);
output so;
input sd, ck;
reg so_l;
    assign so = ~so_l;
    always @ ( ck or sd )
       if (~ck) so_l <= ~sd ;
endmodule
module bw_u1_syncff_4x (q, so, ck, d, se, sd);
output q, so;
input  ck, d, se, sd;
reg    q_r;
  always @ (posedge ck)
      q_r <= se ? sd : d;
  assign q  = q_r;
  assign so = q_r;
endmodule
module bw_u1_zzeccxor2_5x (z, a, b); 
 output z; 
 input a, b;
    assign z = ( a ^ b );
endmodule
module bw_u1_zzmulcsa42_5x (sum, carry, cout, a, b, c, d, cin);
output sum, carry, cout;
input  a, b, c, d, cin;
wire and_cin_b, or_cin_b, xor_a_c_d, and_or_cin_b_xor_a_c_d;
wire and_a_c, and_a_d, and_c_d;
        assign sum   = cin ^ a ^ b ^ c ^ d;
        assign carry = cin & b | (cin | b) & (a ^ c ^ d);
        assign cout  = a & c | a & d | c & d;
endmodule
module bw_u1_zzmulcsa32_5x (sum, cout, a, b, c);
output sum, cout;
input  a, b, c;
wire and_a_b, and_a_c, and_b_c;
        assign sum  = a ^ b ^ c ;
        assign cout = a & b | a & c | b & c ;
endmodule
module bw_u1_zzmulppmuxi21_2x ( z, d0, d1, s );
output  z;
input  d0, d1, s;
    assign z = s ? ~d1 : ~d0;
endmodule
module bw_u1_zzmulnand2_2x ( z, a, b );
output z;
input  a;
input  b;
    assign z = ~( a & b );
endmodule
module zmuxi31d_prim (z, d0, d1, d2, s0, s1, s2);
output z;
input  d0, d1, d2, s0, s1, s2;
wire [2:0] sel = {s0,s1,s2}; 
reg z;
    always @ (s2 or d2 or s1 or d1 or s0 or d0)
        casez ({s2,d2,s1,d1,s0,d0})
            6'b0?0?10: z = 1'b1;  
            6'b0?0?11: z = 1'b0;  
            6'b0?100?: z = 1'b1;  
            6'b0?110?: z = 1'b0;  
            6'b0?1010: z = 1'b1;  
            6'b0?1111: z = 1'b0;  
            6'b100?0?: z = 1'b1;  
            6'b110?0?: z = 1'b0;  
            6'b100?10: z = 1'b1;  
            6'b110?11: z = 1'b0;  
            6'b10100?: z = 1'b1;  
            6'b11110?: z = 1'b0;  
            6'b101010: z = 1'b1;  
            6'b111111: z = 1'b0;  
            default: z = 1'bx;
        endcase
endmodule
module zmuxi41d_prim (z, d0, d1, d2, d3, s0, s1, s2, s3);
output z;
input  d0, d1, d2, d3, s0, s1, s2, s3;
wire [3:0] sel = {s0,s1,s2,s3}; 
reg z;
    always @ (s3 or d3 or s2 or d2 or s1 or d1 or s0 or d0)
        casez ({s3,d3,s2,d2,s1,d1,s0,d0})
            8'b0?0?0?10: z = 1'b1;
            8'b0?0?0?11: z = 1'b0;
            8'b0?0?100?: z = 1'b1;
            8'b0?0?110?: z = 1'b0;
            8'b0?0?1010: z = 1'b1;
            8'b0?0?1111: z = 1'b0;
            8'b0?100?0?: z = 1'b1;
            8'b0?110?0?: z = 1'b0;
            8'b0?100?10: z = 1'b1;
            8'b0?110?11: z = 1'b0;
            8'b0?10100?: z = 1'b1;
            8'b0?11110?: z = 1'b0;
            8'b0?101010: z = 1'b1;
            8'b0?111111: z = 1'b0;
            8'b100?0?0?: z = 1'b1;
            8'b110?0?0?: z = 1'b0;
            8'b100?0?10: z = 1'b1;
            8'b110?0?11: z = 1'b0;
            8'b100?100?: z = 1'b1;
            8'b110?110?: z = 1'b0;
            8'b100?1010: z = 1'b1;
            8'b110?1111: z = 1'b0;
            8'b10100?0?: z = 1'b1;
            8'b11110?0?: z = 1'b0;
            8'b10100?10: z = 1'b1;
            8'b11110?11: z = 1'b0;
            8'b1010100?: z = 1'b1;
            8'b1111110?: z = 1'b0;
            8'b10101010: z = 1'b1;
            8'b11111111: z = 1'b0;
            default: z = 1'bx;
        endcase   
endmodule
module zsoff_prim (q, so, ck, d, se, sd);
output q, so;
input  ck, d, se, sd;
reg    q_r;
  always @ (posedge ck)
      q_r <= se ? sd : d;
  assign q  = q_r;
  assign so = q_r ;
endmodule
module zsoffr_prim (q, so, ck, d, se, sd, r_l);
output q, so;
input  ck, d, se, sd, r_l;
reg    q_r;
  always @ (posedge ck)
      q_r <= se ? sd : (d & r_l) ;
  assign q  = q_r;
  assign so = q_r;
endmodule
module zsoffi_prim (q_l, so, ck, d, se, sd);
output q_l, so;
input  ck, d, se, sd;
reg    q_r;
  always @ (posedge ck)
      q_r <= se ? sd : d;
  assign q_l = ~q_r;
  assign so  = q_r;
endmodule
module zsoffm2_prim (q, so, ck, d0, d1, s, se, sd);
output q, so;
input  ck, d0, d1, s, se, sd;
reg    q_r;
  always @ (posedge ck)
      q_r <= se ? sd : (s ? d1 : d0) ;
  assign q  = q_r;
  assign so = q_r;
endmodule
module zsoffasr_prim (q, so, ck, d, r_l, s_l, se, sd);
  output q, so;
  input ck, d, r_l, s_l, se, sd;
  
  
  reg q;
  wire so;
  always @ (posedge ck or negedge r_l or negedge s_l) begin
		if(~r_l) q <= 1'b0;
		else if (~s_l) q <= r_l;
		else if (se) q <= r_l & s_l & sd;
		else q <= r_l & s_l & (~se) & d;
  end
  assign so = q | ~se;
endmodule
module zckenbuf_prim (clk, rclk, en_l, tm_l);
output clk;
input  rclk, en_l, tm_l;
reg    clken;
  always @ (rclk or en_l or tm_l)
    if (!rclk)  
      clken <= ~en_l | ~tm_l;
  assign clk = clken & rclk;
endmodule
module bw_mckbuf_40x (clk, rclk, en);
output clk;
input  rclk;
input  en;
    assign clk = rclk & en ;
endmodule
module bw_mckbuf_33x (clk, rclk, en);
output clk;
input  rclk;
input  en;
    assign clk = rclk & en ;
endmodule
module bw_mckbuf_30x (clk, rclk, en);
output clk;
input  rclk;
input  en;
    assign clk = rclk & en ;
endmodule
module bw_mckbuf_28x (clk, rclk, en);
output clk;
input  rclk;
input  en;
    assign clk = rclk & en ;
endmodule
module bw_mckbuf_25x (clk, rclk, en);
output clk;
input  rclk;
input  en;
    assign clk = rclk & en ;
endmodule
module bw_mckbuf_22x (clk, rclk, en);
output clk;
input  rclk;
input  en;
    assign clk = rclk & en ;
endmodule
module bw_mckbuf_19x (clk, rclk, en);
output clk;
input  rclk;
input  en;
    assign clk = rclk & en ;
endmodule
module bw_mckbuf_17x (clk, rclk, en);
output clk;
input  rclk;
input  en;
    assign clk = rclk & en ;
endmodule
module bw_mckbuf_14x (clk, rclk, en);
output clk;
input  rclk;
input  en;
    assign clk = rclk & en ;
endmodule
module bw_mckbuf_11x (clk, rclk, en);
output clk;
input  rclk;
input  en;
    assign clk = rclk & en ;
endmodule
module bw_mckbuf_8x (clk, rclk, en);
output clk;
input  rclk;
input  en;
    assign clk = rclk & en ;
endmodule
module bw_mckbuf_7x (clk, rclk, en);
output clk;
input  rclk;
input  en;
    assign clk = rclk & en ;
endmodule
module bw_mckbuf_6x (clk, rclk, en);
output clk;
input  rclk;
input  en;
    assign clk = rclk & en ;
endmodule
module bw_mckbuf_4p5x (clk, rclk, en);
output clk;
input  rclk;
input  en;
    assign clk = rclk & en ;
endmodule
module bw_mckbuf_3x (clk, rclk, en);
output clk;
input  rclk;
input  en;
    assign clk = rclk & en ;
endmodule
module bw_mckbuf_1p5x (clk, rclk, en);
output clk;
input  rclk;
input  en;
    assign clk = rclk & en ;
endmodule
module bw_u1_minbuf_1x (
    z,
    a );
    output z;
    input  a;
    assign z = ( a );
endmodule
module bw_u1_minbuf_4x (
    z,
    a );
    output z;
    input  a;
    assign z = ( a );
endmodule
module bw_u1_minbuf_5x (
    z,
    a );
    output z;
    input  a;
    assign z = ( a );
endmodule
module bw_u1_ckenbuf_4p5x  (clk, rclk, en_l, tm_l);
output clk;
input  rclk, en_l, tm_l;
        zckenbuf_prim i0 ( clk, rclk, en_l, tm_l );
endmodule 
module bw_u1_fill_1x(\vdd! );
input \vdd! ;
endmodule
module bw_u1_fill_2x(\vdd! );
input \vdd! ;
endmodule
module bw_u1_fill_3x(\vdd! );
input \vdd! ;
endmodule
module bw_u1_fill_4x(\vdd! );
input \vdd! ;
endmodule
  
    
    
    
    
    
    
    
        
        
        
        
        
        
        
        
        
        
        
 
        
        
        
        
 
			
module ucb_bus_in (
   
   stall, indata_buf_vld, indata_buf,
   
   rst_l, clk, vld, data, stall_a1
   );
   
   parameter UCB_BUS_WIDTH = 32;
   parameter REG_WIDTH = 64;
   
   input                     rst_l;
   input 		     clk;
   
   input 		     vld;
   input [UCB_BUS_WIDTH-1:0] data;
   output 		     stall;
   
   output 		     indata_buf_vld;
   output [REG_WIDTH+63:0]   indata_buf;
   input 		     stall_a1; 
   
   wire 		     vld_d1;
   wire 		     stall_d1;
   wire [UCB_BUS_WIDTH-1:0]  data_d1;
   wire 		     skid_buf0_en;
   wire 		     vld_buf0;
   wire [UCB_BUS_WIDTH-1:0]  data_buf0;
   wire 		     skid_buf1_en;
   wire 		     vld_buf1;
   wire [UCB_BUS_WIDTH-1:0]  data_buf1;
   wire 		     skid_buf0_sel;
   wire 		     skid_buf1_sel;
   wire 		     vld_mux;
   wire [UCB_BUS_WIDTH-1:0]  data_mux;
   wire [(REG_WIDTH+64)/UCB_BUS_WIDTH-1:0] indata_vec_next;
   wire [(REG_WIDTH+64)/UCB_BUS_WIDTH-1:0] indata_vec;
   wire [REG_WIDTH+63:0]     indata_buf_next;
   wire 		     indata_vec0_d1;
   
   dffrle_ns #(1) vld_d1_ff (.din(vld),
			     .rst_l(rst_l),
			     .en(~stall_d1),
			     .clk(clk),
			     .q(vld_d1));
   dffe_ns #(UCB_BUS_WIDTH) data_d1_ff (.din(data),
					.en(~stall_d1),
					.clk(clk),
					.q(data_d1));
   dffrl_ns #(1) stall_ff (.din(stall_a1),
			   .clk(clk),
			   .rst_l(rst_l),
			   .q(stall));
   dffrl_ns #(1) stall_d1_ff (.din(stall),
			      .clk(clk),
			      .rst_l(rst_l),
			      .q(stall_d1));
   
   
   
   
   
   
   assign 	 skid_buf0_en = stall_a1 & ~stall;
   dffrle_ns #(1) vld_buf0_ff (.din(vld_d1),
			       .rst_l(rst_l),
			       .en(skid_buf0_en),
			       .clk(clk),
			       .q(vld_buf0));
   dffe_ns #(UCB_BUS_WIDTH) data_buf0_ff (.din(data_d1),
					  .en(skid_buf0_en),
					  .clk(clk),
					  .q(data_buf0));
   
   dffrl_ns #(1) skid_buf1_en_ff (.din(skid_buf0_en),
				  .clk(clk),
				  .rst_l(rst_l),
				  .q(skid_buf1_en));
   dffrle_ns #(1) vld_buf1_ff (.din(vld_d1),
			       .rst_l(rst_l),
			       .en(skid_buf1_en),
			       .clk(clk),
			       .q(vld_buf1));
   dffe_ns #(UCB_BUS_WIDTH) data_buf1_ff (.din(data_d1),
					  .en(skid_buf1_en),
					  .clk(clk),
					  .q(data_buf1));
   
   
   
   
   
   assign 	 skid_buf0_sel = ~stall_a1 & stall;
   dffrl_ns #(1) skid_buf1_sel_ff (.din(skid_buf0_sel),
				   .clk(clk),
				   .rst_l(rst_l),
				   .q(skid_buf1_sel));
   assign 	 vld_mux = skid_buf0_sel ? vld_buf0 :
		           skid_buf1_sel ? vld_buf1 :
		                           vld_d1;
   assign 	 data_mux = skid_buf0_sel ? data_buf0 :
		            skid_buf1_sel ? data_buf1 :
		                            data_d1;
   
   
   assign 	 indata_vec_next = {vld_mux,
				    indata_vec[(REG_WIDTH+64)/UCB_BUS_WIDTH-1:1]};
   dffrle_ns #((REG_WIDTH+64)/UCB_BUS_WIDTH) indata_vec_ff (.din(indata_vec_next),
							    .en(~stall_a1),
							    .rst_l(rst_l),
							    .clk(clk),
							    .q(indata_vec));
   
   assign 	 indata_buf_next = {data_mux,
				    indata_buf[REG_WIDTH+63:UCB_BUS_WIDTH]};
   dffe_ns #(REG_WIDTH+64) indata_buf_ff (.din(indata_buf_next),
					  .en(~stall_a1),
					  .clk(clk),
					  .q(indata_buf));
   
   dffrle_ns #(1) indata_vec0_d1_ff (.din(indata_vec[0]),
				     .rst_l(rst_l),
				     .en(~stall_a1),
				     .clk(clk),
				     .q(indata_vec0_d1));
   assign        indata_buf_vld = indata_vec[0] & ~indata_vec0_d1;
endmodule 
  
    
    
    
    
    
    
    
        
        
        
        
        
        
        
        
        
        
        
 
        
        
        
        
 
                        
module ucb_bus_out (
   
   vld, data, outdata_buf_busy,
   
   clk, rst_l, stall, outdata_buf_in, outdata_vec_in, outdata_buf_wr
   );
   
   parameter UCB_BUS_WIDTH = 32;
   parameter REG_WIDTH = 64;            
                                        
   
   input                                clk;
   input 				rst_l;
   
   output 				vld;
   output [UCB_BUS_WIDTH-1:0] 		data;
   input 				stall;
   
   output 				outdata_buf_busy;  
   input [REG_WIDTH+63:0] 		outdata_buf_in;
   input [(REG_WIDTH+64)/UCB_BUS_WIDTH-1:0] outdata_vec_in; 
   input 				outdata_buf_wr;
   
   wire 				stall_d1;
   wire [(REG_WIDTH+64)/UCB_BUS_WIDTH-1:0] 	outdata_vec;
   wire [(REG_WIDTH+64)/UCB_BUS_WIDTH-1:0] 	outdata_vec_next;
   wire [REG_WIDTH+63:0] 		outdata_buf;
   reg [REG_WIDTH+63:0] 		outdata_buf_next;
   wire 				load_outdata;
   wire 				shift_outdata;
   
   assign 	 vld = outdata_vec[0];
   
   assign    data = outdata_buf[UCB_BUS_WIDTH-1:0];
   dffrl_ns #(1) stall_d1_ff (.din(stall),
                              .clk(clk),
                              .rst_l(rst_l),
                              .q(stall_d1));
   
   
   assign 	 load_outdata = outdata_buf_wr & ~outdata_buf_busy;
   assign 	 outdata_buf_busy = outdata_vec[0] | stall_d1;
   
   assign 	 shift_outdata = outdata_vec[0] & ~stall_d1;
   assign 	 outdata_vec_next =
		 load_outdata  ? outdata_vec_in:
		 shift_outdata ? outdata_vec >> 1:
	                         outdata_vec;
   dffrl_ns #((REG_WIDTH+64)/UCB_BUS_WIDTH) outdata_vec_ff (.din(outdata_vec_next),
							    .clk(clk),
							    .rst_l(rst_l),
							    .q(outdata_vec));
   
		 
		 
	  
   always @ *
   begin
      if (load_outdata)
         outdata_buf_next = outdata_buf_in;
      else if (shift_outdata)
      begin
         outdata_buf_next = outdata_buf >> UCB_BUS_WIDTH;
         if (outdata_vec[1] == 1'b0)
            outdata_buf_next[UCB_BUS_WIDTH-1:0] = 0;
      end
      else
         outdata_buf_next = outdata_buf; 
   end
   dff_ns #(REG_WIDTH+64) outdata_buf_ff (.din(outdata_buf_next),
					  .clk(clk),
					  .q(outdata_buf));
endmodule 
module valrdy_to_credit (
            clk,
            reset,
                
            
            data_in,
            valid_in,
            ready_in,
			
            data_out,
            valid_out,
		    yummy_out);
parameter BUFFER_SIZE = 4;
parameter BUFFER_BITS = 3;
   
input clk;
input reset;
 
input [64-1:0]	 data_in;
 input valid_in;			
 input yummy_out;			
output [64-1:0]  data_out;
 output valid_out;
 output ready_in;		
 reg yummy_out_f;
 reg valid_temp_f;
 reg [BUFFER_BITS-1:0] count_f;
reg is_one_f;
 reg is_two_or_more_f;
 wire [BUFFER_BITS-1:0] count_plus_1;
 wire [BUFFER_BITS-1:0] count_minus_1;
 wire up;
 wire down;
 wire valid_temp;
  reg [BUFFER_BITS-1:0] count_temp;
assign data_out = data_in;
assign valid_temp = valid_in & ready_in;
assign valid_out = valid_temp;
assign count_plus_1 = count_f + 1'b1;
assign count_minus_1 = count_f - 1'b1;
assign ready_in = is_two_or_more_f;
assign up = yummy_out_f & ~valid_temp_f;
assign down = ~yummy_out_f & valid_temp_f;
always @ (count_f or count_plus_1 or count_minus_1 or up or down)
begin
	case (count_f)
	0:
		begin
			if(up)
			begin
				count_temp <= count_plus_1;
			end
			else
			begin
				count_temp <= count_f;
			end
		end
	BUFFER_SIZE:
		begin
			if(down)
			begin
				count_temp <= count_minus_1;
			end
			else
			begin
				count_temp <= count_f;
			end
		end
	default:
		begin
			case ({up, down})
				2'b10:	count_temp <= count_plus_1;
				2'b01:	count_temp <= count_minus_1;
				default:	count_temp <= count_f;
			endcase
		end
	endcase
end
 wire top_bits_zero_temp = count_temp < 3 ? 1 : 0;
always @ (posedge clk)
begin
	if(reset)
	begin
	   count_f <= BUFFER_SIZE;
	   yummy_out_f <= 1'b0;
	   valid_temp_f <= 1'b0;
	   is_one_f <= (BUFFER_SIZE == 1);
	   is_two_or_more_f <= (BUFFER_SIZE >= 2);
	end
	else
	begin
	   count_f <= count_temp;
	   yummy_out_f <= yummy_out;
	   valid_temp_f <= valid_temp;
	   is_one_f         <= top_bits_zero_temp & count_temp[0];
   	   is_two_or_more_f <= ~top_bits_zero_temp;
	end
end
endmodule
      
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
module flat_id_to_xy(
    input  [(6-1):0] flat_id,
    output reg [(8-1):0] x_coord,
    output reg [(8-1):0] y_coord
);
    always @*
    begin
        case (flat_id)
        
6'd0: 
begin
    x_coord = 8'd0;
    y_coord = 8'd0;
end
        default:
        begin
            x_coord = 8'dX;
            y_coord = 8'dX;
        end
        endcase
    end
endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
module xy_to_flat_id(
    input  [(8-1):0] x_coord,
    input  [(8-1):0] y_coord,
    output reg [(6-1):0] flat_id
);
    
    
    always @*
    begin
        case (x_coord)
        
8'd0:
begin
     case (y_coord)
    
    8'd0:
    begin
        flat_id = 6'd0;
    end
     default:
     begin
         flat_id = 6'dX;
     end
     endcase
end
        default:
        begin
            flat_id = 6'dX;
        end
        endcase
    end
endmodule
module sync_fifo 
#(
	parameter DSIZE = 64,
	parameter ASIZE = 5,
	parameter MEMSIZE = 16 
)
(
	rdata, 
	empty,
	clk,
	ren,
	wdata,
	full,
	wval,
	reset
	);
output reg [DSIZE-1:0] 	rdata;
output reg			empty;
output reg			full;
input	[DSIZE-1:0]	wdata;
input			wval;
input			ren;
input			clk;
input 			reset;
reg [DSIZE-1:0] sync_buf_mem_f [MEMSIZE-1:0];
reg [ASIZE:0] sync_buf_counter_f;
reg [ASIZE:0] sync_buf_counter_next;
reg [ASIZE-2:0] sync_rd_ptr_f;
reg [ASIZE-2:0] sync_rd_ptr_next;
reg [ASIZE-2:0] sync_wr_ptr_f;
reg [ASIZE-2:0] sync_wr_ptr_next;
always @ *
begin
    empty = (sync_buf_counter_f == 0);
    full =  (sync_buf_counter_f ==  MEMSIZE);
end
always @ *
begin
    if (reset)
    begin
        sync_buf_counter_next = 0;
    end
    else if ((wval && !full) && (ren && !empty))
    begin
        sync_buf_counter_next = sync_buf_counter_f;
    end
    else if (wval && !full)
    begin
        sync_buf_counter_next = sync_buf_counter_f + 1;
    end
    else if (ren && !empty)
    begin
        sync_buf_counter_next = sync_buf_counter_f - 1;
    end
    else
    begin
        sync_buf_counter_next = sync_buf_counter_f;
    end
end
always @ (posedge clk)
begin
    sync_buf_counter_f <= sync_buf_counter_next;
end
always @ *
begin
    if (reset)
    begin   
        sync_rd_ptr_next = 0;
    end
    else if (ren && !empty)
    begin
        sync_rd_ptr_next = sync_rd_ptr_f + 1;
    end
    else
    begin
        sync_rd_ptr_next = sync_rd_ptr_f;
    end
end
always @ (posedge clk)
begin
    sync_rd_ptr_f <= sync_rd_ptr_next;
end
always @ *
begin
    if (reset)
    begin   
        sync_wr_ptr_next = 0;
    end
    else if (wval && !full)
    begin
        sync_wr_ptr_next = sync_wr_ptr_f + 1;
    end
    else
    begin
        sync_wr_ptr_next = sync_wr_ptr_f;
    end
end
always @ (posedge clk)
begin
    sync_wr_ptr_f <= sync_wr_ptr_next;
end
always @ *
begin
    rdata = sync_buf_mem_f[sync_rd_ptr_f];
end
always @ (posedge clk)
begin
    if (wval && !full)
    begin
        sync_buf_mem_f[sync_wr_ptr_f] <= wdata;
    end
    else
    begin 
        sync_buf_mem_f[sync_wr_ptr_f] <= sync_buf_mem_f[sync_wr_ptr_f];
    end
end
endmodule
 
    
    
    
    
    
    
 
 
 
  
    
 
 
    
    
    
    
    
    
    
 
 
module chip_bridge_in (
    rst, 
    wr_clk,
    rd_clk,
    async_mux,
    bout_data_1,
    bout_val_1,
    bout_rdy_1,
    bout_data_2,
    bout_val_2,
    bout_rdy_2,
    bout_data_3,
    bout_val_3,
    bout_rdy_3,
    data_from_fpga,
    data_channel,
    credit_to_fpga
); 
input rst;
input wr_clk;
input rd_clk;
input async_mux;
input bout_rdy_1;
input bout_rdy_2;
input bout_rdy_3;
input [31:0] data_from_fpga;
input [ 1:0] data_channel;
output [63:0]   bout_data_1;
output          bout_val_1;
output [63:0]   bout_data_2;
output          bout_val_2;
output [63:0]   bout_data_3;
output          bout_val_3;
output [2:0]    credit_to_fpga;
wire [63:0] async_bout_data_1;
wire [63:0] async_bout_data_2;
wire [63:0] async_bout_data_3;
wire [63:0] sync_bout_data_1;
wire [63:0] sync_bout_data_2;
wire [63:0] sync_bout_data_3;
wire sort_rdy_1;
wire sort_rdy_2;
wire sort_rdy_3;
wire [63:0] sort_data_1;
wire [63:0] sort_data_2;
wire [63:0] sort_data_3;
wire sort_val_1;
wire sort_val_2;
wire sort_val_3;
wire fifo1_empty;
wire fifo2_empty;
wire fifo3_empty;
wire async_fifo1_empty;
wire async_fifo2_empty;
wire async_fifo3_empty;
wire sync_fifo1_empty;
wire sync_fifo2_empty;
wire sync_fifo3_empty;
wire fifo1_full;
wire fifo2_full;
wire fifo3_full;
wire credit_fifo_full;
wire async_fifo1_full;
wire async_fifo2_full;
wire async_fifo3_full;
wire async_credit_fifo_full;
wire sync_fifo1_full;
wire sync_fifo2_full;
wire sync_fifo3_full;
wire sync_credit_fifo_full;
assign bout_val_1 = ~fifo1_empty & ~credit_fifo_full;
assign bout_val_2 = ~fifo2_empty & ~credit_fifo_full;
assign bout_val_3 = ~fifo3_empty & ~credit_fifo_full;
reg [31:0] channel_buffer;
reg [0:0]  channel_buffer_count;
wire [63:0] buffered_data;
reg [1:0] buffered_channel;
assign sort_data_1 = (buffered_channel == 2'b01 && channel_buffer_count == 1'b1) ? buffered_data : 64'd0;
assign sort_data_2 = (buffered_channel == 2'b10 && channel_buffer_count == 1'b1) ? buffered_data : 64'd0;
assign sort_data_3 = (buffered_channel == 2'b11 && channel_buffer_count == 1'b1) ? buffered_data : 64'd0;
assign sort_val_1  = (buffered_channel == 2'b01 && channel_buffer_count == 1'b1) ? 1'b1 : 1'b0;
assign sort_val_2  = (buffered_channel == 2'b10 && channel_buffer_count == 1'b1) ? 1'b1 : 1'b0;
assign sort_val_3  = (buffered_channel == 2'b11 && channel_buffer_count == 1'b1) ? 1'b1 : 1'b0;
assign buffered_data = {data_from_fpga, channel_buffer};
always @(posedge wr_clk) begin
 
    if(rst) begin
        channel_buffer <= 32'd0;
        channel_buffer_count <= 0;
    end
    else begin
        if(data_channel != 0) begin 
            channel_buffer <= data_from_fpga;
            buffered_channel <= data_channel;
            channel_buffer_count <= channel_buffer_count + 1'b1;
        end
        else begin
            buffered_channel <= data_channel;
            channel_buffer_count <= 1'b0;
        end
    end
end
 
async_fifo #(
.DSIZE(64),
.ASIZE(5),
.MEMSIZE(16) )
async_fifo_1(
    .rreset(rst),
    .wreset(rst),
    .wclk(wr_clk),
    .rclk(rd_clk),
    .ren(bout_rdy_1 & ~credit_fifo_full & async_mux),
    .wval(sort_val_1 & async_mux),
    .wdata(sort_data_1),
    .rdata(async_bout_data_1),
    .wfull(async_fifo1_full), 
    .rempty(async_fifo1_empty)
);
 
 
async_fifo #(
.DSIZE(64),
.ASIZE(5),
.MEMSIZE(16) )
async_fifo_2(
    .rreset(rst),
    .wreset(rst),
    .wclk(wr_clk),
    .rclk(rd_clk),
    .ren(bout_rdy_2 & ~credit_fifo_full & async_mux),
    .wval(sort_val_2 & async_mux),
    .wdata(sort_data_2),
    .rdata(async_bout_data_2),
    .wfull(async_fifo2_full), 
    .rempty(async_fifo2_empty)
);
 
 
async_fifo #(
.DSIZE(64),
.ASIZE(5),
.MEMSIZE(16) )
async_fifo_3(
    .rreset(rst),
    .wreset(rst),
    .wclk(wr_clk),
    .rclk(rd_clk),
    .ren(bout_rdy_3 & ~credit_fifo_full & async_mux),
    .wval(sort_val_3 & async_mux),
    .wdata(sort_data_3),
    .rdata(async_bout_data_3),
    .wfull(async_fifo3_full), 
    .rempty(async_fifo3_empty)
);
 
 
sync_fifo #(
.DSIZE(64),
.ASIZE(5),
.MEMSIZE(16) )
sync_fifo_1(
    .reset(rst),
    .clk(wr_clk),
    .ren(bout_rdy_1 & ~credit_fifo_full & ~async_mux),
    .wval(sort_val_1 & ~async_mux),
    .wdata(sort_data_1),
    .rdata(sync_bout_data_1),
    .full(sync_fifo1_full), 
    .empty(sync_fifo1_empty)
);
 
 
sync_fifo #(
.DSIZE(64),
.ASIZE(5),
.MEMSIZE(16) )
sync_fifo_2(
    .reset(rst),
    .clk(wr_clk),
    .ren(bout_rdy_2 & ~credit_fifo_full & ~async_mux),
    .wval(sort_val_2 & ~async_mux),
    .wdata(sort_data_2),
    .rdata(sync_bout_data_2),
    .full(sync_fifo2_full), 
    .empty(sync_fifo2_empty)
);
 
 
sync_fifo #(
.DSIZE(64),
.ASIZE(5),
.MEMSIZE(16) )
sync_fifo_3(
    .reset(rst),
    .clk(wr_clk),
    .ren(bout_rdy_3 & ~credit_fifo_full & ~async_mux),
    .wval(sort_val_3 & ~async_mux),
    .wdata(sort_data_3),
    .rdata(sync_bout_data_3),
    .full(sync_fifo3_full), 
    .empty(sync_fifo3_empty)
);
 
assign fifo1_full = async_mux ? async_fifo1_full : sync_fifo1_full;
assign fifo2_full = async_mux ? async_fifo2_full : sync_fifo2_full;
assign fifo3_full = async_mux ? async_fifo3_full : sync_fifo3_full;
assign fifo1_empty = async_mux ? async_fifo1_empty : sync_fifo1_empty;
assign fifo2_empty = async_mux ? async_fifo2_empty : sync_fifo2_empty;
assign fifo3_empty = async_mux ? async_fifo3_empty : sync_fifo3_empty;
assign bout_data_1 = async_mux ? async_bout_data_1 : sync_bout_data_1;
assign bout_data_2 = async_mux ? async_bout_data_2 : sync_bout_data_2;
assign bout_data_3 = async_mux ? async_bout_data_3 : sync_bout_data_3;
wire [2:0] credit_gather;
wire credit_empty;
wire async_credit_empty;
wire sync_credit_empty;
wire [2:0] credit_fifo_out;
wire [2:0] async_credit_fifo_out;
wire [2:0] sync_credit_fifo_out;
reg  [2:0] credit_to_fpga_r ;
 
async_fifo #(
.DSIZE(3),
.ASIZE(5),
.MEMSIZE(16) )
async_credit_fifo(
    .rreset(rst),
    .wreset(rst),
    .wclk(rd_clk),
    .rclk(wr_clk),
    .ren(~rst & async_mux),
    .wval(~(rst) & (| credit_gather) & async_mux),
    .wdata(credit_gather),
    .rdata(async_credit_fifo_out),
    .wfull(async_credit_fifo_full),   
    .rempty(async_credit_empty)
);
 
 
sync_fifo #(
.DSIZE(3),
.ASIZE(5),
.MEMSIZE(16) )
sync_credit_fifo(
    .reset(rst),
    .clk(wr_clk),
    .ren(~rst & ~async_mux),
    .wval(~(rst) & (| credit_gather) & ~async_mux),
    .wdata(credit_gather),
    .rdata(sync_credit_fifo_out),
    .full(sync_credit_fifo_full),   
    .empty(sync_credit_empty)
);
 
assign credit_fifo_out = async_mux ? async_credit_fifo_out : sync_credit_fifo_out;
assign credit_fifo_full = async_mux ? async_credit_fifo_full : sync_credit_fifo_full;
assign credit_empty = async_mux ? async_credit_empty: sync_credit_empty;
assign credit_to_fpga = credit_to_fpga_r;
assign credit_gather[0] = bout_rdy_1 & bout_val_1;
assign credit_gather[1] = bout_rdy_2 & bout_val_2;
assign credit_gather[2] = bout_rdy_3 & bout_val_3;
always@(posedge wr_clk) begin
 
   if(rst) begin
 
        credit_to_fpga_r <= 3'b000;       
   end
   else begin
       if(~credit_empty) begin 
           credit_to_fpga_r <= credit_fifo_out;
       end
       else
           credit_to_fpga_r <= 3'b000;       
   end 
end
endmodule
    
    
 
    
    
    
    
    
    
 
 
 
  
    
 
 
    
    
    
    
    
    
    
 
 
module chip_bridge_out (
    rst, 
    wr_clk,
    rd_clk,
    async_mux,
    bin_data_1,
    bin_val_1,
    bin_rdy_1,
    bin_data_2,
    bin_val_2,
    bin_rdy_2,
    bin_data_3,
    bin_val_3,
    bin_rdy_3,
    data_to_fpga,
    data_channel,
    credit_from_fpga
);  
input rst;
input wr_clk;
input rd_clk;
input async_mux;
output          bin_rdy_1;
output          bin_rdy_2;
output          bin_rdy_3;
output [31:0]   data_to_fpga;
output [ 1:0]    data_channel;
input [63:0]    bin_data_1;
input           bin_val_1;
input [63:0]    bin_data_2;
input           bin_val_2;
input [63:0]    bin_data_3;
input           bin_val_3;
input [2:0]     credit_from_fpga;
wire network_rdy_1;
wire network_rdy_2;
wire network_rdy_3;
wire fifo1_full;
wire fifo2_full;
wire fifo3_full;
wire [63:0] network_data_1;
wire [63:0] network_data_2;
wire [63:0] network_data_3;
wire network_val_1;
wire network_val_2;
wire network_val_3;
wire async_fifo1_full;
wire async_fifo2_full;
wire async_fifo3_full;
wire [63:0] async_network_data_1;
wire [63:0] async_network_data_2;
wire [63:0] async_network_data_3;
wire async_network_val_1;
wire async_network_val_2;
wire async_network_val_3;
wire sync_fifo1_full;
wire sync_fifo2_full;
wire sync_fifo3_full;
wire [63:0] sync_network_data_1;
wire [63:0] sync_network_data_2;
wire [63:0] sync_network_data_3;
wire sync_network_val_1;
wire sync_network_val_2;
wire sync_network_val_3;
wire [63:0] data_to_serial_buffer;
reg  [31:0] serial_buffer_data;
reg  [31:0] serial_buffer_data_f ;
reg   [0:0] serial_buffer_data_counter;
wire  [1:0] channel_to_serial_buffer;
reg   [1:0] serial_buffer_channel ;
reg   [1:0] serial_buffer_channel_dup ;
assign bin_rdy_1 = ~fifo1_full; 
assign bin_rdy_2 = ~fifo2_full; 
assign bin_rdy_3 = ~fifo3_full; 
assign data_to_fpga = serial_buffer_data_f;
assign data_channel = serial_buffer_channel;
bridge_network_chooser separator(
 
    .rst    (rst),
    .clk    (rd_clk),
    .data_out(data_to_serial_buffer),
    .data_channel(channel_to_serial_buffer),
    .din_1  (network_data_1),
    .rdy_1  (network_rdy_1),
    .val_1  (~network_val_1),
    .din_2  (network_data_2),
    .rdy_2  (network_rdy_2),
    .val_2  (~network_val_2),
    .din_3  (network_data_3),
    .rdy_3  (network_rdy_3),
    .val_3  (~network_val_3),
    .credit_from_fpga(credit_from_fpga)
);
 
async_fifo #(
.DSIZE(64),
.ASIZE(4),
.MEMSIZE(8) )
async_fifo_1(
    .rreset(rst),
    .wreset(rst),
    .wclk(wr_clk),
    .rclk(rd_clk),
    .ren(network_rdy_1 && async_mux),
    .wval(bin_val_1 && async_mux),
    .wdata(bin_data_1),
    .rdata(async_network_data_1),
    .wfull(async_fifo1_full),
    .rempty(async_network_val_1)
);
 
 
async_fifo #(
.DSIZE(64),
.ASIZE(4),
.MEMSIZE(8) )
async_fifo_2(
    .rreset(rst),
    .wreset(rst),
    .wclk(wr_clk),
    .rclk(rd_clk),
    .ren(network_rdy_2 && async_mux),
    .wval(bin_val_2 && async_mux),
    .wdata(bin_data_2),
    .rdata(async_network_data_2),
    .wfull(async_fifo2_full),
    .rempty(async_network_val_2)
);
 
 
async_fifo #(
.DSIZE(64),
.ASIZE(4),
.MEMSIZE(8) )
async_fifo_3(
    .rreset(rst),
    .wreset(rst),
    .wclk(wr_clk),
    .rclk(rd_clk),
    .ren(network_rdy_3 && async_mux),
    .wval(bin_val_3 && async_mux),
    .wdata(bin_data_3),
    .rdata(async_network_data_3),
    .wfull(async_fifo3_full),
    .rempty(async_network_val_3)
);
 
 
sync_fifo #(
.DSIZE(64),
.ASIZE(4),
.MEMSIZE(8) )
sync_fifo_1(
    .reset(rst),
    .clk(rd_clk),
    .ren(network_rdy_1 && ~async_mux),
    .wval(bin_val_1 && ~async_mux),
    .wdata(bin_data_1),
    .rdata(sync_network_data_1),
    .full(sync_fifo1_full),
    .empty(sync_network_val_1)
);
 
 
sync_fifo #(
.DSIZE(64),
.ASIZE(4),
.MEMSIZE(8) )
sync_fifo_2(
    .reset(rst),
    .clk(rd_clk),
    .ren(network_rdy_2 && ~async_mux),
    .wval(bin_val_2 && ~async_mux),
    .wdata(bin_data_2),
    .rdata(sync_network_data_2),
    .full(sync_fifo2_full),
    .empty(sync_network_val_2)
);
 
 
sync_fifo #(
.DSIZE(64),
.ASIZE(4),
.MEMSIZE(8) )
sync_fifo_3(
    .reset(rst),
    .clk(rd_clk),
    .ren(network_rdy_3 && ~async_mux),
    .wval(bin_val_3 && ~async_mux),
    .wdata(bin_data_3),
    .rdata(sync_network_data_3),
    .full(sync_fifo3_full),
    .empty(sync_network_val_3)
);
 
assign network_val_1  = async_mux ? async_network_val_1 : sync_network_val_1;
assign network_val_2  = async_mux ? async_network_val_2 : sync_network_val_2;
assign network_val_3  = async_mux ? async_network_val_3 : sync_network_val_3;
assign network_data_1  = async_mux ? async_network_data_1 : sync_network_data_1;
assign network_data_2  = async_mux ? async_network_data_2 : sync_network_data_2;
assign network_data_3  = async_mux ? async_network_data_3 : sync_network_data_3;
assign fifo1_full = async_mux ? async_fifo1_full : sync_fifo1_full;
assign fifo2_full = async_mux ? async_fifo2_full : sync_fifo2_full;
assign fifo3_full = async_mux ? async_fifo3_full : sync_fifo3_full;
always @(posedge rd_clk) begin
 
    if(rst) begin
 
        serial_buffer_data <= 32'd0;
        serial_buffer_data_f <= 32'd0;
        serial_buffer_channel <= 2'd0;
        serial_buffer_channel_dup <= 2'd0;
        serial_buffer_data_counter <= 1'b1;
    end
    else begin
        if( channel_to_serial_buffer != 0 && serial_buffer_data_counter == 1) begin
            
            serial_buffer_data_f <= data_to_serial_buffer[31:0];
            serial_buffer_data <= data_to_serial_buffer[63:32];
            serial_buffer_channel <= channel_to_serial_buffer;
            serial_buffer_channel_dup <= channel_to_serial_buffer;
            serial_buffer_data_counter <= serial_buffer_data_counter + 1'b1;
        end
        else if( serial_buffer_channel_dup != 0 && serial_buffer_data_counter != 1'b1) begin
            serial_buffer_data_f <= serial_buffer_data;
            serial_buffer_data_counter <= serial_buffer_data_counter + 1'b1;
        end
        else begin
            serial_buffer_data_counter <= 1'b1;
            serial_buffer_channel <= channel_to_serial_buffer;
            serial_buffer_channel_dup <= channel_to_serial_buffer;
        end
    end
end 
endmodule
module bridge_network_chooser(
    rst,
    clk,
    data_out,
    data_channel,
    din_1,
    rdy_1,
    val_1,
    din_2,
    rdy_2,
    val_2,
    din_3,
    rdy_3,
    val_3,
    credit_from_fpga
);
input rst;
input clk;
input [63:0] din_1;
input [63:0] din_2;
input [63:0] din_3;
input        val_1;
input        val_2;
input        val_3;
input [ 2:0] credit_from_fpga;
output [63:0] data_out;
output [ 1:0] data_channel;
output        rdy_1;
output        rdy_2;
output        rdy_3;
reg [8:0] credit_1; 
reg [8:0] credit_2;
reg [8:0] credit_3;
wire [1:0] select;
reg  [1:0] select_reg;
reg  [0:0] select_counter;
reg sel_23;
reg sel_13;
reg sel_12;
reg [1:0] sel_123;
assign data_out =   rdy_1 ? din_1 :
                    rdy_2 ? din_2 :
                    rdy_3 ? din_3 : 64'd0;
assign data_channel = select; 
assign rdy_1 = (select == 2'b01 && select_counter == 1'b0) ? 1'b1 : 1'b0;
assign rdy_2 = (select == 2'b10 && select_counter == 1'b0) ? 1'b1 : 1'b0;
assign rdy_3 = (select == 2'b11 && select_counter == 1'b0) ? 1'b1 : 1'b0;
assign select = ( (select_counter != 1'b0         ) )   ? select_reg :
                ( (credit_1 == 9'd255 || ~val_1) &&            
                  (credit_2 == 9'd255 || ~val_2) && 
                  (credit_3 == 9'd255 || ~val_3) )   ? 2'b00  :
                ( (credit_2 == 9'd255 || ~val_2) &&            
                  (credit_3 == 9'd255 || ~val_3) )   ? 2'b01  :
                ( (credit_1 == 9'd255 || ~val_1) &&
                  (credit_3 == 9'd255 || ~val_3) )   ? 2'b10  :
                ( (credit_1 == 9'd255 || ~val_1) &&
                  (credit_2 == 9'd255 || ~val_2) )   ? 2'b11  :
                ( (credit_1 == 9'd255 || ~val_1) )   ? (sel_23 ? 2'b11 : 2'b10) : 
                ( (credit_2 == 9'd255 || ~val_2) )   ? (sel_13 ? 2'b11 : 2'b01) :
                ( (credit_3 == 9'd255 || ~val_3) )   ? (sel_12 ? 2'b10 : 2'b01) :
                                                sel_123; 
always @(posedge clk) begin
    if(rst) begin
        select_reg <= 2'd0;
    end
    else begin
        select_reg <= select;
    end
end
always @(posedge clk) begin
    if(rst) begin
        credit_1 <= 9'd0;
        credit_2 <= 9'd0;
        credit_3 <= 9'd0;
        sel_23 <= 0;
        sel_13 <= 0;
        sel_12 <= 0;
        sel_123 <= 0;
        select_counter <= 0;
    end
    else begin
        
        if(select == 0) begin
            select_counter <= 0;
        end
        else begin
            select_counter <= select_counter + 2'b01; 
        end
        
        if(credit_from_fpga[0] & ~(rdy_1 & val_1)) begin
            credit_1 <= credit_1 - 9'd1;
        end
        if(credit_from_fpga[1] & ~(rdy_2 & val_2)) begin
            credit_2 <= credit_2 - 9'd1;
        end
        if(credit_from_fpga[2] & ~(rdy_3 & val_3)) begin
            credit_3 <= credit_3 - 9'd1;
        end
        
        if((credit_1 < 9'd255) &&
           (credit_2 < 9'd255) &&
           (credit_3 < 9'd255) &&
           (sel_123 == 0)         )
            sel_123 <= 2'b01;
        
        if(rdy_1 & val_1) begin
            sel_13 <= 1;
            sel_12 <= 1;
            if (sel_123 == 2'b01) begin
                sel_123 <= 2'b10;
            end
            if(~credit_from_fpga[0]) begin
                credit_1 <= credit_1 + 9'd1;
            end
        end 
        if(rdy_2 & val_2) begin
            sel_23 <= 1;
            sel_12 <= 0;
            if (sel_123 == 2'b10) begin
                sel_123 <= 2'b11;
            end
            if( ~credit_from_fpga[1]) begin
                credit_2 <= credit_2 + 9'd1;
            end
        end
        if(rdy_3 & val_3) begin
            sel_23 <= 0;
            sel_13 <= 0;
            if (sel_123 == 2'b11) begin
                sel_123 <= 2'b01;
            end
            if (~credit_from_fpga[2]) begin
                credit_3 <= credit_3 + 9'd1;
            end
        end
    end
end 
endmodule
module chip_bridge(
    rst_n,
    chip_clk,
    intcnct_clk,
    async_mux,
    network_out_1,
    network_out_2,
    network_out_3,
    data_out_val_1,
    data_out_val_2,
    data_out_val_3,
    data_out_rdy_1,
    data_out_rdy_2,
    data_out_rdy_3,
    intcnct_data_in,
    intcnct_channel_in,
    intcnct_credit_back_in,
    network_in_1,
    network_in_2,
    network_in_3,
    data_in_val_1,
    data_in_val_2,
    data_in_val_3,
    data_in_rdy_1,
    data_in_rdy_2,
    data_in_rdy_3,
    intcnct_data_out,
    intcnct_channel_out,
    intcnct_credit_back_out
);
input           rst_n;
input           chip_clk;
input           intcnct_clk;
input           async_mux;
input  [63:0]   network_out_1;
input  [63:0]   network_out_2;
input  [63:0]   network_out_3;
input           data_out_val_1;
input           data_out_val_2;
input           data_out_val_3;
output          data_out_rdy_1;
output          data_out_rdy_2;
output          data_out_rdy_3;
output [31:0]   intcnct_data_out;
output [1:0]    intcnct_channel_out;
input  [2:0]    intcnct_credit_back_out;
output [63:0]   network_in_1;
output [63:0]   network_in_2;
output [63:0]   network_in_3;
output          data_in_val_1;
output          data_in_val_2;
output          data_in_val_3;
input           data_in_rdy_1;
input           data_in_rdy_2;
input           data_in_rdy_3;
input  [31:0]   intcnct_data_in;
input  [1:0]    intcnct_channel_in;
output [2:0]    intcnct_credit_back_in;
chip_bridge_out chip_fpga_out(
    .rst(~rst_n), 
    .wr_clk(chip_clk),
    .rd_clk(intcnct_clk),
    .async_mux(async_mux),
    .bin_data_1(network_out_1),
    .bin_val_1(data_out_val_1),
    .bin_rdy_1(data_out_rdy_1),
    .bin_data_2(network_out_2),
    .bin_val_2(data_out_val_2),
    .bin_rdy_2(data_out_rdy_2),
    .bin_data_3(network_out_3),
    .bin_val_3(data_out_val_3),
    .bin_rdy_3(data_out_rdy_3),
    .data_to_fpga(intcnct_data_out),
    .data_channel(intcnct_channel_out),
    .credit_from_fpga(intcnct_credit_back_out)
    );  
chip_bridge_in chip_fpga_in(
    .rst(~rst_n), 
    .wr_clk(intcnct_clk),
    .rd_clk(chip_clk),
    .async_mux(async_mux),
    .bout_data_1(network_in_1),
    .bout_val_1(data_in_val_1),
    .bout_rdy_1(data_in_rdy_1),
    .bout_data_2(network_in_2),
    .bout_val_2(data_in_val_2),
    .bout_rdy_2(data_in_rdy_2),
    .bout_data_3(network_in_3),
    .bout_val_3(data_in_val_3),
    .bout_rdy_3(data_in_rdy_3),
    .data_from_fpga(intcnct_data_in),
    .data_channel(intcnct_channel_in),
    .credit_to_fpga(intcnct_credit_back_in)
    );
endmodule
 
 
 
 
 
 
 
module dynamic_input_control(thanks_all_temp_out,
                             route_req_n_out, route_req_e_out, route_req_s_out, route_req_w_out, route_req_p_out,
                             default_ready_n, default_ready_e, default_ready_s, default_ready_w, default_ready_p,
                             tail_out, clk, reset,
                             my_loc_x_in, my_loc_y_in, my_chip_id_in,
                             abs_x, abs_y, abs_chip_id, final_bits, valid_in,
                             thanks_n, thanks_e, thanks_s, thanks_w, thanks_p,
                             length);
output thanks_all_temp_out;
output route_req_n_out;
output route_req_e_out;
output route_req_s_out;
output route_req_w_out;
output route_req_p_out;
output default_ready_n;
output default_ready_e;
output default_ready_s;
output default_ready_w;
output default_ready_p;
output tail_out;
input clk;
input reset;
input [8-1:0] my_loc_x_in;
input [8-1:0] my_loc_y_in;
input [14-1:0] my_chip_id_in;
input [8-1:0] abs_x;
input [8-1:0] abs_y;
input [14-1:0] abs_chip_id;
input [2:0] final_bits;
input valid_in;
input thanks_n;
input thanks_e;
input thanks_s;
input thanks_w;
input thanks_p;
input [8-1:0] length;
reg [8-1:0] count_f;
reg header_last_f;
reg thanks_all_f;
reg count_zero_f;
reg count_one_f;
reg tail_last_f;
reg [8-1:0] count_temp;
wire header_last_temp;
wire thanks_all_temp;
wire count_zero_temp;
wire count_one_temp;
wire tail_last_temp;
wire header;
wire [8-1:0] count_minus_one;
wire length_zero; 
                  
wire tail;
reg header_temp;
assign thanks_all_temp = thanks_n | thanks_e | thanks_s | thanks_w | thanks_p;
assign header = valid_in & header_temp;
assign count_zero_temp = count_temp == 0;
assign count_one_temp = count_temp == 1;
assign thanks_all_temp_out = thanks_all_temp;
assign tail_out = tail;
assign count_minus_one = count_f - 1;
assign length_zero = length == 0;
assign header_last_temp = header_temp;
assign tail = (header & length_zero) | ((~thanks_all_f) & tail_last_f) | (thanks_all_f & count_one_f);
assign tail_last_temp = tail;
dynamic_input_route_request_calc tail_calc(.route_req_n(route_req_n_out),
                                           .route_req_e(route_req_e_out),
                                           .route_req_s(route_req_s_out),
                                           .route_req_w(route_req_w_out),
                                           .route_req_p(route_req_p_out),
                                           .default_ready_n(default_ready_n),
                                           .default_ready_e(default_ready_e),
                                           .default_ready_s(default_ready_s),
                                           .default_ready_w(default_ready_w),
                                           .default_ready_p(default_ready_p),
                                           .my_loc_x_in(my_loc_x_in),
                                           .my_loc_y_in(my_loc_y_in),
                                           .my_chip_id_in(my_chip_id_in),
                                           .abs_x(abs_x),
                                           .abs_y(abs_y),
                                           .abs_chip_id(abs_chip_id),
                                           .final_bits(final_bits),
                                           .length(length),
                                           .header_in(header));
always @ (header_last_f or thanks_all_f or count_zero_f)
begin
        case({header_last_f, count_zero_f, thanks_all_f})
        3'b000: header_temp <= 1'b0;
        3'b001: header_temp <= 1'b0;
        3'b010: header_temp <= 1'b0;
        3'b011: header_temp <= 1'b1;
        3'b100: header_temp <= 1'b1;
        
        3'b101: header_temp <= 1'b0;
        3'b110: header_temp <= 1'b1;
        3'b111: header_temp <= 1'b1;
        default:
                header_temp <= 1'b1;
        endcase
end
always @ (header or thanks_all_f or count_f or count_minus_one or length)
begin
        if(header)
        begin
                count_temp <= length;
        end
        else
        begin
                if(thanks_all_f)
                begin
                        count_temp <= count_minus_one;
                end
                else
                begin
                        count_temp <= count_f;
                end
        end
end
always @ (posedge clk)
begin
        if(reset)
        begin
                count_f <= 5'd0;
                header_last_f <= 1'b1;
                thanks_all_f <= 1'b0;
                count_zero_f <= 1'b1; 
                count_one_f <= 1'b0;
                tail_last_f <= 1'b0;
        end
        else
        begin
                count_f <= count_temp;
                header_last_f <= header_last_temp;
                thanks_all_f <= thanks_all_temp;
                count_zero_f <= count_zero_temp;
                count_one_f <= count_one_temp;
                tail_last_f <= tail_last_temp;
        end
end
endmodule
 
 
 
 
 
 
 
module dynamic_input_route_request_calc(route_req_n, route_req_e, route_req_s, route_req_w, route_req_p, 
                                        default_ready_n, default_ready_e, default_ready_s, default_ready_w, default_ready_p, 
                                        my_loc_x_in, my_loc_y_in, my_chip_id_in, abs_x, abs_y, abs_chip_id, final_bits, length, header_in);
output route_req_n;
output route_req_e;
output route_req_s;
output route_req_w;
output route_req_p;
output default_ready_n;
output default_ready_e;
output default_ready_s;
output default_ready_w;
output default_ready_p;
input [8-1:0] my_loc_x_in;
input [8-1:0] my_loc_y_in;
input [14-1:0] my_chip_id_in;
input [8-1:0] abs_x;
input [8-1:0] abs_y;
input [14-1:0] abs_chip_id;
input [2:0] final_bits;
input [8-1:0] length;
input header_in;
   
wire more_x;
wire more_y;
wire less_x;
wire less_y;
wire done_x;
wire done_y;
wire off_chip;
wire done;
wire north;
wire east;
wire south;
wire west;
wire proc;
wire north_calc;
wire south_calc;
assign off_chip = abs_chip_id != my_chip_id_in;
assign more_x = off_chip ? 0 > my_loc_x_in : abs_x > my_loc_x_in;
assign more_y = off_chip ? 0 > my_loc_y_in : abs_y > my_loc_y_in;
assign less_x = off_chip ? 0 < my_loc_x_in : abs_x < my_loc_x_in;
assign less_y = off_chip ? 0 < my_loc_y_in : abs_y < my_loc_y_in;
assign done_x = off_chip ? 0 == my_loc_x_in : abs_x == my_loc_x_in;
assign done_y = off_chip ? 0 == my_loc_y_in : abs_y == my_loc_y_in;
assign done = done_x & done_y;
assign north_calc = done_x & less_y;
assign south_calc = done_x & more_y;
assign north = north_calc | ((final_bits == 3'b101) & done);
assign south = south_calc | ((final_bits == 3'b011) & done);
assign east = more_x | ((final_bits == 3'b100) & done);
assign west = less_x | ((final_bits == 3'b010) & done);
assign proc = ((final_bits == 3'b000) & done);
assign route_req_n = header_in & north;
assign route_req_e = header_in & east;
assign route_req_s = header_in & south;
assign route_req_w = header_in & west;
assign route_req_p = header_in & proc;
assign default_ready_n = route_req_n;
assign default_ready_e = route_req_e;
assign default_ready_s = route_req_s;
assign default_ready_w = route_req_w;
assign default_ready_p = route_req_p;
endmodule
   
 
 
 
 
 
 
 
module dynamic_input_top_16(route_req_n_out, route_req_e_out, route_req_s_out, route_req_w_out, route_req_p_out, default_ready_n_out, default_ready_e_out, default_ready_s_out, default_ready_w_out, default_ready_p_out, tail_out, yummy_out, data_out, valid_out, clk, reset, my_loc_x_in, my_loc_y_in, my_chip_id_in, valid_in, data_in, thanks_n, thanks_e, thanks_s, thanks_w, thanks_p);
output route_req_n_out;
output route_req_e_out;
output route_req_s_out;
output route_req_w_out;
output route_req_p_out;
output default_ready_n_out;
output default_ready_e_out;
output default_ready_s_out;
output default_ready_w_out;
output default_ready_p_out;
output tail_out;
output yummy_out;
output [64-1:0] data_out;
output valid_out;
input clk;
input reset;
input [8-1:0] my_loc_x_in;
input [8-1:0] my_loc_y_in;
input [14-1:0] my_chip_id_in;
input valid_in;
input [64-1:0] data_in;
input thanks_n;
input thanks_e;
input thanks_s;
input thanks_w;
input thanks_p;
   
wire thanks_all_temp;
wire valid_out_internal;
wire [64-1:0] data_out_internal;
wire [64-1:0] data_out_internal_pre;
assign valid_out = valid_out_internal;
assign data_out = data_out_internal;
network_input_blk_multi_out #(.LOG2_NUMBER_FIFO_ELEMENTS(4)) NIB(.clk(clk), .reset(reset), .data_in(data_in), .valid_in(valid_in), .yummy_out(yummy_out), .thanks_in(thanks_all_temp), .data_val(data_out_internal_pre), .data_val1(), .data_avail(valid_out_internal));
assign data_out_internal = data_out_internal_pre;
dynamic_input_control control(.thanks_all_temp_out(thanks_all_temp), .route_req_n_out(route_req_n_out), .route_req_e_out(route_req_e_out), .route_req_s_out(route_req_s_out), .route_req_w_out(route_req_w_out), .route_req_p_out(route_req_p_out), .default_ready_n(default_ready_n_out), .default_ready_e(default_ready_e_out), .default_ready_s(default_ready_s_out), .default_ready_w(default_ready_w_out), .default_ready_p(default_ready_p_out), .tail_out(tail_out), .clk(clk), .reset(reset), .my_loc_x_in(my_loc_x_in), .my_loc_y_in(my_loc_y_in), 
    .my_chip_id_in(my_chip_id_in), .abs_x(data_out_internal[64-14-1:64-14-8]), .abs_y(data_out_internal[64-14-8-1:64-14-2*8]), .abs_chip_id(data_out_internal[64-1:64-14]),.final_bits(data_out_internal[64-14-2*8-2:64-14-2*8-4]), .valid_in(valid_out_internal), .thanks_n(thanks_n), .thanks_e(thanks_e), .thanks_s(thanks_s), .thanks_w(thanks_w), .thanks_p(thanks_p), .length(data_out_internal[64-14-2*8-5:64-14-2*8-4-8]));
endmodule
 
 
 
 
 
 
 
module dynamic_input_top_4(route_req_n_out, route_req_e_out, route_req_s_out, route_req_w_out, route_req_p_out,
                           default_ready_n_out, default_ready_e_out, default_ready_s_out, default_ready_w_out, default_ready_p_out,
                           tail_out, yummy_out, data_out, valid_out, clk, reset,
                           my_loc_x_in, my_loc_y_in, my_chip_id_in,  valid_in, data_in,
                           thanks_n, thanks_e, thanks_s, thanks_w, thanks_p);
output route_req_n_out;
output route_req_e_out;
output route_req_s_out;
output route_req_w_out;
output route_req_p_out;
output default_ready_n_out;
output default_ready_e_out;
output default_ready_s_out;
output default_ready_w_out;
output default_ready_p_out;
output tail_out;
output yummy_out;
output [64-1:0] data_out;
output valid_out;
input clk;
input reset;
input [8-1:0] my_loc_x_in;
input [8-1:0] my_loc_y_in;
input [14-1:0] my_chip_id_in;
input valid_in;
input [64-1:0] data_in;
input thanks_n;
input thanks_e;
input thanks_s;
input thanks_w;
input thanks_p;
wire thanks_all_temp;
wire [64-1:0] data_internal;
wire valid_out_internal;
assign valid_out = valid_out_internal;
network_input_blk_multi_out #(.LOG2_NUMBER_FIFO_ELEMENTS(2)) NIB(.clk(clk),
                                      .reset(reset),
                                      .data_in(data_in),
                                      .valid_in(valid_in),
                                      .yummy_out(yummy_out),
                                      .thanks_in(thanks_all_temp),
                                      .data_val(data_out),
                                      .data_val1(data_internal), 
                                      .data_avail(valid_out_internal));
dynamic_input_control control(.thanks_all_temp_out(thanks_all_temp),
                              .route_req_n_out(route_req_n_out), 
                              .route_req_e_out(route_req_e_out), 
                              .route_req_s_out(route_req_s_out), 
                              .route_req_w_out(route_req_w_out), 
                              .route_req_p_out(route_req_p_out),
                              .default_ready_n(default_ready_n_out), 
                              .default_ready_e(default_ready_e_out), 
                              .default_ready_s(default_ready_s_out), 
                              .default_ready_w(default_ready_w_out), 
                              .default_ready_p(default_ready_p_out),
                              .tail_out(tail_out),
                              .clk(clk), .reset(reset),
                              .my_loc_x_in(my_loc_x_in), 
                              .my_loc_y_in(my_loc_y_in), 
                              .my_chip_id_in(my_chip_id_in),
                              .abs_x(data_internal[64-14-1:64-14-8]), 
                              .abs_y(data_internal[64-14-8-1:64-14-2*8]), 
                              .abs_chip_id(data_internal[64-1:64-14]),
                              .final_bits(data_internal[64-14-2*8-2:64-14-2*8-4]),
                              .valid_in(valid_out_internal),
                              .thanks_n(thanks_n), .thanks_e(thanks_e), .thanks_s(thanks_s), .thanks_w(thanks_w), .thanks_p(thanks_p),
                              .length(data_internal[64-14-2*8-5:64-14-2*8-4-8]));
endmodule
 
 
 
 
 
 
 
module dynamic_output_control(thanks_a, thanks_b, thanks_c, thanks_d, thanks_x, valid_out, current_route, ec_wants_to_send_but_cannot, clk, reset, route_req_a_in, route_req_b_in, route_req_c_in, route_req_d_in, route_req_x_in, tail_a_in, tail_b_in, tail_c_in, tail_d_in, tail_x_in, valid_out_temp, default_ready, space_avail);
output thanks_a;
output thanks_b;
output thanks_c;
output thanks_d;
output thanks_x;
output valid_out;
output [2:0] current_route;
output    ec_wants_to_send_but_cannot;
input clk;
input reset;
input route_req_a_in;
input route_req_b_in;
input route_req_c_in;
input route_req_d_in;
input route_req_x_in;
input tail_a_in;
input tail_b_in;
input tail_c_in;
input tail_d_in;
input tail_x_in;
input valid_out_temp;
input default_ready;
input space_avail;
reg [2:0]current_route_f;
reg planned_f;
wire [2:0] current_route_temp;
wire planned_or_default;
wire route_req_all_or_with_planned;
wire route_req_all_but_default;
wire valid_out_internal;
reg new_route_needed;
reg planned_temp;
reg [2:0] new_route;
reg tail_current_route;
reg route_req_a_mask;
reg route_req_b_mask;
reg route_req_c_mask;
reg route_req_d_mask;
reg route_req_x_mask;
reg thanks_a;
reg thanks_b;
reg thanks_c;
reg thanks_d;
reg thanks_x;
reg    ec_wants_to_send_but_cannot;
assign planned_or_default = planned_f | default_ready;
assign valid_out_internal = valid_out_temp & planned_or_default & space_avail;
always @(posedge clk)
  begin
     ec_wants_to_send_but_cannot <= valid_out_temp & planned_or_default & ~space_avail;
  end
assign current_route_temp = (new_route_needed) ? new_route : current_route_f;
assign current_route = current_route_f;
assign route_req_all_or_with_planned = (route_req_a_in & route_req_a_mask) | (route_req_b_in & route_req_b_mask) | (route_req_c_in & route_req_c_mask) | (route_req_d_in & route_req_d_mask) | (route_req_x_in & route_req_x_mask);
assign route_req_all_but_default = route_req_b_in | route_req_c_in | route_req_d_in | route_req_x_in;
assign valid_out = valid_out_internal;
always @ (current_route_f or tail_a_in or tail_b_in or tail_c_in or tail_d_in or tail_x_in)
begin
	case(current_route_f) 
	3'b000:
	begin
		tail_current_route <= tail_a_in;
	end
	3'b001:
	begin
		tail_current_route <= tail_b_in;
	end
	3'b010:
	begin
		tail_current_route <= tail_c_in;
	end
	3'b011:
	begin
		tail_current_route <= tail_d_in;
	end
	3'b100:
	begin
		tail_current_route <= tail_x_in;
	end
	default:
	begin
		tail_current_route <= 1'bx; 
					    
					    
					    
					    
	end
	endcase
end
always @ (current_route_f or valid_out_internal)
begin
	case(current_route_f)
	3'b000:
	begin
		thanks_a <= valid_out_internal;
		thanks_b <= 1'b0;
		thanks_c <= 1'b0;
		thanks_d <= 1'b0;
		thanks_x <= 1'b0;
	end
	3'b001:
	begin
		thanks_a <= 1'b0;
		thanks_b <= valid_out_internal;
		thanks_c <= 1'b0;
		thanks_d <= 1'b0;
		thanks_x <= 1'b0;
	end
	3'b010:
	begin
		thanks_a <= 1'b0;
		thanks_b <= 1'b0;
		thanks_c <= valid_out_internal;
		thanks_d <= 1'b0;
		thanks_x <= 1'b0;
	end
	3'b011:
	begin
		thanks_a <= 1'b0;
		thanks_b <= 1'b0;
		thanks_c <= 1'b0;
		thanks_d <= valid_out_internal;
		thanks_x <= 1'b0;
	end
	3'b100:
	begin
		thanks_a <= 1'b0;
		thanks_b <= 1'b0;
		thanks_c <= 1'b0;
		thanks_d <= 1'b0;
		thanks_x <= valid_out_internal;
	end
	default:
	begin
		thanks_a <= 1'bx;
		thanks_b <= 1'bx;
		thanks_c <= 1'bx;
		thanks_d <= 1'bx;
		thanks_x <= 1'bx;
					
					
					
	end
	endcase
end
always @(current_route_f or route_req_a_in or route_req_b_in or route_req_c_in or route_req_d_in or route_req_x_in)
begin
	case(current_route_f)
	3'b000:
	begin
		new_route <= (route_req_b_in)?3'b001:((route_req_c_in)?3'b010:((route_req_d_in)?3'b011:((route_req_x_in)?3'b100:3'b000)));
	end
	3'b001:
	begin
		new_route <= (route_req_c_in)?3'b010:((route_req_d_in)?3'b011:((route_req_x_in)?3'b100:((route_req_a_in)?3'b000:3'b000)));
	end
	3'b010:
	begin
		new_route <= (route_req_d_in)?3'b011:((route_req_x_in)?3'b100:((route_req_a_in)?3'b000:((route_req_b_in)?3'b001:3'b000)));
	end
	3'b011:
	begin
		new_route <= (route_req_x_in)?3'b100:((route_req_a_in)?3'b000:((route_req_b_in)?3'b001:((route_req_c_in)?3'b010:3'b000)));
	end
	3'b100:
	begin
		new_route <= (route_req_a_in)?3'b000:((route_req_b_in)?3'b001:((route_req_c_in)?3'b010:((route_req_d_in)?3'b011:3'b000)));
	end
	default:
	begin
		new_route <= 3'b000;
			
	end
	endcase
end
always @(current_route_f or planned_f)
begin
	if(planned_f)
	begin
		case(current_route_f)
		3'b000:	
			begin
				route_req_a_mask <= 1'b0;
				route_req_b_mask <= 1'b1;
				route_req_c_mask <= 1'b1;
				route_req_d_mask <= 1'b1;
				route_req_x_mask <= 1'b1;
			end
		3'b001:
			begin
				route_req_a_mask <= 1'b1;
				route_req_b_mask <= 1'b0;
				route_req_c_mask <= 1'b1;
				route_req_d_mask <= 1'b1;
				route_req_x_mask <= 1'b1;
			end
		3'b010:
			begin
				route_req_a_mask <= 1'b1;
				route_req_b_mask <= 1'b1;
				route_req_c_mask <= 1'b0;
				route_req_d_mask <= 1'b1;
				route_req_x_mask <= 1'b1;
			end
		3'b011:
			begin
				route_req_a_mask <= 1'b1;
				route_req_b_mask <= 1'b1;
				route_req_c_mask <= 1'b1;
				route_req_d_mask <= 1'b0;
				route_req_x_mask <= 1'b1;
			end
		3'b100:
			begin
				route_req_a_mask <= 1'b1;
				route_req_b_mask <= 1'b1;
				route_req_c_mask <= 1'b1;
				route_req_d_mask <= 1'b1;
				route_req_x_mask <= 1'b0;
			end
		default:
			begin
				route_req_a_mask <= 1'b1;
				route_req_b_mask <= 1'b1;
				route_req_c_mask <= 1'b1;
				route_req_d_mask <= 1'b1;
				route_req_x_mask <= 1'b1;
			end
		endcase
	end
	else
	begin
		route_req_a_mask <= 1'b1;
		route_req_b_mask <= 1'b1;
		route_req_c_mask <= 1'b1;
		route_req_d_mask <= 1'b1;
		route_req_x_mask <= 1'b1;
	end
end
always @ (planned_f or tail_current_route or valid_out_internal or default_ready)
begin
	case({default_ready, valid_out_internal, tail_current_route, planned_f}) 
	4'b0000:	new_route_needed <= 1'b1;
	4'b0001:	new_route_needed <= 1'b0;
	4'b0010:	new_route_needed <= 1'b1;
	4'b0011:	new_route_needed <= 1'b0;
	4'b0100:	new_route_needed <= 1'b0;	
	4'b0101:	new_route_needed <= 1'b0;	
	4'b0110:	new_route_needed <= 1'b1;
	4'b0111:	new_route_needed <= 1'b1;
	4'b1000:	new_route_needed <= 1'b1;
	4'b1001:	new_route_needed <= 1'b0;
	4'b1010:	new_route_needed <= 1'b1;	
    
	4'b1011:	new_route_needed <= 1'b0;
	4'b1100:	new_route_needed <= 1'b0;
	4'b1101:	new_route_needed <= 1'b0;
	4'b1110:	new_route_needed <= 1'b1;
	4'b1111:	new_route_needed <= 1'b1;
	default:	new_route_needed <= 1'b1;
			
	endcase
end
always @ (planned_f or tail_current_route or valid_out_internal or default_ready or route_req_all_or_with_planned or route_req_all_but_default)
begin
	case({route_req_all_or_with_planned, default_ready, valid_out_internal, tail_current_route, planned_f}) 
	5'b00000:	planned_temp <= 1'b0;
	5'b00001:	planned_temp <= 1'b1;
	5'b00010:	planned_temp <= 1'b0;
	5'b00011:	planned_temp <= 1'b1;
	5'b00100:	planned_temp <= 1'b0;	
	5'b00101:	planned_temp <= 1'b1;
	5'b00110:	planned_temp <= 1'b0;	
	5'b00111:	planned_temp <= 1'b0;
	5'b01000:	planned_temp <= 1'b0;	
	5'b01001:	planned_temp <= 1'b1;
	5'b01010:	planned_temp <= 1'b0;	
	5'b01011:	planned_temp <= 1'b1;
	5'b01100:	planned_temp <= 1'b0;	
	5'b01101:	planned_temp <= 1'b1;
	5'b01110:	planned_temp <= 1'b0;	
	5'b01111:	planned_temp <= 1'b0;	
						
						
						
						
						
	5'b10000:	planned_temp <= 1'b1;
	5'b10001:	planned_temp <= 1'b1;
	5'b10010:	planned_temp <= 1'b1;
	5'b10011:	planned_temp <= 1'b1;
	5'b10100:	planned_temp <= 1'b1;
	5'b10101:	planned_temp <= 1'b1;
	5'b10110:	planned_temp <= 1'b1;
	5'b10111:	planned_temp <= 1'b1;
	5'b11000:	planned_temp <= 1'b1;
	5'b11001:	planned_temp <= 1'b1;
	5'b11010:	planned_temp <= 1'b1;
	5'b11011:	planned_temp <= 1'b1;
	5'b11100:	planned_temp <= 1'b1;
	5'b11101:	planned_temp <= 1'b1;
						
						
						
						
						
	5'b11110:	planned_temp <= route_req_all_but_default;
	5'b11111:	planned_temp <= 1'b1;
	default:	planned_temp <= 1'b0;
	endcase
end
always @(posedge clk)
begin
	if(reset)
	begin
		current_route_f <= 3'd0;
		planned_f <= 1'd0;
	end
	else
	begin
		current_route_f <= current_route_temp;
		planned_f <= planned_temp;
	end
end
endmodule
 
 
 
 
 
 
 
module dynamic_output_datapath(data_out, valid_out_temp, data_a_in, data_b_in, data_c_in, data_d_in, data_x_in, valid_a_in, valid_b_in, valid_c_in, valid_d_in, valid_x_in, current_route_in);
output [64-1:0] data_out;
output valid_out_temp;
input [64-1:0] data_a_in;
input [64-1:0] data_b_in;
input [64-1:0] data_c_in;
input [64-1:0] data_d_in;
input [64-1:0] data_x_in;
input valid_a_in;
input valid_b_in;
input valid_c_in;
input valid_d_in;
input valid_x_in;
input [2:0] current_route_in;
one_of_five #(64) data_mux(.in0(data_a_in), .in1(data_b_in), .in2(data_c_in), .in3(data_d_in), .in4(data_x_in), .sel(current_route_in), .out(data_out));
one_of_five #(1) valid_mux(.in0(valid_a_in), .in1(valid_b_in), .in2(valid_c_in), .in3(valid_d_in), .in4(valid_x_in), .sel(current_route_in), .out(valid_out_temp));
endmodule
 
 
 
 
 
 
 
module dynamic_output_top(data_out, thanks_a_out, thanks_b_out, thanks_c_out, thanks_d_out, thanks_x_out, valid_out, popped_interrupt_mesg_out, popped_memory_ack_mesg_out, popped_memory_ack_mesg_out_sender, ec_wants_to_send_but_cannot, clk, reset, route_req_a_in, route_req_b_in, route_req_c_in, route_req_d_in, route_req_x_in, tail_a_in, tail_b_in, tail_c_in, tail_d_in, tail_x_in, data_a_in, data_b_in, data_c_in, data_d_in, data_x_in, valid_a_in, valid_b_in, valid_c_in, valid_d_in, valid_x_in, default_ready_in, yummy_in);
parameter KILL_HEADERS = 1'b0;
output [64-1:0] data_out;
output thanks_a_out;
output thanks_b_out;
output thanks_c_out;
output thanks_d_out;
output thanks_x_out;
output valid_out;
output popped_interrupt_mesg_out;
output popped_memory_ack_mesg_out;
output [9:0] popped_memory_ack_mesg_out_sender;
output ec_wants_to_send_but_cannot;
input clk;
input reset;
input route_req_a_in;
input route_req_b_in;
input route_req_c_in;
input route_req_d_in;
input route_req_x_in;
input tail_a_in;
input tail_b_in;
input tail_c_in;
input tail_d_in;
input tail_x_in;
input [64-1:0] data_a_in;
input [64-1:0] data_b_in;
input [64-1:0] data_c_in;
input [64-1:0] data_d_in;
input [64-1:0] data_x_in;
input valid_a_in;
input valid_b_in;
input valid_c_in;
input valid_d_in;
input valid_x_in;
input default_ready_in;
input yummy_in;
wire valid_out_temp_connection;
wire [2:0] current_route_connection;
wire space_avail_connection;
wire valid_out_pre;
wire data_out_len_zero;
wire data_out_interrupt_user_bits_set;
wire data_out_memory_ack_user_bits_set;
wire [64-1:0] data_out_internal;
wire valid_out_internal;
reg current_route_req;
assign valid_out_internal = valid_out_pre & ~(KILL_HEADERS & current_route_req);
assign data_out_len_zero = data_out_internal[64-14-2*8-4:64-14-2*8-3-8] == 8'd0;
assign data_out_interrupt_user_bits_set = data_out_internal[23:20] == 4'b1111;
assign data_out_memory_ack_user_bits_set = data_out_internal[23:20] == 4'b1110;
assign popped_interrupt_mesg_out = data_out_interrupt_user_bits_set & data_out_len_zero & valid_out_pre & (KILL_HEADERS & current_route_req);
assign popped_memory_ack_mesg_out = data_out_memory_ack_user_bits_set & data_out_len_zero & valid_out_pre & (KILL_HEADERS & current_route_req);
assign popped_memory_ack_mesg_out_sender = data_out_internal[19:10] & { 10 { KILL_HEADERS} };
assign data_out = data_out_internal;
assign valid_out = valid_out_internal;
space_avail_top space(.valid(valid_out_internal), .clk(clk), .reset(reset), .yummy(yummy_in),.spc_avail(space_avail_connection));
dynamic_output_datapath datapath(.data_out(data_out_internal), .valid_out_temp(valid_out_temp_connection), .data_a_in(data_a_in), .data_b_in(data_b_in), .data_c_in(data_c_in), .data_d_in(data_d_in), .data_x_in(data_x_in), .valid_a_in(valid_a_in), .valid_b_in(valid_b_in), .valid_c_in(valid_c_in), .valid_d_in(valid_d_in), .valid_x_in(valid_x_in), .current_route_in(current_route_connection));
dynamic_output_control control(.thanks_a(thanks_a_out), .thanks_b(thanks_b_out), .thanks_c(thanks_c_out), .thanks_d(thanks_d_out), .thanks_x(thanks_x_out), .valid_out(valid_out_pre), .current_route(current_route_connection), .ec_wants_to_send_but_cannot(ec_wants_to_send_but_cannot), .clk(clk), .reset(reset), .route_req_a_in(route_req_a_in), .route_req_b_in(route_req_b_in), .route_req_c_in(route_req_c_in), .route_req_d_in(route_req_d_in), .route_req_x_in(route_req_x_in), .tail_a_in(tail_a_in), .tail_b_in(tail_b_in), .tail_c_in(tail_c_in), .tail_d_in(tail_d_in), .tail_x_in(tail_x_in), .valid_out_temp(valid_out_temp_connection), .default_ready(default_ready_in), .space_avail(space_avail_connection));
always @ (current_route_connection or route_req_a_in or route_req_b_in or route_req_c_in or route_req_d_in or route_req_x_in)
begin
	case(current_route_connection)
	3'b000:	current_route_req <= route_req_a_in;
	3'b001:	current_route_req <= route_req_b_in;
	3'b010:	current_route_req <= route_req_c_in;
	3'b011:	current_route_req <= route_req_d_in;
	3'b100:	current_route_req <= route_req_x_in;
	default:	current_route_req <= 1'bx;
	endcase
end
endmodule
 
 
 
 
 
 
 
module dynamic_input_control_para(thanks_all_temp_out,
                             route_req_0_out, route_req_1_out, 
                             default_ready_0, default_ready_1, 
                             tail_out, clk, reset,
                             my_loc_x_in, my_loc_y_in, my_chip_id_in,
                             abs_x, abs_y, abs_chip_id, final_bits, valid_in,
                             thanks_0, thanks_1, 
                             length);
output thanks_all_temp_out;
output route_req_0_out;
output route_req_1_out;
output default_ready_0;
output default_ready_1;
output tail_out;
input clk;
input reset;
input [8-1:0] my_loc_x_in;
input [8-1:0] my_loc_y_in;
input [14-1:0] my_chip_id_in;
input [8-1:0] abs_x;
input [8-1:0] abs_y;
input [14-1:0] abs_chip_id;
input [2:0] final_bits;
input valid_in;
input thanks_0;
input thanks_1;
input [8-1:0] length;
reg [8-1:0] count_f;
reg header_last_f;
reg thanks_all_f;
reg count_zero_f;
reg count_one_f;
reg tail_last_f;
reg [8-1:0] count_temp;
wire header_last_temp;
wire thanks_all_temp;
wire count_zero_temp;
wire count_one_temp;
wire tail_last_temp;
wire header;
wire [8-1:0] count_minus_one;
wire length_zero; 
                  
wire tail;
reg header_temp;
assign thanks_all_temp = thanks_0 | thanks_1;
assign header = valid_in & header_temp;
assign count_zero_temp = count_temp == 0;
assign count_one_temp = count_temp == 1;
assign thanks_all_temp_out = thanks_all_temp;
assign tail_out = tail;
assign count_minus_one = count_f - 1;
assign length_zero = length == 0;
assign header_last_temp = header_temp;
assign tail = (header & length_zero) | ((~thanks_all_f) & tail_last_f) | (thanks_all_f & count_one_f);
assign tail_last_temp = tail;
dynamic_input_route_request_calc_para tail_calc(.route_req_0(route_req_0_out),
                                           .route_req_1(route_req_1_out),
                                           .default_ready_0(default_ready_0),
                                           .default_ready_1(default_ready_1),
                                           .my_loc_x_in(my_loc_x_in),
                                           .my_loc_y_in(my_loc_y_in),
                                           .my_chip_id_in(my_chip_id_in),
                                           .abs_x(abs_x),
                                           .abs_y(abs_y),
                                           .abs_chip_id(abs_chip_id),
                                           .final_bits(final_bits),
                                           .length(length),
                                           .header_in(header));
always @ (header_last_f or thanks_all_f or count_zero_f)
begin
        case({header_last_f, count_zero_f, thanks_all_f})
        3'b000: header_temp <= 1'b0;
        3'b001: header_temp <= 1'b0;
        3'b010: header_temp <= 1'b0;
        3'b011: header_temp <= 1'b1;
        3'b100: header_temp <= 1'b1;
        
        3'b101: header_temp <= 1'b0;
        3'b110: header_temp <= 1'b1;
        3'b111: header_temp <= 1'b1;
        default:
                header_temp <= 1'b1;
        endcase
end
always @ (header or thanks_all_f or count_f or count_minus_one or length)
begin
        if(header)
        begin
                count_temp <= length;
        end
        else
        begin
                if(thanks_all_f)
                begin
                        count_temp <= count_minus_one;
                end
                else
                begin
                        count_temp <= count_f;
                end
        end
end
always @ (posedge clk)
begin
        if(reset)
        begin
                count_f <= 5'd0;
                header_last_f <= 1'b1;
                thanks_all_f <= 1'b0;
                count_zero_f <= 1'b1; 
                count_one_f <= 1'b0;
                tail_last_f <= 1'b0;
        end
        else
        begin
                count_f <= count_temp;
                header_last_f <= header_last_temp;
                thanks_all_f <= thanks_all_temp;
                count_zero_f <= count_zero_temp;
                count_one_f <= count_one_temp;
                tail_last_f <= tail_last_temp;
        end
end
endmodule
 
 
 
 
 
 
 
module dynamic_input_route_request_calc_para(route_req_0, route_req_1, 
                                        default_ready_0, default_ready_1, 
                                        my_loc_x_in, my_loc_y_in, my_chip_id_in, abs_x, abs_y, abs_chip_id, final_bits, length, header_in);
output route_req_0;
output route_req_1;
output default_ready_0;
output default_ready_1;
input [8-1:0] my_loc_x_in;
input [8-1:0] my_loc_y_in;
input [14-1:0] my_chip_id_in;
input [8-1:0] abs_x;
input [8-1:0] abs_y;
input [14-1:0] abs_chip_id;
input [2:0] final_bits;
input [8-1:0] length;
input header_in;
wire off_chip;
wire [8*3+3-1:0]              stub;
assign off_chip = abs_chip_id != my_chip_id_in;
assign route_req_0 = header_in & (!off_chip) & (abs_x == 8'd0);
assign route_req_1 = header_in & (off_chip);
assign default_ready_0 = route_req_0;
assign default_ready_1 = route_req_1;
assign stub = {my_loc_x_in, my_loc_y_in, abs_y, final_bits};
endmodule
   
 
 
 
 
 
 
 
module dynamic_input_top_16_para(route_req_0_out, route_req_1_out, default_ready_0_out, default_ready_1_out, tail_out, yummy_out, data_out, valid_out, clk, reset, my_loc_x_in, my_loc_y_in, my_chip_id_in, valid_in, data_in,thanks_0, thanks_1);
output route_req_0_out;
output route_req_1_out;
output default_ready_0_out;
output default_ready_1_out;
output tail_out;
output yummy_out;
output [64-1:0] data_out;
output valid_out;
input clk;
input reset;
input [8-1:0] my_loc_x_in;
input [8-1:0] my_loc_y_in;
input [14-1:0] my_chip_id_in;
input valid_in;
input [64-1:0] data_in;
input thanks_0;
input thanks_1;
   
wire thanks_all_temp;
wire valid_out_internal;
wire [64-1:0] data_out_internal;
wire [64-1:0] data_out_internal_pre;
assign valid_out = valid_out_internal;
assign data_out = data_out_internal;
network_input_blk_multi_out #(.LOG2_NUMBER_FIFO_ELEMENTS(4)) NIB(.clk(clk), .reset(reset), .data_in(data_in), .valid_in(valid_in), .yummy_out(yummy_out), .thanks_in(thanks_all_temp), .data_val(data_out_internal_pre), .data_val1(), .data_avail(valid_out_internal));
assign data_out_internal = data_out_internal_pre;
dynamic_input_control_para control(.thanks_all_temp_out(thanks_all_temp), .route_req_0_out(route_req_0_out), .route_req_1_out(route_req_1_out), .default_ready_0(default_ready_0_out), .default_ready_1(default_ready_1_out), .tail_out(tail_out), .clk(clk), .reset(reset), .my_loc_x_in(my_loc_x_in), .my_loc_y_in(my_loc_y_in), 
    .my_chip_id_in(my_chip_id_in), .abs_x(data_out_internal[64-14-1:64-14-8]), .abs_y(data_out_internal[64-14-8-1:64-14-2*8]), .abs_chip_id(data_out_internal[64-1:64-14]),.final_bits(data_out_internal[64-14-2*8-2:64-14-2*8-4]), .valid_in(valid_out_internal), .thanks_0(thanks_0), .thanks_1(thanks_1), .length(data_out_internal[64-14-2*8-5:64-14-2*8-4-8]));
endmodule
 
 
 
 
 
 
 
module dynamic_input_top_4_para(route_req_0_out, route_req_1_out, 
                           default_ready_0_out, default_ready_1_out, 
                           tail_out, yummy_out, data_out, valid_out, clk, reset,
                           my_loc_x_in, my_loc_y_in, my_chip_id_in,  valid_in, data_in,
                           thanks_0, thanks_1);
output route_req_0_out;
output route_req_1_out;
output default_ready_0_out;
output default_ready_1_out;
output tail_out;
output yummy_out;
output [64-1:0] data_out;
output valid_out;
input clk;
input reset;
input [8-1:0] my_loc_x_in;
input [8-1:0] my_loc_y_in;
input [14-1:0] my_chip_id_in;
input valid_in;
input [64-1:0] data_in;
input thanks_0;
input thanks_1;
wire thanks_all_temp;
wire [64-1:0] data_internal;
wire valid_out_internal;
assign valid_out = valid_out_internal;
network_input_blk_multi_out #(.LOG2_NUMBER_FIFO_ELEMENTS(2)) NIB(.clk(clk),
                                      .reset(reset),
                                      .data_in(data_in),
                                      .valid_in(valid_in),
                                      .yummy_out(yummy_out),
                                      .thanks_in(thanks_all_temp),
                                      .data_val(data_out),
                                      .data_val1(data_internal), 
                                      .data_avail(valid_out_internal));
dynamic_input_control_para control(.thanks_all_temp_out(thanks_all_temp),
                              .route_req_0_out(route_req_0_out), .route_req_1_out(route_req_1_out), 
                              .default_ready_0(default_ready_0_out), .default_ready_1(default_ready_1_out), 
                              .tail_out(tail_out),
                              .clk(clk), .reset(reset),
                              .my_loc_x_in(my_loc_x_in), 
                              .my_loc_y_in(my_loc_y_in), 
                              .my_chip_id_in(my_chip_id_in),
                              .abs_x(data_internal[64-14-1:64-14-8]), 
                              .abs_y(data_internal[64-14-8-1:64-14-2*8]), 
                              .abs_chip_id(data_internal[64-1:64-14]),
                              .final_bits(data_internal[64-14-2*8-2:64-14-2*8-4]),
                              .valid_in(valid_out_internal),
                              .thanks_0(thanks_0), .thanks_1(thanks_1), 
                              .length(data_internal[64-14-2*8-5:64-14-2*8-4-8]));
endmodule
 
 
 
 
 
 
 
module dynamic_output_control_para(thanks_0, thanks_1, 
                              valid_out, current_route, ec_wants_to_send_but_cannot, clk, reset, 
                              route_req_0_in, route_req_1_in, 
                              tail_0_in, tail_1_in, 
                              valid_out_temp, default_ready, space_avail);
output thanks_0;
output thanks_1;
output valid_out;
output [0:0] current_route;
output    ec_wants_to_send_but_cannot;
input clk;
input reset;
input route_req_0_in;
input route_req_1_in;
input tail_0_in;
input tail_1_in;
input valid_out_temp;
input default_ready;
input space_avail;
reg [0:0]current_route_f;
reg planned_f;
wire [0:0] current_route_temp;
wire planned_or_default;
wire route_req_all_or_with_planned;
wire route_req_all_but_default;
wire valid_out_internal;
reg new_route_needed;
reg planned_temp;
reg [0:0] new_route;
reg tail_current_route;
reg route_req_0_mask;
reg route_req_1_mask;
reg thanks_0;
reg thanks_1;
reg    ec_wants_to_send_but_cannot;
assign planned_or_default = planned_f | default_ready;
assign valid_out_internal = valid_out_temp & planned_or_default & space_avail;
always @(posedge clk)
  begin
     ec_wants_to_send_but_cannot <= valid_out_temp & planned_or_default & ~space_avail;
  end
assign current_route_temp = (new_route_needed) ? new_route : current_route_f;
assign current_route = current_route_f;
assign route_req_all_or_with_planned = (route_req_0_in & route_req_0_mask) | (route_req_1_in & route_req_1_mask);
assign route_req_all_but_default = (route_req_1_in);
assign valid_out = valid_out_internal;
always @ (current_route_f or tail_0_in or tail_1_in)
begin
	case(current_route_f) 
	
	1'b0:
	begin
		tail_current_route <= tail_0_in;
	end
	1'b1:
	begin
		tail_current_route <= tail_1_in;
	end
	default:
	begin
		tail_current_route <= 1'bx; 
					    
					    
					    
					    
	end
	endcase
end
always @ (current_route_f or valid_out_internal)
begin
	case(current_route_f)
	
	
	1'b0:
	begin
		thanks_0 <= valid_out_internal;
		thanks_1 <= 1'b0;
	end
	1'b1:
	begin
		thanks_0 <= 1'b0;
		thanks_1 <= valid_out_internal;
	end
	default:
	begin
	
		thanks_0 <= 1'bx;
		thanks_1 <= 1'bx;
	
					
					
					
	end
	endcase
end
always @(current_route_f or route_req_0_in or route_req_1_in)
begin
	case(current_route_f)
	
	
	1'b0:
	begin
		new_route <= (route_req_1_in)?1'b1:1'b0;
	end
	1'b1:
	begin
		new_route <= (route_req_0_in)?1'b0:1'b0;
	end
	default:
	begin
		new_route <= 1'b0;
			
	end
	endcase
end
always @(current_route_f or planned_f)
begin
	if(planned_f)
	begin
		case(current_route_f)
		
		1'b0:
			begin
				route_req_0_mask <= 1'b0;
				route_req_1_mask <= 1'b1;
			end
		1'b1:
			begin
				route_req_0_mask <= 1'b1;
				route_req_1_mask <= 1'b0;
			end
		default:
			begin
				route_req_0_mask <= 1'b1;
				route_req_1_mask <= 1'b1;
			end
		
		endcase
	end
	else
	begin
	
		route_req_0_mask <= 1'b1;
		route_req_1_mask <= 1'b1;
	
	end
end
always @ (planned_f or tail_current_route or valid_out_internal or default_ready)
begin
	case({default_ready, valid_out_internal, tail_current_route, planned_f}) 
	4'b0000:	new_route_needed <= 1'b1;
	4'b0001:	new_route_needed <= 1'b0;
	4'b0010:	new_route_needed <= 1'b1;
	4'b0011:	new_route_needed <= 1'b0;
	4'b0100:	new_route_needed <= 1'b0;	
	4'b0101:	new_route_needed <= 1'b0;	
	4'b0110:	new_route_needed <= 1'b1;
	4'b0111:	new_route_needed <= 1'b1;
	4'b1000:	new_route_needed <= 1'b1;
	4'b1001:	new_route_needed <= 1'b0;
	4'b1010:	new_route_needed <= 1'b1;	
    
	4'b1011:	new_route_needed <= 1'b0;
	4'b1100:	new_route_needed <= 1'b0;
	4'b1101:	new_route_needed <= 1'b0;
	4'b1110:	new_route_needed <= 1'b1;
	4'b1111:	new_route_needed <= 1'b1;
	default:	new_route_needed <= 1'b1;
			
	endcase
end
always @ (planned_f or tail_current_route or valid_out_internal or default_ready or route_req_all_or_with_planned or route_req_all_but_default)
begin
	case({route_req_all_or_with_planned, default_ready, valid_out_internal, tail_current_route, planned_f}) 
	5'b00000:	planned_temp <= 1'b0;
	5'b00001:	planned_temp <= 1'b1;
	5'b00010:	planned_temp <= 1'b0;
	5'b00011:	planned_temp <= 1'b1;
	5'b00100:	planned_temp <= 1'b0;	
	5'b00101:	planned_temp <= 1'b1;
	5'b00110:	planned_temp <= 1'b0;	
	5'b00111:	planned_temp <= 1'b0;
	5'b01000:	planned_temp <= 1'b0;	
	5'b01001:	planned_temp <= 1'b1;
	5'b01010:	planned_temp <= 1'b0;	
	5'b01011:	planned_temp <= 1'b1;
	5'b01100:	planned_temp <= 1'b0;	
	5'b01101:	planned_temp <= 1'b1;
	5'b01110:	planned_temp <= 1'b0;	
	5'b01111:	planned_temp <= 1'b0;	
						
						
						
						
						
	5'b10000:	planned_temp <= 1'b1;
	5'b10001:	planned_temp <= 1'b1;
	5'b10010:	planned_temp <= 1'b1;
	5'b10011:	planned_temp <= 1'b1;
	5'b10100:	planned_temp <= 1'b1;
	5'b10101:	planned_temp <= 1'b1;
	5'b10110:	planned_temp <= 1'b1;
	5'b10111:	planned_temp <= 1'b1;
	5'b11000:	planned_temp <= 1'b1;
	5'b11001:	planned_temp <= 1'b1;
	5'b11010:	planned_temp <= 1'b1;
	5'b11011:	planned_temp <= 1'b1;
	5'b11100:	planned_temp <= 1'b1;
	5'b11101:	planned_temp <= 1'b1;
						
						
						
						
						
	5'b11110:	planned_temp <= route_req_all_but_default;
	5'b11111:	planned_temp <= 1'b1;
	default:	planned_temp <= 1'b0;
	endcase
end
always @(posedge clk)
begin
	if(reset)
	begin
		current_route_f <= 3'd0;
		planned_f <= 1'd0;
	end
	else
	begin
		current_route_f <= current_route_temp;
		planned_f <= planned_temp;
	end
end
endmodule
 
 
 
 
 
 
 
module dynamic_output_datapath_para(data_out, valid_out_temp, data_0_in, data_1_in, valid_0_in, valid_1_in, current_route_in);
output [64-1:0] data_out;
output valid_out_temp;
input [64-1:0] data_0_in;
input [64-1:0] data_1_in;
input valid_0_in;
input valid_1_in;
input [0:0] current_route_in;
one_of_n #(64) data_mux(.in0(data_0_in), .in1(data_1_in), .sel(current_route_in), .out(data_out));
one_of_n #(1) valid_mux(.in0(valid_0_in), .in1(valid_1_in), .sel(current_route_in), .out(valid_out_temp));
endmodule
 
 
 
 
 
 
 
module dynamic_output_top_para(data_out, 
                          thanks_0_out, thanks_1_out, 
                          valid_out, popped_interrupt_mesg_out, popped_memory_ack_mesg_out, popped_memory_ack_mesg_out_sender, ec_wants_to_send_but_cannot, clk, reset, 
                          route_req_0_in, route_req_1_in, 
                          tail_0_in, tail_1_in, 
                          data_0_in, data_1_in, 
                          valid_0_in, valid_1_in, 
                          default_ready_in, yummy_in);
parameter KILL_HEADERS = 1'b0;
output [64-1:0] data_out;
output thanks_0_out;
output thanks_1_out;
output valid_out;
output popped_interrupt_mesg_out;
output popped_memory_ack_mesg_out;
output [9:0] popped_memory_ack_mesg_out_sender;
output ec_wants_to_send_but_cannot;
input clk;
input reset;
input route_req_0_in;
input route_req_1_in;
input tail_0_in;
input tail_1_in;
input [64-1:0] data_0_in;
input [64-1:0] data_1_in;
input valid_0_in;
input valid_1_in;
input default_ready_in;
input yummy_in;
wire valid_out_temp_connection;
wire [0:0] current_route_connection;
wire space_avail_connection;
wire valid_out_pre;
wire data_out_len_zero;
wire data_out_interrupt_user_bits_set;
wire data_out_memory_ack_user_bits_set;
wire [64-1:0] data_out_internal;
wire valid_out_internal;
reg current_route_req;
assign valid_out_internal = valid_out_pre & ~(KILL_HEADERS & current_route_req);
assign data_out_len_zero = data_out_internal[64-14-2*8-4:64-14-2*8-3-8] == 8'd0;
assign data_out_interrupt_user_bits_set = data_out_internal[23:20] == 4'b1111;
assign data_out_memory_ack_user_bits_set = data_out_internal[23:20] == 4'b1110;
assign popped_interrupt_mesg_out = data_out_interrupt_user_bits_set & data_out_len_zero & valid_out_pre & (KILL_HEADERS & current_route_req);
assign popped_memory_ack_mesg_out = data_out_memory_ack_user_bits_set & data_out_len_zero & valid_out_pre & (KILL_HEADERS & current_route_req);
assign popped_memory_ack_mesg_out_sender = data_out_internal[19:10] & { 10 { KILL_HEADERS} };
assign data_out = data_out_internal;
assign valid_out = valid_out_internal;
space_avail_top space(.valid(valid_out_internal), .clk(clk), .reset(reset), .yummy(yummy_in),.spc_avail(space_avail_connection));
dynamic_output_datapath_para datapath(.data_out(data_out_internal), .valid_out_temp(valid_out_temp_connection), .data_0_in(data_0_in), .data_1_in(data_1_in), .valid_0_in(valid_0_in), .valid_1_in(valid_1_in), .current_route_in(current_route_connection));
dynamic_output_control_para control(.thanks_0(thanks_0_out), .thanks_1(thanks_1_out), 
                               .valid_out(valid_out_pre), .current_route(current_route_connection), .ec_wants_to_send_but_cannot(ec_wants_to_send_but_cannot), .clk(clk), .reset(reset), 
                               .route_req_0_in(route_req_0_in), .route_req_1_in(route_req_1_in), 
                               .tail_0_in(tail_0_in), .tail_1_in(tail_1_in), 
                               .valid_out_temp(valid_out_temp_connection), .default_ready(default_ready_in), .space_avail(space_avail_connection));
always @ (current_route_connection or route_req_0_in or route_req_1_in)
begin
	case(current_route_connection)
    
	1'b0:    current_route_req <= route_req_0_in;
	1'b1:    current_route_req <= route_req_1_in;
    
	default:	current_route_req <= 1'bx;
	endcase
end
endmodule
module fpga_bridge(
    
    input                               rst_n,
    input                               fpga_out_clk,
    input                               fpga_in_clk,
    input                               intf_out_clk,
    input                               intf_in_clk,
    
    input  [64-1:0]        fpga_intf_data_noc1,
    input  [64-1:0]        fpga_intf_data_noc2,
    input  [64-1:0]        fpga_intf_data_noc3,
    input                               fpga_intf_val_noc1,
    input                               fpga_intf_val_noc2,
    input                               fpga_intf_val_noc3,
    output                              fpga_intf_rdy_noc1,
    output                              fpga_intf_rdy_noc2,
    output                              fpga_intf_rdy_noc3,
    
    output [31:0]                       fpga_intf_data,
    output [1:0]                        fpga_intf_channel,
    input  [2:0]                        fpga_intf_credit_back,
    
    output [64-1:0]        intf_fpga_data_noc1,
    output [64-1:0]        intf_fpga_data_noc2,
    output [64-1:0]        intf_fpga_data_noc3,
    output                              intf_fpga_val_noc1,
    output                              intf_fpga_val_noc2,
    output                              intf_fpga_val_noc3,
    input                               intf_fpga_rdy_noc1,
    input                               intf_fpga_rdy_noc2,
    input                               intf_fpga_rdy_noc3,
    
    input  [31:0]                       intf_fpga_data,
    input  [1:0]                        intf_fpga_channel,
    output [2:0]                        intf_fpga_credit_back
);
parameter SEND_CREDIT_THRESHOLD = 9'd255;
fpga_bridge_send_32 #(
    .FULL_THRESHOLD(SEND_CREDIT_THRESHOLD)
)fpga_chip_out(
    .rst(~rst_n),
    .wr_clk(fpga_out_clk),
    .rd_clk(intf_out_clk),
    .credit_wr_clk(intf_in_clk),
    .bin_data_1(fpga_intf_data_noc1),
    .bin_val_1(fpga_intf_val_noc1),
    .bin_rdy_1(fpga_intf_rdy_noc1),
    .bin_data_2(fpga_intf_data_noc2),
    .bin_val_2(fpga_intf_val_noc2),
    .bin_rdy_2(fpga_intf_rdy_noc2),
    .bin_data_3(fpga_intf_data_noc3),
    .bin_val_3(fpga_intf_val_noc3),
    .bin_rdy_3(fpga_intf_rdy_noc3),
    .data_to_chip(fpga_intf_data),
    .data_channel(fpga_intf_channel),
    .credit_from_chip(fpga_intf_credit_back)
    );
fpga_bridge_rcv_32 fpga_chip_in (
    .rst(~rst_n),
    .wr_clk(intf_in_clk),
    .rd_clk(fpga_in_clk),
    .credit_rd_clk(intf_out_clk),
    .bout_data_1(intf_fpga_data_noc1),
    .bout_val_1(intf_fpga_val_noc1),
    .bout_rdy_1(intf_fpga_rdy_noc1),
    .bout_data_2(intf_fpga_data_noc2),
    .bout_val_2(intf_fpga_val_noc2),
    .bout_rdy_2(intf_fpga_rdy_noc2),
    .bout_data_3(intf_fpga_data_noc3),
    .bout_val_3(intf_fpga_val_noc3),
    .bout_rdy_3(intf_fpga_rdy_noc3),
    .data_from_chip(intf_fpga_data),
    .data_channel(intf_fpga_channel),
    .credit_to_chip(intf_fpga_credit_back)
);
endmodule
module fpu (
	pcx_fpio_data_rdy_px2,
	pcx_fpio_data_px2,
	arst_l,
	grst_l,
	gclk,
	cluster_cken,
	fp_cpx_req_cq,
	fp_cpx_data_ca,
	ctu_tst_pre_grst_l,
	global_shift_enable,
	ctu_tst_scan_disable,
	ctu_tst_scanmode,
	ctu_tst_macrotest,
	ctu_tst_short_chain,
	si,
	so
);
input		pcx_fpio_data_rdy_px2;	
input [123:0]	pcx_fpio_data_px2;	
input		arst_l;			
input		grst_l;			
input		gclk;			
input		cluster_cken;			
output [7:0]	fp_cpx_req_cq;		
output [144:0]	fp_cpx_data_ca;		
input						ctu_tst_pre_grst_l;
input						global_shift_enable;
input						ctu_tst_scan_disable;
input						ctu_tst_scanmode;
input 					ctu_tst_macrotest;
input 					ctu_tst_short_chain;
input           si;                     
output          so;                     
wire		inq_add;		
wire		inq_mul;		
wire		inq_div;		
wire [4:0]	inq_id;			
wire [1:0]	inq_rnd_mode;		
wire [1:0]	inq_fcc;		
wire [7:0]	inq_op;			
wire		inq_in1_exp_neq_ffs;	
wire		inq_in1_exp_eq_0;	
wire		inq_in1_53_0_neq_0;	
wire		inq_in1_50_0_neq_0;	
wire		inq_in1_53_32_neq_0;	
wire [63:0]	inq_in1;		
wire		inq_in2_exp_neq_ffs;	
wire		inq_in2_exp_eq_0;	
wire		inq_in2_53_0_neq_0;	
wire		inq_in2_50_0_neq_0;	
wire		inq_in2_53_32_neq_0;	
wire [63:0]	inq_in2;		
wire  		fadd_clken_l;		
wire 		fmul_clken_l;		
wire 		fdiv_clken_l;		
wire [4:0] fp_id_in; 
wire [1:0] fp_rnd_mode_in; 
wire [1:0] fp_fcc_in; 
wire [7:0] fp_op_in; 
wire [68:0] fp_src1_in; 
wire [68:0] fp_src2_in; 
wire [3:0] inq_rdaddr; 
wire [3:0] inq_wraddr; 
wire inq_read_en; 
wire inq_we; 
wire [154:0] inq_dout; 
wire [4:0] inq_dout_unused; 
wire		a1stg_step;		
wire		a6stg_fadd_in;		
wire [9:0]	add_id_out_in;		
wire		a6stg_fcmpop;		
wire [4:0]	add_exc_out;		
wire		a6stg_dbl_dst;		
wire		a6stg_sng_dst;		
wire		a6stg_long_dst;		
wire		a6stg_int_dst;		
wire		add_sign_out;		
wire [10:0]	add_exp_out;		
wire [63:0]	add_frac_out;		
wire [1:0]	add_cc_out;		
wire [1:0]	add_fcc_out;		
wire		add_pipe_active;        
wire		m1stg_step;		
wire		m6stg_fmul_in;		
wire [9:0]	m6stg_id_in;		
wire [4:0]	mul_exc_out;		
wire		m6stg_fmul_dbl_dst;	
wire		m6stg_fmuls;		
wire		mul_sign_out;		
wire [10:0]	mul_exp_out;		
wire [51:0]	mul_frac_out;		
wire		mul_pipe_active;        
wire		d1stg_step;		
wire		d8stg_fdiv_in;		
wire [9:0]	div_id_out_in;		
wire [4:0]	div_exc_out;		
wire		d8stg_fdivd;		
wire		d8stg_fdivs;		
wire		div_sign_out;		
wire [10:0]	div_exp_out;		
wire [51:0]	div_frac_out;		
wire		div_pipe_active;        
wire [7:0]	fp_cpx_req_cq_unbuf;		
wire		add_dest_rdy;		
wire		mul_dest_rdy;		
wire		div_dest_rdy;		
wire [144:0]	fp_cpx_data_ca_unbuf;		
wire rclk; 
wire		sehold; 
wire fpu_grst_l;
wire [63:0] inq_in1_add_buf1;
wire [63:0] inq_in1_mul_buf1;
wire [63:0] inq_in1_div_buf1;
wire [63:0] inq_in2_add_buf1;
wire [63:0] inq_in2_mul_buf1;
wire [63:0] inq_in2_div_buf1;
wire [4:0] inq_id_add_buf1;
wire [4:0] inq_id_mul_buf1;
wire [4:0] inq_id_div_buf1;
wire [7:0] inq_op_add_buf1;
wire [7:0] inq_op_mul_buf1;
wire [7:0] inq_op_div_buf1;
wire [1:0] inq_rnd_mode_add_buf1;
wire [1:0] inq_rnd_mode_mul_buf1;
wire [1:0] inq_rnd_mode_div_buf1;
wire inq_in1_50_0_neq_0_add_buf1;
wire inq_in1_50_0_neq_0_mul_buf1;
wire inq_in1_50_0_neq_0_div_buf1;
wire inq_in1_53_0_neq_0_add_buf1;
wire inq_in1_53_0_neq_0_mul_buf1;
wire inq_in1_53_0_neq_0_div_buf1;
wire inq_in1_53_32_neq_0_add_buf1;
wire inq_in1_53_32_neq_0_mul_buf1;
wire inq_in1_53_32_neq_0_div_buf1;
wire inq_in1_exp_eq_0_add_buf1;
wire inq_in1_exp_eq_0_mul_buf1;
wire inq_in1_exp_eq_0_div_buf1;
wire inq_in1_exp_neq_ffs_add_buf1;
wire inq_in1_exp_neq_ffs_mul_buf1;
wire inq_in1_exp_neq_ffs_div_buf1;
wire inq_in2_50_0_neq_0_add_buf1;
wire inq_in2_50_0_neq_0_mul_buf1;
wire inq_in2_50_0_neq_0_div_buf1;
wire inq_in2_53_0_neq_0_add_buf1;
wire inq_in2_53_0_neq_0_mul_buf1;
wire inq_in2_53_0_neq_0_div_buf1;
wire inq_in2_53_32_neq_0_add_buf1;
wire inq_in2_53_32_neq_0_mul_buf1;
wire inq_in2_53_32_neq_0_div_buf1;
wire inq_in2_exp_eq_0_add_buf1;
wire inq_in2_exp_eq_0_mul_buf1;
wire inq_in2_exp_eq_0_div_buf1;
wire inq_in2_exp_neq_ffs_add_buf1;
wire inq_in2_exp_neq_ffs_mul_buf1;
wire inq_in2_exp_neq_ffs_div_buf1;
wire [123:0] pcx_fpio_data_px2_buf1;
wire [155:0] inq_sram_din_buf1;
wire         pcx_fpio_data_rdy_px2_buf1;
wire         arst_l_in_buf3;
wire         fpu_grst_l_in_buf2;
wire         se_in_buf3;
wire         manual_scan_0;
wire         scan_manual_1;
wire         se;
wire         si_buf1;
wire         scan_inq_sram_w;
wire         rst_tri_en;
wire         arst_l_add_buf4;
wire         fpu_grst_l_add_buf3;
wire         se_add_exp_buf2;
wire         se_add_frac_buf2;
wire         scan_manual_2;
wire         fmul_clken_l_buf1;
wire         arst_l_mul_buf2;
wire         fpu_grst_l_mul_buf1;
wire         se_mul_buf4;
wire         se_mul64_buf2;
wire         scan_manual_3;
wire         fdiv_clken_l_div_frac_buf1;
wire         fdiv_clken_l_div_exp_buf1;
wire         arst_l_div_buf2;
wire         se_div_buf5;
wire         scan_manual_4;
wire         arst_l_out_buf3;
wire         se_out_buf2;
wire         scan_manual_5;
wire         ctu_tst_pre_grst_l_buf1;
wire         global_shift_enable_buf1;
wire         ctu_tst_scan_disable_buf1;
wire         ctu_tst_scanmode_buf1;
wire         ctu_tst_macrotest_buf1;
wire         ctu_tst_short_chain_buf1;
wire         scan_manual_6_buf1;
wire         so_unbuf;
wire         scan_manual_6;
wire         grst_l_buf1;
wire         cluster_cken_buf1;
wire         se_cluster_header_buf2;
wire         arst_l_cluster_header_buf2;
fpu_in fpu_in (
	.pcx_fpio_data_rdy_px2		(pcx_fpio_data_rdy_px2_buf1),
	.pcx_fpio_data_px2		(pcx_fpio_data_px2_buf1[123:0]),
	.a1stg_step			(a1stg_step),
	.m1stg_step			(m1stg_step),
	.d1stg_step			(d1stg_step),
	.add_pipe_active		(add_pipe_active),
	.mul_pipe_active		(mul_pipe_active),
	.div_pipe_active		(div_pipe_active),
	.inq_dout    (inq_dout[154:0]),
	.sehold (sehold),
	.arst_l				(arst_l_in_buf3),
	.grst_l				(fpu_grst_l_in_buf2),
	.rclk				(rclk),
	.fadd_clken_l			(fadd_clken_l),
	.fmul_clken_l			(fmul_clken_l),
	.fdiv_clken_l			(fdiv_clken_l),
	.inq_add			(inq_add),
	.inq_mul			(inq_mul),
	.inq_div			(inq_div),
	.inq_id				(inq_id[4:0]),
	.inq_rnd_mode			(inq_rnd_mode[1:0]),
	.inq_fcc			(inq_fcc[1:0]),
	.inq_op				(inq_op[7:0]),
	.inq_in1_exp_neq_ffs		(inq_in1_exp_neq_ffs),
	.inq_in1_exp_eq_0		(inq_in1_exp_eq_0),
	.inq_in1_53_0_neq_0		(inq_in1_53_0_neq_0),
	.inq_in1_50_0_neq_0		(inq_in1_50_0_neq_0),
	.inq_in1_53_32_neq_0		(inq_in1_53_32_neq_0),
	.inq_in1			(inq_in1[63:0]),
	.inq_in2_exp_neq_ffs		(inq_in2_exp_neq_ffs),
	.inq_in2_exp_eq_0		(inq_in2_exp_eq_0),
	.inq_in2_53_0_neq_0		(inq_in2_53_0_neq_0),
	.inq_in2_50_0_neq_0		(inq_in2_50_0_neq_0),
	.inq_in2_53_32_neq_0		(inq_in2_53_32_neq_0),
	.inq_in2			(inq_in2[63:0]),
	.fp_id_in (fp_id_in[4:0]),
	.fp_rnd_mode_in (fp_rnd_mode_in[1:0]),
	.fp_fcc_in (fp_fcc_in[1:0]),
	.fp_op_in (fp_op_in[7:0]),
	.fp_src1_in (fp_src1_in[68:0]),
	.fp_src2_in (fp_src2_in[68:0]),
	.inq_rdaddr (inq_rdaddr[3:0]),
	.inq_wraddr (inq_wraddr[3:0]),
	.inq_read_en (inq_read_en),
	.inq_we (inq_we),
	.se (se_in_buf3),
  .si (manual_scan_0),
  .so (scan_manual_1)
);
bw_r_rf16x160 i_fpu_inq_sram (
	.din ({inq_sram_din_buf1[155:0], 4'b0000}),
	.rd_adr (inq_rdaddr[3:0]),
	.wr_adr (inq_wraddr[3:0]),
	.read_en (inq_read_en),
	.wr_en (inq_we),
	.word_wen (4'hf),
	.byte_wen (20'hfffff),
	.rd_clk (rclk),
	.wr_clk (rclk),
	.se (se),
	.si_r (si_buf1),
	.si_w (scan_inq_sram_w),
	.reset_l (arst_l_in_buf3),
	.sehold (sehold),
	.rst_tri_en (rst_tri_en),
	.dout ({inq_dout[154:0], inq_dout_unused[4:0]}),
	.so_r (scan_inq_sram_w),
	.so_w (manual_scan_0)
);
fpu_add fpu_add (
	.inq_op				(inq_op_add_buf1[7:0]),
	.inq_rnd_mode			(inq_rnd_mode_add_buf1[1:0]),
	.inq_id				(inq_id_add_buf1[4:0]),
	.inq_fcc			(inq_fcc[1:0]),
	.inq_in1			(inq_in1_add_buf1[63:0]),
	.inq_in1_50_0_neq_0		(inq_in1_50_0_neq_0_add_buf1),
	.inq_in1_53_32_neq_0		(inq_in1_53_32_neq_0_add_buf1),
	.inq_in1_exp_eq_0		(inq_in1_exp_eq_0_add_buf1),
	.inq_in1_exp_neq_ffs		(inq_in1_exp_neq_ffs_add_buf1),
	.inq_in2			(inq_in2_add_buf1[63:0]),
	.inq_in2_50_0_neq_0		(inq_in2_50_0_neq_0_add_buf1),
	.inq_in2_53_32_neq_0		(inq_in2_53_32_neq_0_add_buf1),
	.inq_in2_exp_eq_0		(inq_in2_exp_eq_0_add_buf1),
	.inq_in2_exp_neq_ffs		(inq_in2_exp_neq_ffs_add_buf1),
	.inq_add			(inq_add),
	.add_dest_rdy			(add_dest_rdy),
	.fadd_clken_l			(fadd_clken_l),
	.arst_l				(arst_l_add_buf4),
	.grst_l				(fpu_grst_l_add_buf3),
	.rclk				(rclk),
	.add_pipe_active                (add_pipe_active),
	.a1stg_step			(a1stg_step),
	.a6stg_fadd_in			(a6stg_fadd_in),
	.add_id_out_in			(add_id_out_in[9:0]),
	.a6stg_fcmpop			(a6stg_fcmpop),
	.add_exc_out			(add_exc_out[4:0]),
	.a6stg_dbl_dst			(a6stg_dbl_dst),
	.a6stg_sng_dst			(a6stg_sng_dst),
	.a6stg_long_dst			(a6stg_long_dst),
	.a6stg_int_dst			(a6stg_int_dst),
	.add_sign_out			(add_sign_out),
	.add_exp_out			(add_exp_out[10:0]),
	.add_frac_out			(add_frac_out[63:0]),
	.add_cc_out			(add_cc_out[1:0]),
	.add_fcc_out			(add_fcc_out[1:0]),
	.se_add_exp     (se_add_exp_buf2),
	.se_add_frac    (se_add_frac_buf2),
  .si             (scan_manual_1),
  .so             (scan_manual_2)
);
fpu_mul fpu_mul (
	.inq_op				(inq_op_mul_buf1[7:0]),
	.inq_rnd_mode			(inq_rnd_mode_mul_buf1[1:0]),
	.inq_id				(inq_id_mul_buf1[4:0]),
	.inq_in1			(inq_in1_mul_buf1[63:0]),
	.inq_in1_53_0_neq_0		(inq_in1_53_0_neq_0),
	.inq_in1_50_0_neq_0		(inq_in1_50_0_neq_0_mul_buf1),
	.inq_in1_53_32_neq_0		(inq_in1_53_32_neq_0_mul_buf1),
	.inq_in1_exp_eq_0		(inq_in1_exp_eq_0_mul_buf1),
	.inq_in1_exp_neq_ffs		(inq_in1_exp_neq_ffs_mul_buf1),
	.inq_in2			(inq_in2_mul_buf1[63:0]),
	.inq_in2_53_0_neq_0		(inq_in2_53_0_neq_0),
	.inq_in2_50_0_neq_0		(inq_in2_50_0_neq_0_mul_buf1),
	.inq_in2_53_32_neq_0		(inq_in2_53_32_neq_0_mul_buf1),
	.inq_in2_exp_eq_0		(inq_in2_exp_eq_0_mul_buf1),
	.inq_in2_exp_neq_ffs		(inq_in2_exp_neq_ffs_mul_buf1),
	.inq_mul			(inq_mul),
	.mul_dest_rdy			(mul_dest_rdy),
	.mul_dest_rdya			(mul_dest_rdy),
	.fmul_clken_l			(fmul_clken_l),
	.fmul_clken_l_buf1			(fmul_clken_l_buf1),
	.arst_l				(arst_l_mul_buf2),
	.grst_l				(fpu_grst_l_mul_buf1),
	.rclk				(rclk),
	.mul_pipe_active                (mul_pipe_active),
	.m1stg_step			(m1stg_step),
	.m6stg_fmul_in			(m6stg_fmul_in),
	.m6stg_id_in			(m6stg_id_in[9:0]),
	.mul_exc_out			(mul_exc_out[4:0]),
	.m6stg_fmul_dbl_dst		(m6stg_fmul_dbl_dst),
	.m6stg_fmuls			(m6stg_fmuls),
	.mul_sign_out			(mul_sign_out),
	.mul_exp_out			(mul_exp_out[10:0]),
	.mul_frac_out			(mul_frac_out[51:0]),
	.se_mul           (se_mul_buf4),
	.se_mul64 (se_mul64_buf2),
  .si              (scan_manual_2),
  .so              (scan_manual_3)
);
fpu_div fpu_div (
	.inq_op				(inq_op_div_buf1[7:0]),
	.inq_rnd_mode			(inq_rnd_mode_div_buf1[1:0]),
	.inq_id				(inq_id_div_buf1[4:0]),
	.inq_in1			(inq_in1_div_buf1[63:0]),
	.inq_in1_53_0_neq_0		(inq_in1_53_0_neq_0_div_buf1),
	.inq_in1_50_0_neq_0		(inq_in1_50_0_neq_0_div_buf1),
	.inq_in1_53_32_neq_0		(inq_in1_53_32_neq_0_div_buf1),
	.inq_in1_exp_eq_0		(inq_in1_exp_eq_0_div_buf1),
	.inq_in1_exp_neq_ffs		(inq_in1_exp_neq_ffs_div_buf1),
	.inq_in2			(inq_in2_div_buf1[63:0]),
	.inq_in2_53_0_neq_0		(inq_in2_53_0_neq_0_div_buf1),
	.inq_in2_50_0_neq_0		(inq_in2_50_0_neq_0_div_buf1),
	.inq_in2_53_32_neq_0		(inq_in2_53_32_neq_0_div_buf1),
	.inq_in2_exp_eq_0		(inq_in2_exp_eq_0_div_buf1),
	.inq_in2_exp_neq_ffs		(inq_in2_exp_neq_ffs_div_buf1),
	.inq_div			(inq_div),
	.div_dest_rdy			(div_dest_rdy),
  .fdiv_clken_l			(fdiv_clken_l_div_frac_buf1),
  .fdiv_clken_l_div_exp_buf1 (fdiv_clken_l_div_exp_buf1),
	.arst_l				(arst_l_div_buf2),
	.grst_l				(fpu_grst_l),
	.rclk				(rclk),
	.div_pipe_active                (div_pipe_active),
	.d1stg_step			(d1stg_step),
	.d8stg_fdiv_in			(d8stg_fdiv_in),
	.div_id_out_in			(div_id_out_in[9:0]),
	.div_exc_out			(div_exc_out[4:0]),
	.d8stg_fdivd			(d8stg_fdivd),
	.d8stg_fdivs			(d8stg_fdivs),
	.div_sign_out			(div_sign_out),
	.div_exp_outa			(div_exp_out[10:0]),
	.div_frac_outa			(div_frac_out[51:0]),
	.se              (se_div_buf5),
  .si              (scan_manual_3),
  .so              (scan_manual_4)
);
fpu_out fpu_out (
	.d8stg_fdiv_in			(d8stg_fdiv_in),
	.m6stg_fmul_in			(m6stg_fmul_in),
	.a6stg_fadd_in			(a6stg_fadd_in),
	.div_id_out_in			(div_id_out_in[9:0]),
	.m6stg_id_in			(m6stg_id_in[9:0]),
	.add_id_out_in			(add_id_out_in[9:0]),
	.div_exc_out			(div_exc_out[4:0]),
	.d8stg_fdivd			(d8stg_fdivd),
	.d8stg_fdivs			(d8stg_fdivs),
	.div_sign_out			(div_sign_out),
	.div_exp_out			(div_exp_out[10:0]),
	.div_frac_out			(div_frac_out[51:0]),
	.mul_exc_out			(mul_exc_out[4:0]),
	.m6stg_fmul_dbl_dst		(m6stg_fmul_dbl_dst),
	.m6stg_fmuls			(m6stg_fmuls),
	.mul_sign_out			(mul_sign_out),
	.mul_exp_out			(mul_exp_out[10:0]),
	.mul_frac_out			(mul_frac_out[51:0]),
	.add_exc_out			(add_exc_out[4:0]),
	.a6stg_fcmpop			(a6stg_fcmpop),
	.add_cc_out			(add_cc_out[1:0]),
	.add_fcc_out			(add_fcc_out[1:0]),
	.a6stg_dbl_dst			(a6stg_dbl_dst),
	.a6stg_sng_dst			(a6stg_sng_dst),
	.a6stg_long_dst			(a6stg_long_dst),
	.a6stg_int_dst			(a6stg_int_dst),
	.add_sign_out			(add_sign_out),
	.add_exp_out			(add_exp_out[10:0]),
	.add_frac_out			(add_frac_out[63:0]),
	.arst_l				(arst_l_out_buf3),
	.grst_l				(fpu_grst_l_add_buf3),
	.rclk				(rclk),
	.fp_cpx_req_cq			(fp_cpx_req_cq_unbuf[7:0]),
	.add_dest_rdy			(add_dest_rdy),
	.mul_dest_rdy			(mul_dest_rdy),
	.div_dest_rdy			(div_dest_rdy),
	.fp_cpx_data_ca			(fp_cpx_data_ca_unbuf[144:0]),
	.se               (se_out_buf2),
  .si           (scan_manual_4),
  .so           (scan_manual_5)
);
assign se = 1'b0;
assign sehold = 1'b0;
assign rst_tri_en = 1'b0;
assign rclk = gclk;
assign fpu_grst_l = grst_l;
fpu_rptr_groups fpu_rptr_groups (
	.inq_in1 (inq_in1[63:0]),
	.inq_in2 (inq_in2[63:0]),
	.inq_id (inq_id[4:0]),
	.inq_op (inq_op[7:0]),
	.inq_rnd_mode (inq_rnd_mode[1:0]),
	.inq_in1_50_0_neq_0 (inq_in1_50_0_neq_0),
	.inq_in1_53_0_neq_0 (inq_in1_53_0_neq_0),
	.inq_in1_53_32_neq_0 (inq_in1_53_32_neq_0),
	.inq_in1_exp_eq_0 (inq_in1_exp_eq_0),
	.inq_in1_exp_neq_ffs (inq_in1_exp_neq_ffs),
	.inq_in2_50_0_neq_0 (inq_in2_50_0_neq_0),
	.inq_in2_53_0_neq_0 (inq_in2_53_0_neq_0),
	.inq_in2_53_32_neq_0 (inq_in2_53_32_neq_0),
	.inq_in2_exp_eq_0 (inq_in2_exp_eq_0),
	.inq_in2_exp_neq_ffs (inq_in2_exp_neq_ffs),
	.ctu_tst_macrotest (ctu_tst_macrotest),
	.ctu_tst_pre_grst_l (ctu_tst_pre_grst_l),
	.ctu_tst_scan_disable (ctu_tst_scan_disable),
	.ctu_tst_scanmode (ctu_tst_scanmode),
	.ctu_tst_short_chain (ctu_tst_short_chain),
	.global_shift_enable (global_shift_enable),
	.grst_l (grst_l),
	.cluster_cken (cluster_cken),
	.se (se),
	.arst_l (arst_l),
	.fpu_grst_l (fpu_grst_l),
	.fmul_clken_l (fmul_clken_l),
	.fdiv_clken_l (fdiv_clken_l),
	.scan_manual_6 (),
	
	.si (si),
	.so_unbuf (so_unbuf),
	.pcx_fpio_data_px2 (pcx_fpio_data_px2[123:0]),
	.pcx_fpio_data_rdy_px2 (pcx_fpio_data_rdy_px2),
	.fp_cpx_data_ca (fp_cpx_data_ca_unbuf[144:0]),
	.fp_cpx_req_cq (fp_cpx_req_cq_unbuf[7:0]),
	.inq_sram_din_unbuf ({fp_id_in[4:0],
		fp_rnd_mode_in[1:0],
		fp_fcc_in[1:0],
		fp_op_in[7:0],
		fp_src1_in[68:0],
		fp_src2_in[68:0], 1'b0}),
	.inq_in1_add_buf1 (inq_in1_add_buf1[63:0]),
	.inq_in1_mul_buf1 (inq_in1_mul_buf1[63:0]),
	.inq_in1_div_buf1 (inq_in1_div_buf1[63:0]),
	.inq_in2_add_buf1 (inq_in2_add_buf1[63:0]),
	.inq_in2_mul_buf1 (inq_in2_mul_buf1[63:0]),
	.inq_in2_div_buf1 (inq_in2_div_buf1[63:0]),
	.inq_id_add_buf1 (inq_id_add_buf1[4:0]),
	.inq_id_div_buf1 (inq_id_div_buf1[4:0]),
	.inq_id_mul_buf1 (inq_id_mul_buf1[4:0]),
	.inq_op_add_buf1 (inq_op_add_buf1[7:0]),
	.inq_op_mul_buf1 (inq_op_mul_buf1[7:0]),
	.inq_op_div_buf1 (inq_op_div_buf1[7:0]),
	.inq_rnd_mode_add_buf1 (inq_rnd_mode_add_buf1[1:0]),
	.inq_rnd_mode_mul_buf1 (inq_rnd_mode_mul_buf1[1:0]),
	.inq_rnd_mode_div_buf1 (inq_rnd_mode_div_buf1[1:0]),
	.inq_in1_50_0_neq_0_add_buf1 (inq_in1_50_0_neq_0_add_buf1),
	.inq_in1_50_0_neq_0_mul_buf1 (inq_in1_50_0_neq_0_mul_buf1),
	.inq_in1_50_0_neq_0_div_buf1 (inq_in1_50_0_neq_0_div_buf1),
	.inq_in1_53_0_neq_0_add_buf1 (inq_in1_53_0_neq_0_add_buf1),
	.inq_in1_53_0_neq_0_mul_buf1 (inq_in1_53_0_neq_0_mul_buf1),
	.inq_in1_53_0_neq_0_div_buf1 (inq_in1_53_0_neq_0_div_buf1),
	.inq_in1_53_32_neq_0_add_buf1 (inq_in1_53_32_neq_0_add_buf1),
	.inq_in1_53_32_neq_0_mul_buf1 (inq_in1_53_32_neq_0_mul_buf1),
	.inq_in1_53_32_neq_0_div_buf1 (inq_in1_53_32_neq_0_div_buf1),
	.inq_in1_exp_eq_0_add_buf1 (inq_in1_exp_eq_0_add_buf1),
	.inq_in1_exp_eq_0_mul_buf1 (inq_in1_exp_eq_0_mul_buf1),
	.inq_in1_exp_eq_0_div_buf1 (inq_in1_exp_eq_0_div_buf1),
	.inq_in1_exp_neq_ffs_add_buf1 (inq_in1_exp_neq_ffs_add_buf1),
	.inq_in1_exp_neq_ffs_mul_buf1 (inq_in1_exp_neq_ffs_mul_buf1),
	.inq_in1_exp_neq_ffs_div_buf1 (inq_in1_exp_neq_ffs_div_buf1),
	.inq_in2_50_0_neq_0_add_buf1 (inq_in2_50_0_neq_0_add_buf1),
	.inq_in2_50_0_neq_0_mul_buf1 (inq_in2_50_0_neq_0_mul_buf1),
	.inq_in2_50_0_neq_0_div_buf1 (inq_in2_50_0_neq_0_div_buf1),
	.inq_in2_53_0_neq_0_add_buf1 (inq_in2_53_0_neq_0_add_buf1),
	.inq_in2_53_0_neq_0_mul_buf1 (inq_in2_53_0_neq_0_mul_buf1),
	.inq_in2_53_0_neq_0_div_buf1 (inq_in2_53_0_neq_0_div_buf1),
	.inq_in2_53_32_neq_0_add_buf1 (inq_in2_53_32_neq_0_add_buf1),
	.inq_in2_53_32_neq_0_mul_buf1 (inq_in2_53_32_neq_0_mul_buf1),
	.inq_in2_53_32_neq_0_div_buf1 (inq_in2_53_32_neq_0_div_buf1),
	.inq_in2_exp_eq_0_add_buf1 (inq_in2_exp_eq_0_add_buf1),
	.inq_in2_exp_eq_0_mul_buf1 (inq_in2_exp_eq_0_mul_buf1),
	.inq_in2_exp_eq_0_div_buf1 (inq_in2_exp_eq_0_div_buf1),
	.inq_in2_exp_neq_ffs_add_buf1 (inq_in2_exp_neq_ffs_add_buf1),
	.inq_in2_exp_neq_ffs_mul_buf1 (inq_in2_exp_neq_ffs_mul_buf1),
	.inq_in2_exp_neq_ffs_div_buf1 (inq_in2_exp_neq_ffs_div_buf1),
	.ctu_tst_macrotest_buf1 (ctu_tst_macrotest_buf1),
	.ctu_tst_pre_grst_l_buf1 (ctu_tst_pre_grst_l_buf1),
	.ctu_tst_scan_disable_buf1 (ctu_tst_scan_disable_buf1),
	.ctu_tst_scanmode_buf1 (ctu_tst_scanmode_buf1),
	.ctu_tst_short_chain_buf1 (ctu_tst_short_chain_buf1),
	.global_shift_enable_buf1 (global_shift_enable_buf1),
	.grst_l_buf1 (grst_l_buf1),
	.cluster_cken_buf1 (cluster_cken_buf1),
	.se_add_exp_buf2 (se_add_exp_buf2),
	.se_add_frac_buf2 (se_add_frac_buf2),
	.se_out_buf2 (se_out_buf2),
	.se_mul64_buf2 (se_mul64_buf2),
	.se_cluster_header_buf2 (se_cluster_header_buf2),
	.se_in_buf3 (se_in_buf3),
	.se_mul_buf4 (se_mul_buf4),
	.se_div_buf5 (se_div_buf5),
	.arst_l_div_buf2 (arst_l_div_buf2),
	.arst_l_mul_buf2 (arst_l_mul_buf2),
	.arst_l_cluster_header_buf2 (arst_l_cluster_header_buf2),
	.arst_l_in_buf3 (arst_l_in_buf3),
	.arst_l_out_buf3 (arst_l_out_buf3),
	.arst_l_add_buf4 (arst_l_add_buf4),
	.fpu_grst_l_mul_buf1 (fpu_grst_l_mul_buf1),
	.fpu_grst_l_in_buf2 (fpu_grst_l_in_buf2),
	.fpu_grst_l_add_buf3 (fpu_grst_l_add_buf3),
	.fmul_clken_l_buf1 (fmul_clken_l_buf1),
	.fdiv_clken_l_div_exp_buf1 (fdiv_clken_l_div_exp_buf1),
	.fdiv_clken_l_div_frac_buf1 (fdiv_clken_l_div_frac_buf1),
	.scan_manual_6_buf1 (scan_manual_6_buf1),
	.si_buf1 (si_buf1),
	.so (so),
	.pcx_fpio_data_px2_buf1 (pcx_fpio_data_px2_buf1[123:0]),
	.pcx_fpio_data_rdy_px2_buf1 (pcx_fpio_data_rdy_px2_buf1),
	.fp_cpx_data_ca_buf1 (fp_cpx_data_ca[144:0]),
	.fp_cpx_req_cq_buf1 (fp_cpx_req_cq[7:0]),
	.inq_sram_din_buf1 (inq_sram_din_buf1[155:0])
);
endmodule
module fpu_add (
	inq_op,
	inq_rnd_mode,
	inq_id,
	inq_fcc,
	inq_in1,
	inq_in1_50_0_neq_0,
	inq_in1_53_32_neq_0,
	inq_in1_exp_eq_0,
	inq_in1_exp_neq_ffs,
	inq_in2,
	inq_in2_50_0_neq_0,
	inq_in2_53_32_neq_0,
	inq_in2_exp_eq_0,
	inq_in2_exp_neq_ffs,
	inq_add,
	add_dest_rdy,
	fadd_clken_l,
	arst_l,
	grst_l,
	rclk,
	add_pipe_active,	
	a1stg_step,
	a6stg_fadd_in,
	add_id_out_in,
	a6stg_fcmpop,
	add_exc_out,
	a6stg_dbl_dst,
	a6stg_sng_dst,
	a6stg_long_dst,
	a6stg_int_dst,
	add_sign_out,
	add_exp_out,
	add_frac_out,
	add_cc_out,
	add_fcc_out,
	se_add_exp,
	se_add_frac,
	si,
	so
);
input [7:0]	inq_op;			
input [1:0]	inq_rnd_mode;		
input [4:0]	inq_id;			
input [1:0]	inq_fcc;		
input [63:0]	inq_in1;		
input		inq_in1_50_0_neq_0;	
input		inq_in1_53_32_neq_0;	
input		inq_in1_exp_eq_0;	
input		inq_in1_exp_neq_ffs;	
input [63:0]	inq_in2;		
input		inq_in2_50_0_neq_0;	
input		inq_in2_53_32_neq_0;	
input		inq_in2_exp_eq_0;	
input		inq_in2_exp_neq_ffs;	
input		inq_add;		
input		add_dest_rdy;		
input		fadd_clken_l;           
input		arst_l;			
input		grst_l;			
input		rclk;			
output		add_pipe_active;        
output		a1stg_step;		
output		a6stg_fadd_in;		
output [9:0]    add_id_out_in;		
output		a6stg_fcmpop;		
output [4:0]	add_exc_out;		
output		a6stg_dbl_dst;		
output		a6stg_sng_dst;		
output		a6stg_long_dst;		
output		a6stg_int_dst;		
output		add_sign_out;		
output [10:0]	add_exp_out;		
output [63:0]	add_frac_out;		
output [1:0]	add_cc_out;		
output [1:0]	add_fcc_out;		
input           se_add_exp;     
input           se_add_frac;    
input           si;                     
output          so;                     
wire		a1stg_denorm_sng_in1;	
wire		a1stg_denorm_dbl_in1;	
wire		a1stg_denorm_sng_in2;	
wire		a1stg_denorm_dbl_in2;	
wire		a1stg_norm_sng_in1;	
wire		a1stg_norm_dbl_in1;	
wire		a1stg_norm_sng_in2;	
wire		a1stg_norm_dbl_in2;	
wire		a1stg_step;		
wire		a1stg_stepa;		
wire		a1stg_sngop;		
wire		a1stg_intlngop;		
wire		a1stg_fsdtoix;		
wire		a1stg_fstod;		
wire		a1stg_fstoi;		
wire		a1stg_fstox;		
wire		a1stg_fdtoi;		
wire		a1stg_fdtox;		
wire		a1stg_faddsubs;		
wire		a1stg_faddsubd;		
wire		a1stg_fdtos;		
wire		a2stg_faddsubop;	
wire		a2stg_fsdtoix_fdtos;	
wire		a2stg_fitos;		
wire		a2stg_fitod;		
wire		a2stg_fxtos;		
wire		a2stg_fxtod;		
wire		a3stg_faddsubop;	
wire [1:0]	a3stg_faddsubopa;	
wire		a4stg_dblop;		
wire		a6stg_fadd_in;		
wire [9:0]	add_id_out_in;		
wire [1:0]	add_fcc_out;		
wire		a6stg_dbl_dst;		
wire		a6stg_sng_dst;		
wire		a6stg_long_dst;		
wire		a6stg_int_dst;		
wire		a6stg_fcmpop;		
wire		a6stg_step;		
wire		a3stg_sub_in;		
wire		add_sign_out;		
wire [1:0]	add_cc_out;		
wire		a4stg_in_of;		
wire [4:0]	add_exc_out;		
wire		a2stg_frac1_in_frac1;	
wire		a2stg_frac1_in_frac2;	
wire		a1stg_2nan_in_inv;	
wire		a1stg_faddsubop_inv;	
wire		a2stg_frac1_in_qnan;	
wire		a2stg_frac1_in_nv;	
wire		a2stg_frac1_in_nv_dbl;	
wire		a2stg_frac2_in_frac1;	
wire		a2stg_frac2_in_qnan;	
wire [5:0]	a2stg_shr_cnt_in;	
wire 		a2stg_shr_cnt_5_inv_in; 
wire		a2stg_shr_frac2_shr_int; 
wire		a2stg_shr_frac2_shr_dbl; 
wire		a2stg_shr_frac2_shr_sng; 
wire		a2stg_shr_frac2_max;	
wire		a2stg_sub_step;		
wire		a2stg_fracadd_frac2_inv_in; 
wire		a2stg_fracadd_frac2_inv_shr1_in; 
wire		a2stg_fracadd_frac2;	
wire		a2stg_fracadd_cin_in;	
wire		a3stg_exp_7ff;		
wire		a3stg_exp_ff;		
wire		a3stg_exp_add;		
wire		a2stg_expdec_neq_0;	
wire		a3stg_exp10_0_eq0;	
wire		a3stg_exp10_1_eq0;	
wire		a3stg_fdtos_inv;	
wire		a4stg_fixtos_fxtod_inv;	
wire		a4stg_rnd_frac_add_inv;	
wire [9:0]	a4stg_shl_cnt_in;	
wire		a4stg_rnd_sng;		
wire		a4stg_rnd_dbl;		
wire		add_frac_out_rndadd;	
wire		add_frac_out_rnd_frac;	
wire		add_frac_out_shl;	
wire		a4stg_to_0;		
wire		add_exp_out_expinc;	
wire		add_exp_out_exp;	
wire		add_exp_out_exp1;	
wire		add_exp_out_expadd;	
wire		a4stg_to_0_inv;		
wire            add_pipe_active;        
wire        	a1stg_expadd3_11;	
wire [11:0]	a1stg_expadd1_11_0;	
wire [10:0]	a1stg_expadd4_inv;	
wire [5:0]	a1stg_expadd2_5_0;	
wire [11:0]	a2stg_exp;		
wire [12:0]	a2stg_expadd;		
wire [10:0]	a3stg_exp_10_0;		
wire [11:0]	a4stg_exp_11_0;		
wire [10:0]	add_exp_out;		
wire		a1stg_in2_neq_in1_frac;	
wire		a1stg_in2_gt_in1_frac;	
wire		a1stg_in2_eq_in1_exp;	
wire		a2stg_frac2_63;		
wire		a2stg_frac2hi_neq_0;	
wire		a2stg_frac2lo_neq_0;	
wire		a3stg_fsdtoix_nx;	
wire		a3stg_fsdtoi_nx;	
wire		a3stg_denorm;		
wire		a3stg_denorm_inv;	
wire [5:0]	a3stg_lead0;		
wire		a4stg_round;		
wire [5:0]	a4stg_shl_cnt;		
wire		a4stg_denorm_inv;	
wire		a3stg_inc_exp_inv;	
wire		a3stg_same_exp_inv;	
wire		a3stg_dec_exp_inv;	
wire		a4stg_rnd_frac_40;	
wire		a4stg_rnd_frac_39;	
wire		a4stg_rnd_frac_11;	
wire		a4stg_rnd_frac_10;	
wire		a4stg_rndadd_cout;	
wire		a4stg_frac_9_0_nx;	
wire		a4stg_frac_dbl_nx;	
wire		a4stg_frac_38_0_nx;	
wire		a4stg_frac_sng_nx;	
wire		a4stg_frac_neq_0;	
wire		a4stg_shl_data_neq_0;	
wire		add_of_out_cout;	
wire [63:0]	add_frac_out;		
wire        scan_out_fpu_add_ctl;
wire        scan_out_fpu_add_exp_dp;
fpu_add_ctl fpu_add_ctl (
	.inq_in1_51			(inq_in1[51]),
	.inq_in1_54			(inq_in1[54]),
	.inq_in1_63			(inq_in1[63]),
	.inq_in1_50_0_neq_0		(inq_in1_50_0_neq_0),
	.inq_in1_53_32_neq_0		(inq_in1_53_32_neq_0),
	.inq_in1_exp_eq_0		(inq_in1_exp_eq_0),
	.inq_in1_exp_neq_ffs		(inq_in1_exp_neq_ffs),
	.inq_in2_51			(inq_in2[51]),
	.inq_in2_54			(inq_in2[54]),
	.inq_in2_63			(inq_in2[63]),
	.inq_in2_50_0_neq_0		(inq_in2_50_0_neq_0),
	.inq_in2_53_32_neq_0		(inq_in2_53_32_neq_0),
	.inq_in2_exp_eq_0		(inq_in2_exp_eq_0),
	.inq_in2_exp_neq_ffs		(inq_in2_exp_neq_ffs),
	.inq_op				(inq_op[7:0]),
	.inq_rnd_mode			(inq_rnd_mode[1:0]),
	.inq_id				(inq_id[4:0]),
	.inq_fcc			(inq_fcc[1:0]),
	.inq_add			(inq_add),
	.add_dest_rdy			(add_dest_rdy),
	.a1stg_in2_neq_in1_frac		(a1stg_in2_neq_in1_frac),
	.a1stg_in2_gt_in1_frac		(a1stg_in2_gt_in1_frac),
	.a1stg_in2_eq_in1_exp		(a1stg_in2_eq_in1_exp),
	.a1stg_expadd1			(a1stg_expadd1_11_0[11:0]),
	.a2stg_expadd			(a2stg_expadd[11:0]),
	.a2stg_frac2hi_neq_0		(a2stg_frac2hi_neq_0),
	.a2stg_frac2lo_neq_0		(a2stg_frac2lo_neq_0),
	.a2stg_exp			(a2stg_exp[11:0]),
	.a3stg_fsdtoix_nx		(a3stg_fsdtoix_nx),
	.a3stg_fsdtoi_nx		(a3stg_fsdtoi_nx),
	.a2stg_frac2_63			(a2stg_frac2_63),
	.a4stg_exp			(a4stg_exp_11_0[11:0]),
	.add_of_out_cout		(add_of_out_cout),
	.a4stg_frac_neq_0		(a4stg_frac_neq_0),
	.a4stg_shl_data_neq_0		(a4stg_shl_data_neq_0),
	.a4stg_frac_dbl_nx		(a4stg_frac_dbl_nx),
	.a4stg_frac_sng_nx		(a4stg_frac_sng_nx),
	.a1stg_expadd2			(a1stg_expadd2_5_0[5:0]),
	.a1stg_expadd4_inv		(a1stg_expadd4_inv[10:0]),
	.a3stg_denorm			(a3stg_denorm),
	.a3stg_denorm_inv		(a3stg_denorm_inv),
	.a4stg_denorm_inv		(a4stg_denorm_inv),
	.a3stg_exp			(a3stg_exp_10_0[10:0]),
	.a4stg_round			(a4stg_round),
	.a3stg_lead0			(a3stg_lead0[5:0]),
	.a4stg_rnd_frac_40		(a4stg_rnd_frac_40),
	.a4stg_rnd_frac_39		(a4stg_rnd_frac_39),
	.a4stg_rnd_frac_11		(a4stg_rnd_frac_11),
	.a4stg_rnd_frac_10		(a4stg_rnd_frac_10),
	.a4stg_frac_38_0_nx		(a4stg_frac_38_0_nx),
	.a4stg_frac_9_0_nx		(a4stg_frac_9_0_nx),
	.arst_l				(arst_l),
	.grst_l				(grst_l),
	.rclk			(rclk),
	.add_pipe_active                (add_pipe_active),
	.a1stg_denorm_sng_in1		(a1stg_denorm_sng_in1),
	.a1stg_denorm_dbl_in1		(a1stg_denorm_dbl_in1),
	.a1stg_denorm_sng_in2		(a1stg_denorm_sng_in2),
	.a1stg_denorm_dbl_in2		(a1stg_denorm_dbl_in2),
	.a1stg_norm_sng_in1		(a1stg_norm_sng_in1),
	.a1stg_norm_dbl_in1		(a1stg_norm_dbl_in1),
	.a1stg_norm_sng_in2		(a1stg_norm_sng_in2),
	.a1stg_norm_dbl_in2		(a1stg_norm_dbl_in2),
	.a1stg_step			(a1stg_step),
	.a1stg_stepa			(a1stg_stepa),
	.a1stg_sngop			(a1stg_sngop),
	.a1stg_intlngop			(a1stg_intlngop),
	.a1stg_fsdtoix			(a1stg_fsdtoix),
	.a1stg_fstod			(a1stg_fstod),
	.a1stg_fstoi			(a1stg_fstoi),
	.a1stg_fstox			(a1stg_fstox),
	.a1stg_fdtoi			(a1stg_fdtoi),
	.a1stg_fdtox			(a1stg_fdtox),
	.a1stg_faddsubs			(a1stg_faddsubs),
	.a1stg_faddsubd			(a1stg_faddsubd),
	.a1stg_fdtos			(a1stg_fdtos),
	.a2stg_faddsubop		(a2stg_faddsubop),
	.a2stg_fsdtoix_fdtos		(a2stg_fsdtoix_fdtos),
	.a2stg_fitos			(a2stg_fitos),
	.a2stg_fitod			(a2stg_fitod),
	.a2stg_fxtos			(a2stg_fxtos),
	.a2stg_fxtod			(a2stg_fxtod),
	.a3stg_faddsubop		(a3stg_faddsubop),
	.a3stg_faddsubopa		(a3stg_faddsubopa[1:0]),
	.a4stg_dblop			(a4stg_dblop),
	.a6stg_fadd_in			(a6stg_fadd_in),
	.add_id_out_in			(add_id_out_in[9:0]),
	.add_fcc_out			(add_fcc_out[1:0]),
	.a6stg_dbl_dst			(a6stg_dbl_dst),
	.a6stg_sng_dst			(a6stg_sng_dst),
	.a6stg_long_dst			(a6stg_long_dst),
	.a6stg_int_dst			(a6stg_int_dst),
	.a6stg_fcmpop			(a6stg_fcmpop),
	.a6stg_step			(a6stg_step),
	.a3stg_sub_in			(a3stg_sub_in),
	.add_sign_out			(add_sign_out),
	.add_cc_out			(add_cc_out[1:0]),
	.a4stg_in_of			(a4stg_in_of),
	.add_exc_out			(add_exc_out[4:0]),
	.a2stg_frac1_in_frac1		(a2stg_frac1_in_frac1),
	.a2stg_frac1_in_frac2		(a2stg_frac1_in_frac2),
	.a1stg_2nan_in_inv		(a1stg_2nan_in_inv),
	.a1stg_faddsubop_inv		(a1stg_faddsubop_inv),
	.a2stg_frac1_in_qnan		(a2stg_frac1_in_qnan),
	.a2stg_frac1_in_nv		(a2stg_frac1_in_nv),
	.a2stg_frac1_in_nv_dbl		(a2stg_frac1_in_nv_dbl),
	.a2stg_frac2_in_frac1		(a2stg_frac2_in_frac1),
	.a2stg_frac2_in_qnan		(a2stg_frac2_in_qnan),
	.a2stg_shr_cnt_in		(a2stg_shr_cnt_in[5:0]),
	.a2stg_shr_cnt_5_inv_in   (a2stg_shr_cnt_5_inv_in),
	.a2stg_shr_frac2_shr_int	(a2stg_shr_frac2_shr_int),
	.a2stg_shr_frac2_shr_dbl	(a2stg_shr_frac2_shr_dbl),
	.a2stg_shr_frac2_shr_sng	(a2stg_shr_frac2_shr_sng),
	.a2stg_shr_frac2_max		(a2stg_shr_frac2_max),
	.a2stg_sub_step			(a2stg_sub_step),
	.a2stg_fracadd_frac2_inv_in	(a2stg_fracadd_frac2_inv_in),
	.a2stg_fracadd_frac2_inv_shr1_in (a2stg_fracadd_frac2_inv_shr1_in),
	.a2stg_fracadd_frac2		(a2stg_fracadd_frac2),
	.a2stg_fracadd_cin_in		(a2stg_fracadd_cin_in),
	.a3stg_exp_7ff			(a3stg_exp_7ff),
	.a3stg_exp_ff			(a3stg_exp_ff),
	.a3stg_exp_add			(a3stg_exp_add),
	.a2stg_expdec_neq_0		(a2stg_expdec_neq_0),
	.a3stg_exp10_0_eq0		(a3stg_exp10_0_eq0),
	.a3stg_exp10_1_eq0		(a3stg_exp10_1_eq0),
	.a3stg_fdtos_inv		(a3stg_fdtos_inv),
	.a4stg_fixtos_fxtod_inv		(a4stg_fixtos_fxtod_inv),
	.a4stg_rnd_frac_add_inv		(a4stg_rnd_frac_add_inv),
	.a4stg_shl_cnt_in		(a4stg_shl_cnt_in[9:0]),
	.a4stg_rnd_sng			(a4stg_rnd_sng),
	.a4stg_rnd_dbl			(a4stg_rnd_dbl),
	.add_frac_out_rndadd		(add_frac_out_rndadd),
	.add_frac_out_rnd_frac		(add_frac_out_rnd_frac),
	.add_frac_out_shl		(add_frac_out_shl),
	.a4stg_to_0			(a4stg_to_0),
	.add_exp_out_expinc		(add_exp_out_expinc),
	.add_exp_out_exp		(add_exp_out_exp),
	.add_exp_out_exp1		(add_exp_out_exp1),
	.add_exp_out_expadd		(add_exp_out_expadd),
	.a4stg_to_0_inv			(a4stg_to_0_inv),
	.se				(se_add_exp),
	.si				(si),
	.so				(scan_out_fpu_add_ctl)
);
fpu_add_exp_dp fpu_add_exp_dp (
	.inq_in1			(inq_in1[62:52]),
	.inq_in2			(inq_in2[62:52]),
	.inq_op				(inq_op[1:0]),
	.inq_op_7			(inq_op[7]),
	.a1stg_step			(a1stg_stepa),
	.a1stg_faddsubd			(a1stg_faddsubd),
	.a1stg_faddsubs			(a1stg_faddsubs),
	.a1stg_fsdtoix			(a1stg_fsdtoix),
	.a6stg_step			(a6stg_step),
	.a1stg_fstod			(a1stg_fstod),
	.a1stg_fdtos			(a1stg_fdtos),
	.a1stg_fstoi			(a1stg_fstoi),
	.a1stg_fstox			(a1stg_fstox),
	.a1stg_fdtoi			(a1stg_fdtoi),
	.a1stg_fdtox			(a1stg_fdtox),
	.a2stg_fsdtoix_fdtos		(a2stg_fsdtoix_fdtos),
	.a2stg_faddsubop		(a2stg_faddsubop),
	.a2stg_fitos			(a2stg_fitos),
	.a2stg_fitod			(a2stg_fitod),
	.a2stg_fxtos			(a2stg_fxtos),
	.a2stg_fxtod			(a2stg_fxtod),
	.a3stg_exp_7ff			(a3stg_exp_7ff),
	.a3stg_exp_ff			(a3stg_exp_ff),
	.a3stg_exp_add			(a3stg_exp_add),
	.a3stg_inc_exp_inv		(a3stg_inc_exp_inv),
	.a3stg_same_exp_inv		(a3stg_same_exp_inv),
	.a3stg_dec_exp_inv		(a3stg_dec_exp_inv),
	.a3stg_faddsubop		(a3stg_faddsubop),
	.a3stg_fdtos_inv		(a3stg_fdtos_inv),
	.a4stg_fixtos_fxtod_inv		(a4stg_fixtos_fxtod_inv),
	.a4stg_shl_cnt			(a4stg_shl_cnt[5:0]),
	.a4stg_denorm_inv		(a4stg_denorm_inv),
	.a4stg_rndadd_cout		(a4stg_rndadd_cout),
	.add_exp_out_expinc		(add_exp_out_expinc),
	.add_exp_out_exp		(add_exp_out_exp),
	.add_exp_out_exp1		(add_exp_out_exp1),
	.a4stg_in_of			(a4stg_in_of),
	.add_exp_out_expadd		(add_exp_out_expadd),
	.a4stg_dblop			(a4stg_dblop),
	.a4stg_to_0_inv			(a4stg_to_0_inv),
	.fadd_clken_l			(fadd_clken_l),
	.rclk			(rclk),
	.a1stg_expadd3_11		(a1stg_expadd3_11),
	.a1stg_expadd1_11_0		(a1stg_expadd1_11_0[11:0]),
	.a1stg_expadd4_inv		(a1stg_expadd4_inv[10:0]),
	.a1stg_expadd2_5_0		(a1stg_expadd2_5_0[5:0]),
	.a2stg_exp			(a2stg_exp[11:0]),
	.a2stg_expadd			(a2stg_expadd[12:0]),
	.a3stg_exp_10_0			(a3stg_exp_10_0[10:0]),
	.a4stg_exp_11_0			(a4stg_exp_11_0[11:0]),
	.add_exp_out			(add_exp_out[10:0]),
	.se                             (se_add_exp),
        .si                             (scan_out_fpu_add_ctl),
        .so                             (scan_out_fpu_add_exp_dp)
);
fpu_add_frac_dp fpu_add_frac_dp (
	.inq_in1			(inq_in1[62:0]),
	.inq_in2			(inq_in2[63:0]),
	.a1stg_step			(a1stg_stepa),
	.a1stg_sngop			(a1stg_sngop),
	.a1stg_expadd3_11		(a1stg_expadd3_11),
	.a1stg_norm_dbl_in1		(a1stg_norm_dbl_in1),
	.a1stg_denorm_dbl_in1		(a1stg_denorm_dbl_in1),
	.a1stg_norm_sng_in1		(a1stg_norm_sng_in1),
	.a1stg_denorm_sng_in1		(a1stg_denorm_sng_in1),
	.a1stg_norm_dbl_in2		(a1stg_norm_dbl_in2),
	.a1stg_denorm_dbl_in2		(a1stg_denorm_dbl_in2),
	.a1stg_norm_sng_in2		(a1stg_norm_sng_in2),
	.a1stg_denorm_sng_in2		(a1stg_denorm_sng_in2),
	.a1stg_intlngop			(a1stg_intlngop),
	.a2stg_frac1_in_frac1		(a2stg_frac1_in_frac1),
	.a2stg_frac1_in_frac2		(a2stg_frac1_in_frac2),
	.a1stg_2nan_in_inv		(a1stg_2nan_in_inv),
	.a1stg_faddsubop_inv		(a1stg_faddsubop_inv),
	.a2stg_frac1_in_qnan		(a2stg_frac1_in_qnan),
	.a2stg_frac1_in_nv		(a2stg_frac1_in_nv),
	.a2stg_frac1_in_nv_dbl		(a2stg_frac1_in_nv_dbl),
	.a6stg_step			(a6stg_step),
	.a2stg_frac2_in_frac1		(a2stg_frac2_in_frac1),
	.a2stg_frac2_in_qnan		(a2stg_frac2_in_qnan),
	.a2stg_shr_cnt_in		(a2stg_shr_cnt_in[5:0]),
	.a2stg_shr_cnt_5_inv_in (a2stg_shr_cnt_5_inv_in),
	.a2stg_shr_frac2_shr_int	(a2stg_shr_frac2_shr_int),
	.a2stg_shr_frac2_shr_dbl	(a2stg_shr_frac2_shr_dbl),
	.a2stg_shr_frac2_shr_sng	(a2stg_shr_frac2_shr_sng),
	.a2stg_shr_frac2_max		(a2stg_shr_frac2_max),
	.a2stg_expadd_11		(a2stg_expadd[12]),
	.a2stg_sub_step			(a2stg_sub_step),
	.a2stg_fracadd_frac2_inv_in	(a2stg_fracadd_frac2_inv_in),
	.a2stg_fracadd_frac2_inv_shr1_in (a2stg_fracadd_frac2_inv_shr1_in),
	.a2stg_fracadd_frac2		(a2stg_fracadd_frac2),
	.a2stg_fracadd_cin_in		(a2stg_fracadd_cin_in),
	.a2stg_exp			(a2stg_exp[5:0]),
	.a2stg_expdec_neq_0		(a2stg_expdec_neq_0),
	.a3stg_faddsubopa		(a3stg_faddsubopa[1:0]),
	.a3stg_sub_in			(a3stg_sub_in),
	.a3stg_exp10_0_eq0		(a3stg_exp10_0_eq0),
	.a3stg_exp10_1_eq0		(a3stg_exp10_1_eq0),
	.a3stg_exp_0			(a3stg_exp_10_0[0]),
	.a4stg_rnd_frac_add_inv		(a4stg_rnd_frac_add_inv),
	.a3stg_fdtos_inv		(a3stg_fdtos_inv),
	.a4stg_fixtos_fxtod_inv		(a4stg_fixtos_fxtod_inv),
	.a4stg_rnd_sng			(a4stg_rnd_sng),
	.a4stg_rnd_dbl			(a4stg_rnd_dbl),
	.a4stg_shl_cnt_in		(a4stg_shl_cnt_in[9:0]),
	.add_frac_out_rndadd		(add_frac_out_rndadd),
	.add_frac_out_rnd_frac		(add_frac_out_rnd_frac),
	.a4stg_in_of			(a4stg_in_of),
	.add_frac_out_shl		(add_frac_out_shl),
	.a4stg_to_0			(a4stg_to_0),
	.fadd_clken_l			(fadd_clken_l),
	.rclk			(rclk),
	.a1stg_in2_neq_in1_frac		(a1stg_in2_neq_in1_frac),
	.a1stg_in2_gt_in1_frac		(a1stg_in2_gt_in1_frac),
	.a1stg_in2_eq_in1_exp		(a1stg_in2_eq_in1_exp),
	.a2stg_frac2_63			(a2stg_frac2_63),
	.a2stg_frac2hi_neq_0		(a2stg_frac2hi_neq_0),
	.a2stg_frac2lo_neq_0		(a2stg_frac2lo_neq_0),
	.a3stg_fsdtoix_nx		(a3stg_fsdtoix_nx),
	.a3stg_fsdtoi_nx		(a3stg_fsdtoi_nx),
	.a3stg_denorm			(a3stg_denorm),
	.a3stg_denorm_inv		(a3stg_denorm_inv),
	.a3stg_lead0			(a3stg_lead0[5:0]),
	.a4stg_round			(a4stg_round),
	.a4stg_shl_cnt			(a4stg_shl_cnt[5:0]),
	.a4stg_denorm_inv		(a4stg_denorm_inv),
	.a3stg_inc_exp_inv		(a3stg_inc_exp_inv),
	.a3stg_same_exp_inv		(a3stg_same_exp_inv),
	.a3stg_dec_exp_inv		(a3stg_dec_exp_inv),
	.a4stg_rnd_frac_40		(a4stg_rnd_frac_40),
	.a4stg_rnd_frac_39		(a4stg_rnd_frac_39),
	.a4stg_rnd_frac_11		(a4stg_rnd_frac_11),
	.a4stg_rnd_frac_10		(a4stg_rnd_frac_10),
	.a4stg_rndadd_cout		(a4stg_rndadd_cout),
	.a4stg_frac_9_0_nx		(a4stg_frac_9_0_nx),
	.a4stg_frac_dbl_nx		(a4stg_frac_dbl_nx),
	.a4stg_frac_38_0_nx		(a4stg_frac_38_0_nx),
	.a4stg_frac_sng_nx		(a4stg_frac_sng_nx),
	.a4stg_frac_neq_0		(a4stg_frac_neq_0),
	.a4stg_shl_data_neq_0		(a4stg_shl_data_neq_0),
	.add_of_out_cout		(add_of_out_cout),
	.add_frac_out			(add_frac_out[63:0]),
	.se                             (se_add_frac),
        .si                             (scan_out_fpu_add_exp_dp),
        .so                             (so)
);
endmodule
module fpu_add_ctl (
	inq_in1_51,
	inq_in1_54,
	inq_in1_63,
	inq_in1_50_0_neq_0,
	inq_in1_53_32_neq_0,
	inq_in1_exp_eq_0,
	inq_in1_exp_neq_ffs,
	inq_in2_51,
	inq_in2_54,
	inq_in2_63,
	inq_in2_50_0_neq_0,
	inq_in2_53_32_neq_0,
	inq_in2_exp_eq_0,
	inq_in2_exp_neq_ffs,
	inq_op,
	inq_rnd_mode,
	inq_id,
	inq_fcc,
	inq_add,
	add_dest_rdy,
	a1stg_in2_neq_in1_frac,
	a1stg_in2_gt_in1_frac,
	a1stg_in2_eq_in1_exp,
	a1stg_expadd1,
	a2stg_expadd,
	a2stg_frac2hi_neq_0,
	a2stg_frac2lo_neq_0,
	a2stg_exp,
	a3stg_fsdtoix_nx,
	a3stg_fsdtoi_nx,
	a2stg_frac2_63,
	a4stg_exp,
	add_of_out_cout,
	a4stg_frac_neq_0,
	a4stg_shl_data_neq_0,
	a4stg_frac_dbl_nx,
	a4stg_frac_sng_nx,
	a1stg_expadd2,
	a1stg_expadd4_inv,
	a3stg_denorm,
	a3stg_denorm_inv,
	a4stg_denorm_inv,
	a3stg_exp,
	a4stg_round,
	a3stg_lead0,
	a4stg_rnd_frac_40,
	a4stg_rnd_frac_39,
	a4stg_rnd_frac_11,
	a4stg_rnd_frac_10,
	a4stg_frac_38_0_nx,
	a4stg_frac_9_0_nx,
	arst_l,
	grst_l,
	rclk,
	
	add_pipe_active,
	a1stg_denorm_sng_in1,
	a1stg_denorm_dbl_in1,
	a1stg_denorm_sng_in2,
	a1stg_denorm_dbl_in2,
	a1stg_norm_sng_in1,
	a1stg_norm_dbl_in1,
	a1stg_norm_sng_in2,
	a1stg_norm_dbl_in2,
	a1stg_step,
	a1stg_stepa,
	a1stg_sngop,
	a1stg_intlngop,
	a1stg_fsdtoix,
	a1stg_fstod,
	a1stg_fstoi,
	a1stg_fstox,
	a1stg_fdtoi,
	a1stg_fdtox,
	a1stg_faddsubs,
	a1stg_faddsubd,
	a1stg_fdtos,
	a2stg_faddsubop,
	a2stg_fsdtoix_fdtos,
	a2stg_fitos,
	a2stg_fitod,
	a2stg_fxtos,
	a2stg_fxtod,
	a3stg_faddsubop,
	a3stg_faddsubopa,
	a4stg_dblop,
	a6stg_fadd_in,
	add_id_out_in,
	add_fcc_out,
	a6stg_dbl_dst,
	a6stg_sng_dst,
	a6stg_long_dst,
	a6stg_int_dst,
	a6stg_fcmpop,
	a6stg_step,
	a3stg_sub_in,
	add_sign_out,
	add_cc_out,
	a4stg_in_of,
	add_exc_out,
	a2stg_frac1_in_frac1,
	a2stg_frac1_in_frac2,
	a1stg_2nan_in_inv,
	a1stg_faddsubop_inv,
	a2stg_frac1_in_qnan,
	a2stg_frac1_in_nv,
	a2stg_frac1_in_nv_dbl,
	a2stg_frac2_in_frac1,
	a2stg_frac2_in_qnan,
	a2stg_shr_cnt_in,
	a2stg_shr_cnt_5_inv_in,
	a2stg_shr_frac2_shr_int,
	a2stg_shr_frac2_shr_dbl,
	a2stg_shr_frac2_shr_sng,
	a2stg_shr_frac2_max,
	a2stg_sub_step,
	a2stg_fracadd_frac2_inv_in,
	a2stg_fracadd_frac2_inv_shr1_in,
	a2stg_fracadd_frac2,
	a2stg_fracadd_cin_in,
	a3stg_exp_7ff,
	a3stg_exp_ff,
	a3stg_exp_add,
	a2stg_expdec_neq_0,
	a3stg_exp10_0_eq0,
	a3stg_exp10_1_eq0,
	a3stg_fdtos_inv,
	a4stg_fixtos_fxtod_inv,
	a4stg_rnd_frac_add_inv,
	a4stg_shl_cnt_in,
	a4stg_rnd_sng,
	a4stg_rnd_dbl,
	add_frac_out_rndadd,
	add_frac_out_rnd_frac,
	add_frac_out_shl,
	a4stg_to_0,
	add_exp_out_expinc,
	add_exp_out_exp,
	add_exp_out_exp1,
	add_exp_out_expadd,
	a4stg_to_0_inv,
	se,
	si,
	so
);
parameter
		FADDS=	8'h41,
		FADDD=	8'h42,
		FSUBS=	8'h45,
		FSUBD=	8'h46,
		FCMPS=	8'h51,
		FCMPD=	8'h52,
		FCMPES=	8'h55,
		FCMPED=	8'h56,
		FSTOX=	8'h81,
		FDTOX=	8'h82,
		FSTOI=	8'hd1,
		FDTOI=	8'hd2,
		FSTOD=	8'hc9,
		FDTOS=	8'hc6,
		FXTOS=	8'h84,
		FXTOD=	8'h88,
		FITOS=	8'hc4,
		FITOD=	8'hc8;
input		inq_in1_51;		
input		inq_in1_54;		
input		inq_in1_63;		
input		inq_in1_50_0_neq_0;	
input		inq_in1_53_32_neq_0;	
input		inq_in1_exp_eq_0;	
input		inq_in1_exp_neq_ffs;	
input		inq_in2_51;		
input		inq_in2_54;		
input		inq_in2_63;		
input		inq_in2_50_0_neq_0;	
input		inq_in2_53_32_neq_0;	
input		inq_in2_exp_eq_0;	
input		inq_in2_exp_neq_ffs;	
input [7:0]	inq_op;			
input [1:0]	inq_rnd_mode;		
input [4:0]	inq_id;			
input [1:0]	inq_fcc;		
input		inq_add;		
input		add_dest_rdy;		
input		a1stg_in2_neq_in1_frac;	
input		a1stg_in2_gt_in1_frac;	
input		a1stg_in2_eq_in1_exp;	
input [11:0]	a1stg_expadd1;		
input [11:0]	a2stg_expadd;		
input		a2stg_frac2hi_neq_0;	
input		a2stg_frac2lo_neq_0;	
input [11:0]	a2stg_exp;		
input		a3stg_fsdtoix_nx;	
input		a3stg_fsdtoi_nx;	
input		a2stg_frac2_63;		
input [11:0]	a4stg_exp;		
input		add_of_out_cout;	
input		a4stg_frac_neq_0;	
input		a4stg_shl_data_neq_0;	
input		a4stg_frac_dbl_nx;	
input		a4stg_frac_sng_nx;	
input [5:0]	a1stg_expadd2;		
input [10:0]	a1stg_expadd4_inv;	
input		a3stg_denorm;		
input		a3stg_denorm_inv;	
input		a4stg_denorm_inv;	
input [10:0]	a3stg_exp;		
input		a4stg_round;		
input [5:0]	a3stg_lead0;		
input		a4stg_rnd_frac_40;	
input		a4stg_rnd_frac_39;	
input		a4stg_rnd_frac_11;	
input		a4stg_rnd_frac_10;	
input		a4stg_frac_38_0_nx;	
input		a4stg_frac_9_0_nx;	
input		arst_l;			
input		grst_l;			
input		rclk;		
output		add_pipe_active;        
output		a1stg_denorm_sng_in1;	
output		a1stg_denorm_dbl_in1;	
output		a1stg_denorm_sng_in2;	
output		a1stg_denorm_dbl_in2;	
output		a1stg_norm_sng_in1;	
output		a1stg_norm_dbl_in1;	
output		a1stg_norm_sng_in2;	
output		a1stg_norm_dbl_in2;	
output		a1stg_step;		
output		a1stg_stepa;		
output		a1stg_sngop;		
output		a1stg_intlngop;		
output		a1stg_fsdtoix;		
output		a1stg_fstod;		
output		a1stg_fstoi;		
output		a1stg_fstox;		
output		a1stg_fdtoi;		
output		a1stg_fdtox;		
output		a1stg_faddsubs;		
output		a1stg_faddsubd;		
output		a1stg_fdtos;		
output		a2stg_faddsubop;	
output		a2stg_fsdtoix_fdtos;	
output		a2stg_fitos;		
output		a2stg_fitod;		
output		a2stg_fxtos;		
output		a2stg_fxtod;		
output		a3stg_faddsubop;	
output [1:0]	a3stg_faddsubopa;	
output		a4stg_dblop;		
output		a6stg_fadd_in;		
output [9:0]	add_id_out_in;		
output [1:0]	add_fcc_out;		
output		a6stg_dbl_dst;		
output		a6stg_sng_dst;		
output		a6stg_long_dst;		
output		a6stg_int_dst;		
output		a6stg_fcmpop;		
output		a6stg_step;		
output		a3stg_sub_in;		
output		add_sign_out;		
output [1:0]	add_cc_out;		
output		a4stg_in_of;		
output [4:0]	add_exc_out;		
output		a2stg_frac1_in_frac1;	
output		a2stg_frac1_in_frac2;	
output		a1stg_2nan_in_inv;	
output		a1stg_faddsubop_inv;	
output		a2stg_frac1_in_qnan;	
output		a2stg_frac1_in_nv;	
output		a2stg_frac1_in_nv_dbl;	
output		a2stg_frac2_in_frac1;	
output		a2stg_frac2_in_qnan;	
output [5:0]	a2stg_shr_cnt_in;	
output    a2stg_shr_cnt_5_inv_in; 
output		a2stg_shr_frac2_shr_int; 
output		a2stg_shr_frac2_shr_dbl; 
output		a2stg_shr_frac2_shr_sng; 
output		a2stg_shr_frac2_max;	
output		a2stg_sub_step;		
output		a2stg_fracadd_frac2_inv_in; 
output		a2stg_fracadd_frac2_inv_shr1_in; 
output		a2stg_fracadd_frac2;	
output		a2stg_fracadd_cin_in;	
output		a3stg_exp_7ff;		
output		a3stg_exp_ff;		
output		a3stg_exp_add;		
output		a2stg_expdec_neq_0;	
output		a3stg_exp10_0_eq0;	
output		a3stg_exp10_1_eq0;	
output		a3stg_fdtos_inv;	
output		a4stg_fixtos_fxtod_inv;	
output		a4stg_rnd_frac_add_inv; 
output [9:0]	a4stg_shl_cnt_in;	
output		a4stg_rnd_sng;		
output		a4stg_rnd_dbl;		
output		add_frac_out_rndadd;	
output		add_frac_out_rnd_frac;	
output		add_frac_out_shl;	
output		a4stg_to_0;		
output		add_exp_out_expinc;	
output		add_exp_out_exp;	
output		add_exp_out_exp1;	
output		add_exp_out_expadd;	
output		a4stg_to_0_inv;		
input		se;			
input		si;			
output		so;			
wire		reset;
wire		a1stg_in1_51;
wire		a1stg_in1_54;
wire		a1stg_in1_63;
wire		a1stg_in1_50_0_neq_0;
wire		a1stg_in1_53_32_neq_0;
wire		a1stg_in1_exp_eq_0;
wire		a1stg_in1_exp_neq_ffs;
wire		a1stg_in2_51;
wire		a1stg_in2_54;
wire		a1stg_in2_63;
wire		a1stg_in2_50_0_neq_0;
wire		a1stg_in2_53_32_neq_0;
wire		a1stg_in2_exp_eq_0;
wire		a1stg_in2_exp_neq_ffs;
wire		a1stg_denorm_sng_in1;
wire		a1stg_denorm_dbl_in1;
wire		a1stg_denorm_sng_in2;
wire		a1stg_denorm_dbl_in2;
wire		a1stg_norm_sng_in1;
wire		a1stg_norm_dbl_in1;
wire		a1stg_norm_sng_in2;
wire		a1stg_norm_dbl_in2;
wire		a1stg_snan_sng_in1;
wire		a1stg_snan_dbl_in1;
wire		a1stg_snan_sng_in2;
wire		a1stg_snan_dbl_in2;
wire		a1stg_qnan_sng_in1;
wire		a1stg_qnan_dbl_in1;
wire		a1stg_qnan_sng_in2;
wire		a1stg_qnan_dbl_in2;
wire		a1stg_snan_in1;
wire		a1stg_snan_in2;
wire		a1stg_qnan_in1;
wire		a1stg_qnan_in2;
wire		a1stg_nan_sng_in1;
wire		a1stg_nan_dbl_in1;
wire		a1stg_nan_sng_in2;
wire		a1stg_nan_dbl_in2;
wire		a1stg_nan_in1;
wire		a1stg_nan_in2;
wire		a1stg_nan_in;
wire		a1stg_2nan_in;
wire		a1stg_inf_sng_in1;
wire		a1stg_inf_dbl_in1;
wire		a1stg_inf_sng_in2;
wire		a1stg_inf_dbl_in2;
wire		a1stg_inf_in1;
wire		a1stg_inf_in2;
wire		a1stg_2inf_in;
wire		a1stg_infnan_sng_in1;
wire		a1stg_infnan_dbl_in1;
wire		a1stg_infnan_sng_in2;
wire		a1stg_infnan_dbl_in2;
wire		a1stg_infnan_in1;
wire		a1stg_infnan_in2;
wire		a1stg_infnan_in;
wire		a1stg_2zero_in;
wire		a1stg_step;
wire		a1stg_stepa;
wire [7:0]	a1stg_op_in;
wire [7:0]	a1stg_op;
wire		a1stg_sngop;
wire [3:0]	a1stg_sngopa;
wire		a1stg_dblop;
wire [3:0]	a1stg_dblopa;
wire [1:0]	a1stg_rnd_mode;
wire [4:0]	a1stg_id;
wire [1:0]	a1stg_fcc;
wire		a1stg_fadd;
wire		a1stg_dbl_dst;
wire		a1stg_sng_dst;
wire		a1stg_long_dst;
wire		a1stg_int_dst;
wire		a1stg_intlngop;
wire		a1stg_faddsubop;
wire		a1stg_fsubop;
wire		a1stg_fsdtox;
wire		a1stg_fcmpesd;
wire		a1stg_fcmpsd;
wire		a1stg_faddsub_dtosop;
wire		a1stg_fdtoix;
wire		a1stg_fstoix;
wire		a1stg_fsdtoix;
wire		a1stg_fixtosd;
wire		a1stg_fstod;
wire		a1stg_fstoi;
wire		a1stg_fstox;
wire		a1stg_fdtoi;
wire		a1stg_fdtox;
wire		a1stg_fsdtoix_fdtos;
wire		a1stg_fitos;
wire		a1stg_fitod;
wire		a1stg_fxtos;
wire		a1stg_fcmpop;
wire		a1stg_f4cycop;
wire		a1stg_fixtos_fxtod;
wire		a1stg_faddsubs_fdtos;
wire		a1stg_faddsubs;
wire		a1stg_faddsubd;
wire		a1stg_fdtos;
wire		a1stg_fistod;
wire		a1stg_fixtos;
wire		a1stg_fxtod;
wire            a1stg_opdec_36;
wire [34:28]	a1stg_opdec;
wire [3:0]      a1stg_opdec_24_21;
wire [8:0]      a1stg_opdec_19_11;
wire [9:0]      a1stg_opdec_9_0;
wire		fixtosd_hold;
wire [30:0]	a2stg_opdec_in;
wire            a2stg_opdec_36;
wire [34:28]	a2stg_opdec;
wire [3:0]      a2stg_opdec_24_21;
wire [8:0]      a2stg_opdec_19_11;
wire [9:0]      a2stg_opdec_9_0;
wire [1:0]	a2stg_rnd_mode;
wire [4:0]	a2stg_id;
wire [1:0]	a2stg_fcc;
wire		a2stg_fadd;
wire		a2stg_long_dst;
wire		a2stg_faddsubop;
wire		a2stg_fsubop;
wire		a2stg_faddsub_dtosop;
wire		a2stg_fdtoix;
wire		a2stg_fstoix;
wire		a2stg_fsdtoix;
wire		a2stg_fstod;
wire		a2stg_fstoi;
wire		a2stg_fstox;
wire		a2stg_fdtoi;
wire		a2stg_fdtox;
wire		a2stg_fsdtoix_fdtos;
wire		a2stg_fitos;
wire		a2stg_fitod;
wire		a2stg_fxtos;
wire		a2stg_fcmpop;
wire		a2stg_fixtos_fxtod;
wire		a2stg_fdtos;
wire		a2stg_fxtod;
wire            a3stg_opdec_36;
wire [34:29]	a3stg_opdec;
wire            a3stg_opdec_24;
wire            a3stg_opdec_21;
wire [9:0]      a3stg_opdec_9_0;
wire [1:0]	a3stg_rnd_mode;
wire [4:0]	a3stg_id;
wire [1:0]	a3stg_fcc;
wire		a3stg_fadd;
wire		a3stg_int_dst;
wire		a3stg_faddsubop;
wire [1:0]	a3stg_faddsubopa;
wire		a3stg_fsdtoix;
wire		a3stg_f4cycop;
wire		a3stg_fixtos_fxtod;
wire		a3stg_fdtos;
wire            a4stg_opdec_36;
wire [34:29]	a4stg_opdec;
wire            a4stg_opdec_24;
wire            a4stg_opdec_21;
wire            a4stg_opdec_9;
wire [7:0]      a4stg_opdec_7_0;
wire [1:0]	a4stg_rnd_mode_in;
wire [1:0]	a4stg_rnd_mode;
wire [1:0]	a4stg_rnd_mode2;
wire [9:0]	a4stg_id_in;
wire [9:0]	a4stg_id;
wire [1:0]	a4stg_fcc;
wire		a4stg_dblop;
wire		a4stg_fadd;
wire		a4stg_faddsubop;
wire		a4stg_faddsub_dtosop;
wire		a4stg_fsdtoix;
wire		a4stg_fcmpop;
wire		a4stg_fixtos_fxtod;
wire		a4stg_faddsubs_fdtos;
wire		a4stg_faddsubs;
wire		a4stg_faddsubd;
wire		a4stg_fdtos;
wire		a4stg_fistod;
wire [34:30]	a5stg_opdec;
wire            a5stg_opdec_9;
wire            a5stg_opdec_7;
wire            a5stg_opdec_1;
wire            a5stg_opdec_0;
wire [9:0]	a5stg_id;
wire		a5stg_fadd;
wire		a5stg_fixtos_fxtod;
wire		a5stg_fixtos;
wire		a5stg_fxtod;
wire [34:30]	a6stg_opdec_in;
wire            a6stg_opdec_in_9;
wire		a6stg_fadd_in;
wire [34:30]	a6stg_opdec;
wire            a6stg_opdec_9;
wire [9:0]	add_id_out_in;
wire [9:0]	add_id_out;
wire [1:0]	add_fcc_out_in;
wire [1:0]	add_fcc_out;
wire		a6stg_fadd;
wire		a6stg_dbl_dst;
wire		a6stg_sng_dst;
wire		a6stg_long_dst;
wire		a6stg_int_dst;
wire		a6stg_fcmpop;
wire		a6stg_hold;
wire		a6stg_step;
wire		a1stg_sub;
wire		a2stg_sign1;
wire		a2stg_sign2;
wire		a2stg_sub;
wire		a2stg_in2_neq_in1_frac;
wire		a2stg_in2_gt_in1_frac;
wire		a2stg_in2_eq_in1_exp;
wire		a2stg_in2_gt_in1_exp;
wire		a2stg_nan_in;
wire		a2stg_nan_in2;
wire		a2stg_snan_in2;
wire		a2stg_qnan_in2;
wire		a2stg_snan_in1;
wire		a2stg_qnan_in1;
wire		a2stg_2zero_in;
wire		a2stg_2inf_in;
wire		a2stg_in2_eq_in1;
wire		a2stg_in2_gt_in1;
wire		a3stg_sub_in;
wire		a2stg_faddsub_sign;
wire		a3stg_sign_in;
wire		a3stg_sign;
wire		a2stg_cc_1;
wire		a2stg_cc_0;
wire [1:0]	a2stg_cc;
wire [1:0]	a3stg_cc;
wire		a4stg_sign_in;
wire		a4stg_sign;
wire		a4stg_sign2;
wire [1:0]	a4stg_cc;
wire		add_sign_out;
wire [1:0]	add_cc_out_in;
wire [1:0]	add_cc_out;
wire		a1stg_nv;
wire		a2stg_nv;
wire		a1stg_of_mask;
wire		a2stg_of_mask;
wire		a3stg_nv_in;
wire		a3stg_nv;
wire		a3stg_of_mask;
wire		a2stg_nx_tmp1;
wire		a2stg_nx_tmp2;
wire		a2stg_nx_tmp3;
wire		a3stg_a2_expadd_11;
wire		a3stg_nx_tmp1;
wire		a3stg_nx_tmp2;
wire		a3stg_nx_tmp3;
wire		a3stg_nx;
wire		a4stg_nv_in;
wire		a4stg_nv;
wire		a4stg_nv2;
wire		a4stg_of_mask_in;
wire		a4stg_of_mask;
wire		a4stg_of_mask2;
wire		a4stg_nx_in;
wire		a4stg_nx;
wire		a4stg_nx2;
wire		add_nv_out;
wire		a4stg_in_of;
wire		add_of_out_tmp1_in;
wire		add_of_out_tmp1;
wire		add_of_out_tmp2;
wire		add_of_out;
wire		a4stg_uf;
wire		add_uf_out;
wire		add_nx_out_in;
wire		add_nx_out;
wire [4:0]	add_exc_out;
wire		a2stg_frac1_in_frac1;
wire		a2stg_frac1_in_frac2;
wire		a1stg_2nan_in_inv;
wire		a1stg_faddsubop_inv;
wire		a2stg_frac1_in_qnan;
wire		a2stg_frac1_in_nv;
wire		a2stg_frac1_in_nv_dbl;
wire		a2stg_frac2_in_frac1;
wire		a2stg_frac2_in_qnan;
wire		a1stg_exp_diff_add1;
wire		a1stg_exp_diff_add2;
wire		a1stg_exp_diff_5;
wire [10:0]	a1stg_exp_diff;
wire [5:0]	a1stg_clamp63;
wire [5:0]	a2stg_shr_cnt_in;
wire    a2stg_shr_cnt_5_inv_in;
wire		a2stg_shr_frac2_shr_int;
wire		a2stg_shr_frac2_shr_dbl;
wire		a2stg_shr_frac2_shr_sng;
wire		a2stg_shr_frac2_max;
wire		a2stg_sub_step;
wire		a1stg_faddsub_clamp63_0;
wire		a2stg_fracadd_frac2_inv_in;
wire		a2stg_fracadd_frac2_inv_shr1_in;
wire		a2stg_fracadd_frac2_in;
wire		a2stg_fracadd_frac2;
wire		a2stg_fracadd_cin_in;
wire		a3stg_exp_7ff;
wire		a3stg_exp_ff;
wire		a3stg_exp_add;
wire		a2stg_expdec_neq_0;
wire		a3stg_exp10_0_eq0;
wire		a3stg_exp10_1_eq0;
wire		a3stg_fdtos_inv;
wire		a4stg_fixtos_fxtod_inv;
wire		a4stg_rnd_frac_add_inv;
wire [9:0]	a4stg_shl_cnt_in;
wire		a4stg_rnd_sng;
wire		a4stg_rnd_dbl;
wire		a4stg_rndup_sng;
wire		a4stg_rndup_dbl;
wire		a4stg_rndup;
wire		a5stg_rndup;
wire		add_frac_out_rndadd;
wire		add_frac_out_rnd_frac;
wire		add_frac_out_shl;
wire		a4stg_to_0;
wire		add_exp_out_expinc;
wire		add_exp_out_exp;
wire		add_exp_out_exp1;
wire		add_exp_out_expadd;
wire		a4stg_to_0_inv;
wire		add_pipe_active_in;
wire		add_pipe_active;
wire        add_ctl_rst_l;
dffrl_async #(1)  dffrl_add_ctl (
  .din  (grst_l),
  .clk  (rclk),
  .rst_l(arst_l),
  .q    (add_ctl_rst_l),
	.se (se),
	.si (),
	.so ()
  );
assign reset= (!add_ctl_rst_l);
dffe_s #(1) i_a1stg_in1_51 (
	.din	(inq_in1_51),
	.en     (a1stg_step),
        .clk    (rclk),
 
        .q      (a1stg_in1_51),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a1stg_in1_54 (
	.din	(inq_in1_54),
	.en     (a1stg_step),
        .clk    (rclk),
 
        .q      (a1stg_in1_54),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a1stg_in1_63 (
        .din	(inq_in1_63),
        .en	(a1stg_step),
        .clk	(rclk),
 
        .q	(a1stg_in1_63),
 
        .se	(se),
        .si	(),
        .so	()
);
dffe_s #(1) i_a1stg_in1_50_0_neq_0 (
	.din	(inq_in1_50_0_neq_0),
	.en	(a1stg_step),
	.clk	(rclk),
	.q	(a1stg_in1_50_0_neq_0),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_a1stg_in1_53_32_neq_0 (
	.din	(inq_in1_53_32_neq_0),
	.en	(a1stg_step),
	.clk	(rclk),
	.q	(a1stg_in1_53_32_neq_0),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_a1stg_in1_exp_eq_0 (
        .din	(inq_in1_exp_eq_0),
        .en	(a1stg_step),
        .clk	(rclk),
 
        .q	(a1stg_in1_exp_eq_0),
 
        .se	(se),
        .si	(),
        .so	()
);
dffe_s #(1) i_a1stg_in1_exp_neq_ffs (
	.din	(inq_in1_exp_neq_ffs),
	.en	(a1stg_step),
	.clk	(rclk),
	.q	(a1stg_in1_exp_neq_ffs),
   	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_a1stg_in2_51 (
	.din	(inq_in2_51),
	.en	(a1stg_step),
	.clk	(rclk),
	.q	(a1stg_in2_51),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_a1stg_in2_54 (
	.din	(inq_in2_54),
	.en	(a1stg_step),
	.clk	(rclk),
	.q	(a1stg_in2_54),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_a1stg_in2_63 (
        .din	(inq_in2_63),
        .en	(a1stg_step),
        .clk	(rclk),
 
        .q	(a1stg_in2_63),
 
        .se	(se),
        .si	(),
        .so	()
);
dffe_s #(1) i_a1stg_in2_50_0_neq_0 (
	.din	(inq_in2_50_0_neq_0),
	.en	(a1stg_step),
	.clk	(rclk),
	.q	(a1stg_in2_50_0_neq_0),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_a1stg_in2_53_32_neq_0 (
	.din	(inq_in2_53_32_neq_0),
	.en	(a1stg_step),
	.clk	(rclk),
	.q	(a1stg_in2_53_32_neq_0),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_a1stg_in2_exp_eq_0 (
	.din	(inq_in2_exp_eq_0),
	 .en	(a1stg_step),
	.clk	(rclk),
	.q	(a1stg_in2_exp_eq_0),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_a1stg_in2_exp_neq_ffs (
        .din	(inq_in2_exp_neq_ffs),
        .en	(a1stg_step),
        .clk	(rclk),
 
        .q	(a1stg_in2_exp_neq_ffs),
 
        .se	(se),
        .si	(),
        .so	()
);
assign a1stg_denorm_sng_in1= a1stg_in1_exp_eq_0 && a1stg_sngopa[0];
assign a1stg_denorm_dbl_in1= a1stg_in1_exp_eq_0 && a1stg_dblopa[0];
assign a1stg_denorm_sng_in2= a1stg_in2_exp_eq_0 && a1stg_sngopa[0];
assign a1stg_denorm_dbl_in2= a1stg_in2_exp_eq_0 && a1stg_dblopa[0];
assign a1stg_norm_sng_in1= (!a1stg_in1_exp_eq_0) && a1stg_sngopa[0];
assign a1stg_norm_dbl_in1= (!a1stg_in1_exp_eq_0) && a1stg_dblopa[0];
assign a1stg_norm_sng_in2= (!a1stg_in2_exp_eq_0) && a1stg_sngopa[0];
assign a1stg_norm_dbl_in2= (!a1stg_in2_exp_eq_0) && a1stg_dblopa[0];
assign a1stg_snan_sng_in1= (!a1stg_in1_exp_neq_ffs) && (!a1stg_in1_54)
		&& a1stg_in1_53_32_neq_0 && a1stg_sngopa[1];
assign a1stg_snan_dbl_in1= (!a1stg_in1_exp_neq_ffs) && (!a1stg_in1_51)
		&& a1stg_in1_50_0_neq_0 && a1stg_dblopa[1];
assign a1stg_snan_sng_in2= (!a1stg_in2_exp_neq_ffs) && (!a1stg_in2_54)
                && a1stg_in2_53_32_neq_0 && a1stg_sngopa[1];
assign a1stg_snan_dbl_in2= (!a1stg_in2_exp_neq_ffs) && (!a1stg_in2_51)
                && a1stg_in2_50_0_neq_0 && a1stg_dblopa[1];
assign a1stg_qnan_sng_in1= (!a1stg_in1_exp_neq_ffs) && a1stg_in1_54
		&& a1stg_sngopa[1];
assign a1stg_qnan_dbl_in1= (!a1stg_in1_exp_neq_ffs) && a1stg_in1_51
		&& a1stg_dblopa[1];
assign a1stg_qnan_sng_in2= (!a1stg_in2_exp_neq_ffs) && a1stg_in2_54
                && a1stg_sngopa[1];
assign a1stg_qnan_dbl_in2= (!a1stg_in2_exp_neq_ffs) && a1stg_in2_51
                && a1stg_dblopa[1];
assign a1stg_snan_in1= a1stg_snan_sng_in1 || a1stg_snan_dbl_in1;
assign a1stg_snan_in2= a1stg_snan_sng_in2 || a1stg_snan_dbl_in2;
assign a1stg_qnan_in1= a1stg_qnan_sng_in1 || a1stg_qnan_dbl_in1;
 
assign a1stg_qnan_in2= a1stg_qnan_sng_in2 || a1stg_qnan_dbl_in2;
assign a1stg_nan_sng_in1= (!a1stg_in1_exp_neq_ffs)
		&& (a1stg_in1_54 || a1stg_in1_53_32_neq_0)
		&& a1stg_sngopa[2];
assign a1stg_nan_dbl_in1= (!a1stg_in1_exp_neq_ffs)
		&& (a1stg_in1_51 || a1stg_in1_50_0_neq_0)
		&& a1stg_dblopa[2];
assign a1stg_nan_sng_in2= (!a1stg_in2_exp_neq_ffs)
		&& (a1stg_in2_54 || a1stg_in2_53_32_neq_0)
		&& a1stg_sngopa[2];
assign a1stg_nan_dbl_in2= (!a1stg_in2_exp_neq_ffs)
		&& (a1stg_in2_51 || a1stg_in2_50_0_neq_0)
		&& a1stg_dblopa[2];
assign a1stg_nan_in1= a1stg_nan_sng_in1 || a1stg_nan_dbl_in1;
assign a1stg_nan_in2= a1stg_nan_sng_in2 || a1stg_nan_dbl_in2;
assign a1stg_nan_in= a1stg_nan_in1 || a1stg_nan_in2;
assign a1stg_2nan_in= a1stg_nan_in1 && a1stg_nan_in2;
assign a1stg_inf_sng_in1= (!a1stg_in1_exp_neq_ffs)
		&& (!a1stg_in1_54) && (!a1stg_in1_53_32_neq_0)
		&& a1stg_sngopa[2];
assign a1stg_inf_dbl_in1= (!a1stg_in1_exp_neq_ffs)
		&& (!a1stg_in1_51) && (!a1stg_in1_50_0_neq_0)
		&& a1stg_dblopa[2];
assign a1stg_inf_sng_in2= (!a1stg_in2_exp_neq_ffs)
		&& (!a1stg_in2_54) && (!a1stg_in2_53_32_neq_0)
		&& a1stg_sngopa[2];
assign a1stg_inf_dbl_in2= (!a1stg_in2_exp_neq_ffs)
		&& (!a1stg_in2_51) && (!a1stg_in2_50_0_neq_0)
		&& a1stg_dblopa[2];
assign a1stg_inf_in1= a1stg_inf_sng_in1 || a1stg_inf_dbl_in1;
assign a1stg_inf_in2= a1stg_inf_sng_in2 || a1stg_inf_dbl_in2;
assign a1stg_2inf_in= a1stg_inf_in1 && a1stg_inf_in2;
assign a1stg_infnan_sng_in1= (!a1stg_in1_exp_neq_ffs) && a1stg_sngopa[3];
assign a1stg_infnan_dbl_in1= (!a1stg_in1_exp_neq_ffs) && a1stg_dblopa[3];
assign a1stg_infnan_sng_in2= (!a1stg_in2_exp_neq_ffs) && a1stg_sngopa[3];
assign a1stg_infnan_dbl_in2= (!a1stg_in2_exp_neq_ffs) && a1stg_dblopa[3];
assign a1stg_infnan_in1= a1stg_infnan_sng_in1 || a1stg_infnan_dbl_in1;
assign a1stg_infnan_in2= a1stg_infnan_sng_in2 || a1stg_infnan_dbl_in2;
assign a1stg_infnan_in= a1stg_infnan_in1 || a1stg_infnan_in2;
assign a1stg_2zero_in =
		a1stg_in1_exp_eq_0                          &&
                (!a1stg_in1_54          || a1stg_dblopa[3]) &&  
                (!a1stg_in1_53_32_neq_0 || a1stg_dblopa[3]) &&  
                (!a1stg_in1_51)                             &&
                (!a1stg_in1_50_0_neq_0)                     &&
                a1stg_in2_exp_eq_0                          &&
                (!a1stg_in2_54          || a1stg_dblopa[3]) &&  
                (!a1stg_in2_53_32_neq_0 || a1stg_dblopa[3]) &&  
                (!a1stg_in2_51)                             &&
                (!a1stg_in2_50_0_neq_0);
assign a1stg_step= (!fixtosd_hold) && (!a6stg_hold);
assign a1stg_stepa= a1stg_step;
assign a1stg_op_in[7:0]= ({8{inq_add}}
			    & inq_op[7:0]);
dffre_s #(8) i_a1stg_op (
        .din    (a1stg_op_in[7:0]),
        .en     (a1stg_step),
        .rst    (reset),
        .clk    (rclk),
        .q      (a1stg_op[7:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a1stg_sngop (
	.din	(inq_op[0]),
        .en     (a1stg_step),
        .clk    (rclk),
        .q      (a1stg_sngop),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(4) i_a1stg_sngopa (
        .din	({4{inq_op[0]}}),
        .en	(a1stg_step),
        .clk	(rclk),
 
        .q	(a1stg_sngopa[3:0]),
 
        .se	(se),
        .si	(),
        .so	()
);
dffe_s #(1) i_a1stg_dblop (
	.din	(inq_op[1]),
        .en     (a1stg_step),
        .clk    (rclk),
 
        .q      (a1stg_dblop),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(4) i_a1stg_dblopa (
 	.din	({4{inq_op[1]}}),
	.en	(a1stg_step),
	.clk	(rclk),
	.q	(a1stg_dblopa[3:0]),
 
        .se	(se),
        .si	(),
        .so	()
);
dffe_s #(2) i_a1stg_rnd_mode (
        .din    (inq_rnd_mode[1:0]),
        .en     (a1stg_step),
        .clk    (rclk),
        .q      (a1stg_rnd_mode[1:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(5) i_a1stg_id (
        .din    (inq_id[4:0]),
        .en     (a1stg_step),
        .clk    (rclk),
 
        .q      (a1stg_id[4:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(2) i_a1stg_fcc (
        .din    (inq_fcc[1:0]),
        .en     (a1stg_step),
        .clk    (rclk),
        .q      (a1stg_fcc[1:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign a1stg_fadd= (a1stg_op[7:0]==FADDS) || (a1stg_op[7:0]==FADDD)
		|| (a1stg_op[7:0]==FSUBS) || (a1stg_op[7:0]==FSUBD)
		|| (a1stg_op[7:0]==FCMPES) || (a1stg_op[7:0]==FCMPED)
		|| (a1stg_op[7:0]==FCMPS) || (a1stg_op[7:0]==FCMPD)
		|| (a1stg_op[7:0]==FITOS) || (a1stg_op[7:0]==FITOD)
		|| (a1stg_op[7:0]==FXTOS) || (a1stg_op[7:0]==FXTOD)
		|| (a1stg_op[7:0]==FSTOI) || (a1stg_op[7:0]==FSTOX)
		|| (a1stg_op[7:0]==FDTOI) || (a1stg_op[7:0]==FDTOX)
		|| (a1stg_op[7:0]==FSTOD) || (a1stg_op[7:0]==FDTOS);
assign a1stg_dbl_dst= (a1stg_op[7:0]==FADDD) || (a1stg_op[7:0]==FSUBD)
		|| (a1stg_op[7:0]==FITOD) || (a1stg_op[7:0]==FXTOD)
		|| (a1stg_op[7:0]==FSTOD);
assign a1stg_sng_dst= (a1stg_op[7:0]==FADDS) || (a1stg_op[7:0]==FSUBS)
		|| (a1stg_op[7:0]==FITOS) || (a1stg_op[7:0]==FXTOS)
		|| (a1stg_op[7:0]==FDTOS);
assign a1stg_long_dst= (a1stg_op[7:0]==FSTOX) || (a1stg_op[7:0]==FDTOX);
assign a1stg_int_dst= (a1stg_op[7:0]==FSTOI) || (a1stg_op[7:0]==FDTOI);
assign a1stg_intlngop= (!(a1stg_sngopa[3] || a1stg_dblop));
assign a1stg_faddsubop= (a1stg_op[7:0]==FADDS) || (a1stg_op[7:0]==FADDD)
		|| (a1stg_op[7:0]==FSUBS) || (a1stg_op[7:0]==FSUBD);
assign a1stg_fsubop= (a1stg_op[7:0]==FSUBS) || (a1stg_op[7:0]==FSUBD);
assign a1stg_fsdtox= (a1stg_op[7:0]==FSTOX) || (a1stg_op[7:0]==FDTOX);
assign a1stg_fcmpesd= (a1stg_op[7:0]==FCMPES) || (a1stg_op[7:0]==FCMPED);
assign a1stg_fcmpsd= (a1stg_op[7:0]==FCMPS) || (a1stg_op[7:0]==FCMPD);
assign a1stg_faddsub_dtosop= (a1stg_op[7:0]==FADDS) || (a1stg_op[7:0]==FADDD)
                || (a1stg_op[7:0]==FSUBS) || (a1stg_op[7:0]==FSUBD)
		|| (a1stg_op[7:0]==FDTOS);
assign a1stg_fdtoix= (a1stg_op[7:0]==FDTOI) || (a1stg_op[7:0]==FDTOX);
assign a1stg_fstoix= (a1stg_op[7:0]==FSTOI) || (a1stg_op[7:0]==FSTOX);
assign a1stg_fsdtoix= (a1stg_op[7:0]==FSTOI) || (a1stg_op[7:0]==FSTOX)
		|| (a1stg_op[7:0]==FDTOI) || (a1stg_op[7:0]==FDTOX);
assign a1stg_fixtosd= (a1stg_op[7:0]==FITOS) || (a1stg_op[7:0]==FITOD)
		|| (a1stg_op[7:0]==FXTOS) || (a1stg_op[7:0]==FXTOD);
assign a1stg_fstod= (a1stg_op[7:0]==FSTOD);
assign a1stg_fstoi= (a1stg_op[7:0]==FSTOI);
assign a1stg_fstox= (a1stg_op[7:0]==FSTOX);
assign a1stg_fdtoi= (a1stg_op[7:0]==FDTOI);
assign a1stg_fdtox= (a1stg_op[7:0]==FDTOX);
assign a1stg_fsdtoix_fdtos= (a1stg_op[7:0]==FSTOI) || (a1stg_op[7:0]==FSTOX)
                || (a1stg_op[7:0]==FDTOI) || (a1stg_op[7:0]==FDTOX)
		|| (a1stg_op[7:0]==FDTOS);
assign a1stg_fitos= (a1stg_op[7:0]==FITOS);
assign a1stg_fitod= (a1stg_op[7:0]==FITOD);
assign a1stg_fxtos= (a1stg_op[7:0]==FXTOS);
assign a1stg_fcmpop= (a1stg_op[7:0]==FCMPS) || (a1stg_op[7:0]==FCMPD)
		|| (a1stg_op[7:0]==FCMPES) || (a1stg_op[7:0]==FCMPED);
assign a1stg_f4cycop= (a1stg_op[7:0]==FADDS) || (a1stg_op[7:0]==FADDD)
                || (a1stg_op[7:0]==FSUBS) || (a1stg_op[7:0]==FSUBD)
                || (a1stg_op[7:0]==FDTOS) || (a1stg_op[7:0]==FSTOD)
		|| (a1stg_op[7:0]==FITOD);
assign a1stg_fixtos_fxtod= (a1stg_op[7:0]==FITOS) || (a1stg_op[7:0]==FXTOS)
		|| (a1stg_op[7:0]==FXTOD);
assign a1stg_faddsubs_fdtos= (a1stg_op[7:0]==FADDS) || (a1stg_op[7:0]==FSUBS)
		|| (a1stg_op[7:0]==FDTOS);
assign a1stg_faddsubs= (a1stg_op[7:0]==FADDS) || (a1stg_op[7:0]==FSUBS);
assign a1stg_faddsubd= (a1stg_op[7:0]==FADDD) || (a1stg_op[7:0]==FSUBD);
assign a1stg_fdtos= (a1stg_op[7:0]==FDTOS);
assign a1stg_fistod= (a1stg_op[7:0]==FITOD) || (a1stg_op[7:0]==FSTOD);
assign a1stg_fixtos= (a1stg_op[7:0]==FITOS) || (a1stg_op[7:0]==FXTOS);
assign a1stg_fxtod= (a1stg_op[7:0]==FXTOD);
assign a1stg_opdec_36 = a1stg_dblop;
assign a1stg_opdec[34:28] =
			 {a1stg_fadd,
			  a1stg_dbl_dst,
			  a1stg_sng_dst,
			  a1stg_long_dst,
			  a1stg_int_dst,
			  a1stg_faddsubop,
			  a1stg_fsubop};
assign a1stg_opdec_24_21[3:0] =
			 {a1stg_faddsub_dtosop,
			  a1stg_fdtoix,
			  a1stg_fstoix,
			  a1stg_fsdtoix};
assign a1stg_opdec_19_11[8:0] =
			 {a1stg_fstod,
			  a1stg_fstoi,
			  a1stg_fstox,
			  a1stg_fdtoi,
			  a1stg_fdtox,
			  a1stg_fsdtoix_fdtos,
			  a1stg_fitos,
			  a1stg_fitod,
			  a1stg_fxtos};
 
assign a1stg_opdec_9_0[9:0] = 
			 {a1stg_fcmpop,
			  a1stg_f4cycop,
			  a1stg_fixtos_fxtod,
			  a1stg_faddsubs_fdtos,
			  a1stg_faddsubs,
			  a1stg_faddsubd,
			  a1stg_fdtos,
			  a1stg_fistod,
			  a1stg_fixtos,
			  a1stg_fxtod};
assign fixtosd_hold= a2stg_fixtos_fxtod
		&& (!(a1stg_op[7] && (!a1stg_op[1]) && (!a1stg_op[0])
			&& (a1stg_op[2] || (!a1stg_op[6]))));
assign a2stg_opdec_in[30:0]= {31{(!fixtosd_hold)}}
			    & {a1stg_opdec_36, a1stg_opdec[34:28],
                               a1stg_opdec_24_21[3:0], a1stg_opdec_19_11[8:0],
                               a1stg_opdec_9_0[9:0]};
dffre_s #(31) i_a2stg_opdec (
	.din	(a2stg_opdec_in[30:0]),
	.en	(a6stg_step),
	.rst    (reset),
        .clk    (rclk),
        .q      ({a2stg_opdec_36, a2stg_opdec[34:28], a2stg_opdec_24_21[3:0],
                  a2stg_opdec_19_11[8:0], a2stg_opdec_9_0[9:0]}),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(2) i_a2stg_rnd_mode (
        .din    (a1stg_rnd_mode[1:0]),
        .en     (a6stg_step),
        .clk    (rclk),
        .q      (a2stg_rnd_mode[1:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(5) i_a2stg_id (
        .din    (a1stg_id[4:0]),
        .en     (a6stg_step),
        .clk    (rclk),
 
        .q      (a2stg_id[4:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(2) i_a2stg_fcc (
        .din    (a1stg_fcc[1:0]),
        .en     (a6stg_step),
        .clk    (rclk),
        .q      (a2stg_fcc[1:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign a2stg_fadd= a2stg_opdec[34];
assign a2stg_long_dst= a2stg_opdec[31];
assign a2stg_faddsubop= a2stg_opdec[29];
assign a2stg_fsubop= a2stg_opdec[28];
assign a2stg_faddsub_dtosop= a2stg_opdec_24_21[3];
assign a2stg_fdtoix= a2stg_opdec_24_21[2];
assign a2stg_fstoix= a2stg_opdec_24_21[1];
assign a2stg_fsdtoix= a2stg_opdec_24_21[0];
assign a2stg_fstod= a2stg_opdec_19_11[8];
assign a2stg_fstoi= a2stg_opdec_19_11[7];
assign a2stg_fstox= a2stg_opdec_19_11[6];
assign a2stg_fdtoi= a2stg_opdec_19_11[5];
assign a2stg_fdtox= a2stg_opdec_19_11[4];
assign a2stg_fsdtoix_fdtos= a2stg_opdec_19_11[3];
assign a2stg_fitos= a2stg_opdec_19_11[2];
assign a2stg_fitod= a2stg_opdec_19_11[1];
assign a2stg_fxtos= a2stg_opdec_19_11[0];
assign a2stg_fcmpop= a2stg_opdec_9_0[9];
assign a2stg_fixtos_fxtod= a2stg_opdec_9_0[7];
assign a2stg_fdtos= a2stg_opdec_9_0[3];
assign a2stg_fxtod= a2stg_opdec_9_0[0];
dffre_s #(19) i_a3stg_opdec (
        .din    ({a2stg_opdec_36, a2stg_opdec[34:29], a2stg_opdec_24_21[3],
                  a2stg_opdec_24_21[0], a2stg_opdec_9_0[9:0]}),
        .en     (a6stg_step),
        .rst    (reset),
        .clk    (rclk),
        .q      ({a3stg_opdec_36, a3stg_opdec[34:29], a3stg_opdec_24,
                  a3stg_opdec_21, a3stg_opdec_9_0[9:0]}),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(2) i_a3stg_faddsubopa (
	.din	({2{a2stg_faddsubop}}),
	.en	(a6stg_step),
	.rst	(reset),
	.clk	(rclk),
	.q	(a3stg_faddsubopa[1:0]),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(2) i_a3stg_rnd_mode (
        .din    (a2stg_rnd_mode[1:0]),
        .en     (a6stg_step),
        .clk    (rclk),
        .q      (a3stg_rnd_mode[1:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(5) i_a3stg_id (
        .din    (a2stg_id[4:0]),
        .en     (a6stg_step),
        .clk    (rclk),
        .q      (a3stg_id[4:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(2) i_a3stg_fcc (
        .din    (a2stg_fcc[1:0]),
        .en     (a6stg_step),
        .clk    (rclk),
        .q      (a3stg_fcc[1:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign a3stg_fadd= a3stg_opdec[34];
assign a3stg_int_dst= a3stg_opdec[30];
assign a3stg_faddsubop= a3stg_opdec[29];
assign a3stg_fsdtoix= a3stg_opdec_21;
assign a3stg_f4cycop= a3stg_opdec_9_0[8];
assign a3stg_fixtos_fxtod= a3stg_opdec_9_0[7];
assign a3stg_fdtos= a3stg_opdec_9_0[3];
dffre_s #(18) i_a4stg_opdec (
        .din    ({a3stg_opdec_36, a3stg_opdec[34:29], a3stg_opdec_24,
                  a3stg_opdec_21, a3stg_opdec_9_0[9], a3stg_opdec_9_0[7:0]}),
        .en     (a6stg_step),
        .rst    (reset),
        .clk    (rclk),
        .q      ({a4stg_opdec_36, a4stg_opdec[34:29], a4stg_opdec_24,
                  a4stg_opdec_21, a4stg_opdec_9, a4stg_opdec_7_0[7:0]}),
        .se     (se),
        .si     (),
        .so     ()
);
assign a4stg_rnd_mode_in[1:0]= ({2{a3stg_f4cycop}}
			    & a3stg_rnd_mode[1:0])
		| ({2{(!a3stg_f4cycop)}}
			    & a4stg_rnd_mode2[1:0]);
dffe_s #(2) i_a4stg_rnd_mode (
	.din	(a4stg_rnd_mode_in[1:0]),
	.en     (a6stg_step),
	.clk    (rclk),
        .q      (a4stg_rnd_mode[1:0]),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(2) i_a4stg_rnd_mode2 (
	.din	(a3stg_rnd_mode[1:0]),
	.en     (a6stg_step),
        .clk    (rclk),
 
        .q      (a4stg_rnd_mode2[1:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign a4stg_id_in[9:0]= {(a3stg_id[4:2]==3'o7),
				(a3stg_id[4:2]==3'o6),
				(a3stg_id[4:2]==3'o5),
				(a3stg_id[4:2]==3'o4),
				(a3stg_id[4:2]==3'o3),
				(a3stg_id[4:2]==3'o2),
				(a3stg_id[4:2]==3'o1),
				(a3stg_id[4:2]==3'o0),
				a3stg_id[1:0]};
dffe_s #(10) i_a4stg_id (
        .din    (a4stg_id_in[9:0]),
        .en     (a6stg_step),
        .clk    (rclk),
        .q      (a4stg_id[9:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(2) i_a4stg_fcc (
        .din    (a3stg_fcc[1:0]),
        .en     (a6stg_step),
        .clk    (rclk),
        .q      (a4stg_fcc[1:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign a4stg_dblop= a4stg_opdec_36;
assign a4stg_fadd= a4stg_opdec[34];
assign a4stg_faddsubop= a4stg_opdec[29];
assign a4stg_faddsub_dtosop= a4stg_opdec_24;
assign a4stg_fsdtoix= a4stg_opdec_21;
assign a4stg_fcmpop= a4stg_opdec_9;
assign a4stg_fixtos_fxtod= a4stg_opdec_7_0[7];
assign a4stg_faddsubs_fdtos= a4stg_opdec_7_0[6];
assign a4stg_faddsubs= a4stg_opdec_7_0[5];
assign a4stg_faddsubd= a4stg_opdec_7_0[4];
assign a4stg_fdtos= a4stg_opdec_7_0[3];
assign a4stg_fistod= a4stg_opdec_7_0[2];
dffre_s #(9) i_a5stg_opdec (
        .din    ({a4stg_opdec[34:30], a4stg_opdec_9, a4stg_opdec_7_0[7],
                  a4stg_opdec_7_0[1], a4stg_opdec_7_0[0]}),
        .en     (a6stg_step),
        .rst    (reset),
        .clk    (rclk),
        .q      ({a5stg_opdec[34:30], a5stg_opdec_9, a5stg_opdec_7,
                  a5stg_opdec_1, a5stg_opdec_0}),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(10) i_a5stg_id (
        .din    (a4stg_id[9:0]),
        .en     (a6stg_step),
        .clk    (rclk),
        .q      (a5stg_id[9:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign a5stg_fadd= a5stg_opdec[34];
assign a5stg_fixtos_fxtod= a5stg_opdec_7;
assign a5stg_fixtos= a5stg_opdec_1;
assign a5stg_fxtod= a5stg_opdec_0;
assign a6stg_opdec_in[34:30] = ({5{a5stg_fixtos_fxtod}}
			    & a5stg_opdec[34:30])
		| ({5{((!a4stg_fixtos_fxtod) && (!a5stg_fixtos_fxtod))}}
			    & a4stg_opdec[34:30]);
assign a6stg_opdec_in_9 = (a5stg_fixtos_fxtod
			    & a5stg_opdec_9)
		| (((!a4stg_fixtos_fxtod) && (!a5stg_fixtos_fxtod))
			    & a4stg_opdec_9);
assign a6stg_fadd_in= (a5stg_fixtos_fxtod && a6stg_step && (!reset)
			&& a5stg_fadd)
		|| ((!a4stg_fixtos_fxtod) && (!a5stg_fixtos_fxtod)
			&& a6stg_step && (!reset) && a4stg_fadd)
		|| ((!a6stg_step) && (!reset) && a6stg_fadd);
dffre_s #(6) i_a6stg_opdec (
	.din	({a6stg_opdec_in[34:30], a6stg_opdec_in_9}),
	.en     (a6stg_step),
        .rst    (reset),
        .clk    (rclk),
        .q      ({a6stg_opdec[34:30], a6stg_opdec_9}),
        .se     (se),
        .si     (),
        .so     ()
);
assign add_id_out_in[9:0]= ({10{((!a5stg_fixtos_fxtod) && a6stg_step)}}
			    & a4stg_id[9:0])
		| ({10{(a5stg_fixtos_fxtod && a6stg_step)}}
			    & a5stg_id[9:0])
		| ({10{(!a6stg_step)}}
			    & add_id_out[9:0]);
dff_s #(10) i_add_id_out (
	.din	(add_id_out_in[9:0]),
        .clk    (rclk),
        .q      (add_id_out[9:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign add_fcc_out_in[1:0]= ({2{a4stg_fcmpop}}
			    & a4stg_fcc);
dffe_s #(2) i_add_fcc_out (
	.din    (add_fcc_out_in[1:0]),
        .en     (a6stg_step),
        .clk    (rclk),
        .q      (add_fcc_out[1:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign a6stg_fadd= a6stg_opdec[34];
assign a6stg_dbl_dst= a6stg_opdec[33];
assign a6stg_sng_dst= a6stg_opdec[32];
assign a6stg_long_dst= a6stg_opdec[31];
assign a6stg_int_dst= a6stg_opdec[30];
assign a6stg_fcmpop= a6stg_opdec_9;
assign a6stg_hold= a6stg_fadd && (!add_dest_rdy);
assign a6stg_step= (!a6stg_hold);
assign add_pipe_active_in =  
   a1stg_fadd || a2stg_fadd || a3stg_fadd || a4stg_fadd || a5stg_fadd || a6stg_fadd;
dffre_s #(1) i_add_pipe_active (
	.din	(add_pipe_active_in),
	.en     (1'b1),
        .rst    (reset),
        .clk    (rclk),
        .q      (add_pipe_active),
        .se     (se),
        .si     (),
        .so     ()
);
assign a1stg_sub= (a1stg_fsubop ^ (a1stg_in1_63 ^ a1stg_in2_63))
		&& (!a1stg_fdtos)
		&& (!(a1stg_faddsubop && a1stg_nan_in));
dffe_s #(1) i_a2stg_sign1 (
	.din	(a1stg_in1_63),
	.en	(a6stg_step),
	.clk    (rclk),
        .q      (a2stg_sign1),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a2stg_sign2 (
	.din    (a1stg_in2_63),
        .en     (a6stg_step),
        .clk    (rclk),
 
        .q      (a2stg_sign2),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a2stg_sub (
        .din    (a1stg_sub),
        .en     (a6stg_step),
        .clk    (rclk),
 
        .q      (a2stg_sub),
 
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a2stg_in2_neq_in1_frac (
        .din    (a1stg_in2_neq_in1_frac),
        .en     (a6stg_step),
        .clk    (rclk),
 
        .q      (a2stg_in2_neq_in1_frac),
 
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a2stg_in2_gt_in1_frac (
        .din    (a1stg_in2_gt_in1_frac),
        .en     (a6stg_step),
        .clk    (rclk),
 
        .q      (a2stg_in2_gt_in1_frac),
 
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a2stg_in2_eq_in1_exp (
        .din    (a1stg_in2_eq_in1_exp),
        .en     (a6stg_step),
        .clk    (rclk),
 
        .q      (a2stg_in2_eq_in1_exp),
 
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a2stg_in2_gt_in1_exp (
        .din    (a1stg_expadd1[11]),
        .en     (a6stg_step),
        .clk    (rclk),
 
        .q      (a2stg_in2_gt_in1_exp),
 
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a2stg_nan_in (
        .din    (a1stg_nan_in),
        .en     (a6stg_step),
        .clk    (rclk),
 
        .q      (a2stg_nan_in),
 
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a2stg_nan_in2 (
        .din    (a1stg_nan_in2),
        .en     (a6stg_step),
        .clk    (rclk),
 
        .q      (a2stg_nan_in2),
 
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a2stg_snan_in2 (
        .din    (a1stg_snan_in2),
        .en     (a6stg_step),
        .clk    (rclk),
 
        .q      (a2stg_snan_in2),
 
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a2stg_qnan_in2 (
        .din    (a1stg_qnan_in2),
        .en     (a6stg_step),
        .clk    (rclk),
 
        .q      (a2stg_qnan_in2),
 
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a2stg_snan_in1 (
        .din    (a1stg_snan_in1),
        .en     (a6stg_step),
        .clk    (rclk),
 
        .q      (a2stg_snan_in1),
 
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a2stg_qnan_in1 (
        .din    (a1stg_qnan_in1),
        .en     (a6stg_step),
        .clk    (rclk),
 
        .q      (a2stg_qnan_in1),
 
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a2stg_2zero_in (
        .din    (a1stg_2zero_in),
        .en     (a6stg_step),
        .clk    (rclk),
 
        .q      (a2stg_2zero_in),
 
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a2stg_2inf_in (
        .din    (a1stg_2inf_in),
        .en     (a6stg_step),
        .clk    (rclk),
 
        .q      (a2stg_2inf_in),
 
        .se     (se),
        .si     (),
        .so     ()
);
assign a2stg_in2_eq_in1= a2stg_in2_eq_in1_exp && (!a2stg_in2_neq_in1_frac);
assign a2stg_in2_gt_in1= a2stg_in2_gt_in1_exp
		|| (a2stg_in2_eq_in1_exp && a2stg_in2_neq_in1_frac
			&& a2stg_in2_gt_in1_frac);
assign a3stg_sub_in= a2stg_sub
		&& (!a2stg_nan_in)
		&& (!(a2stg_fsdtoix && (!a2stg_expadd[11])));
assign a2stg_faddsub_sign= (a2stg_sign1
			&& (!a2stg_nan_in)
			&& (a2stg_sign2 ^ a2stg_fsubop)
			&& (!(a2stg_2inf_in && a2stg_sub)))
		|| (a2stg_sign1
			&& (!a2stg_nan_in)
			&& (!a2stg_in2_eq_in1)
			&& (!a2stg_in2_gt_in1)
			&& (!(a2stg_2inf_in && a2stg_sub)))
		|| ((!a2stg_in2_eq_in1)
			&& a2stg_in2_gt_in1
			&& (!a2stg_nan_in)
			&& (a2stg_sign2 ^ a2stg_fsubop)
			&& (!(a2stg_2inf_in && a2stg_sub)))
		|| (a2stg_sign2
			&& (a2stg_snan_in2
				|| (a2stg_qnan_in2 && (!a2stg_snan_in1))))
		|| (a2stg_sign1
			&& ((a2stg_snan_in1 && (!a2stg_snan_in2))
				|| (a2stg_qnan_in1 && (!a2stg_nan_in2))))
		|| ((a2stg_rnd_mode[1:0]==2'b11)
			&& a2stg_in2_eq_in1
			&& (a2stg_sign1 ^ (a2stg_sign2 ^ a2stg_fsubop))
			&& (!a2stg_nan_in)
			&& (!a2stg_2inf_in));
assign a3stg_sign_in= (a2stg_faddsubop && a2stg_faddsub_sign)
		|| ((!a2stg_faddsubop) && a2stg_sign2);
dffe_s #(1) i_a3stg_sign (
	.din	(a3stg_sign_in),
	.en     (a6stg_step),
        .clk    (rclk),
        .q      (a3stg_sign),
	.se     (se),
        .si     (),
        .so     ()
);
assign a2stg_cc_1= ((a2stg_sign2 && (!a2stg_2zero_in) && a2stg_sub)
			|| ((!a2stg_in2_eq_in1) && (!a2stg_sub)
				&& (a2stg_in2_gt_in1 ^ (!a2stg_sign2)))
			|| a2stg_nan_in)
		&& a2stg_fcmpop;
assign a2stg_cc_0= (((!a2stg_sign2) && (!a2stg_2zero_in) && a2stg_sub)
			|| ((!a2stg_in2_eq_in1) && (!a2stg_sub)
				&& (a2stg_in2_gt_in1 ^ a2stg_sign2))
			|| a2stg_nan_in)
		&& a2stg_fcmpop;
assign a2stg_cc[1:0]= {a2stg_cc_1, a2stg_cc_0};
dffe_s #(2) i_a3stg_cc (
	.din	(a2stg_cc[1:0]),
	.en     (a6stg_step),
        .clk    (rclk),
        .q      (a3stg_cc[1:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign a4stg_sign_in= (a3stg_f4cycop && a3stg_sign)
		|| ((!a3stg_f4cycop) && a4stg_sign2);
dffe_s #(1) i_a4stg_sign (
	.din	(a4stg_sign_in),
	.en     (a6stg_step),
        .clk    (rclk),
        .q      (a4stg_sign),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a4stg_sign2 (
	.din	(a3stg_sign),
	.en     (a6stg_step),
        .clk    (rclk),
        .q      (a4stg_sign2),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(2) i_a4stg_cc (
        .din    (a3stg_cc[1:0]),
        .en     (a6stg_step),
        .clk    (rclk),
        .q      (a4stg_cc[1:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_add_sign_out (
	.din	(a4stg_sign),
	.en     (a6stg_step),
        .clk    (rclk),
        .q      (add_sign_out),
	.se     (se),
        .si     (),
        .so     ()
);
assign add_cc_out_in[1:0]= ({2{a4stg_fcmpop}}
			    & a4stg_cc[1:0]);
dffe_s #(2) i_add_cc_out (
	.din	(add_cc_out_in[1:0]),
	.en     (a6stg_step),
        .clk    (rclk),
        .q      (add_cc_out[1:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign a1stg_nv= (a1stg_faddsubop
			&& ((a1stg_2inf_in && a1stg_sub)
				|| a1stg_snan_in1
				|| a1stg_snan_in2))
		|| (a1stg_fstod && a1stg_snan_in2)
		|| (a1stg_fdtos && a1stg_snan_in2)
		|| (a1stg_fcmpesd && a1stg_nan_in)
		|| (a1stg_fcmpsd
			&& (a1stg_snan_in1 || a1stg_snan_in2));
dffe_s #(1) i_a2stg_nv (
	.din	(a1stg_nv),
	.en     (a6stg_step),
        .clk    (rclk),
        .q      (a2stg_nv),
        .se     (se),
        .si     (),
        .so     ()
);
assign a1stg_of_mask= (!(a1stg_faddsub_dtosop && a1stg_infnan_in));
dffe_s #(1) i_a2stg_of_mask (
        .din    (a1stg_of_mask),
        .en     (a6stg_step),
        .clk    (rclk),
        .q      (a2stg_of_mask),
        .se     (se),
        .si     (),
        .so     ()
);
assign a3stg_nv_in= ((!a2stg_expadd[11])
			&& a2stg_fsdtoix
			&& ((!a2stg_sign2)
				|| (|a2stg_expadd[10:0])
				|| a2stg_frac2hi_neq_0
				|| (a2stg_long_dst && a2stg_frac2lo_neq_0)))
		|| a2stg_nv;
dffe_s #(1) i_a3stg_nv (
	.din	(a3stg_nv_in),
	.en     (a6stg_step),
        .clk    (rclk),
        .q      (a3stg_nv),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a3stg_of_mask (
        .din    (a2stg_of_mask),
        .en     (a6stg_step),
        .clk    (rclk),
        .q      (a3stg_of_mask),
        .se     (se),
        .si     (),
        .so     ()
);
assign a2stg_nx_tmp1= (a2stg_fdtoix && (|a2stg_exp[11:10]))
		|| (a2stg_fstoix && (|a2stg_exp[11:7]));
assign a2stg_nx_tmp2= ((a2stg_fdtoix && (!(|a2stg_exp[11:10])))
			|| (a2stg_fstoix && (!(|a2stg_exp[11:7]))))
		&& ((|a2stg_exp[10:1])
			|| a2stg_frac2hi_neq_0
			|| a2stg_frac2lo_neq_0
			|| a2stg_frac2_63);
assign a2stg_nx_tmp3= (a2stg_exp[11:0]==12'h41f)
		&& a2stg_sign2
		&& (!a2stg_frac2hi_neq_0)
		&& a2stg_frac2lo_neq_0
		&& a2stg_fdtoi;
dffe_s #(1) i_a3stg_a2_expadd_11 (
	.din	(a2stg_expadd[11]),
	.en	(a6stg_step),
	.clk	(rclk),
	.q	(a3stg_a2_expadd_11),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_a3stg_nx_tmp1 (
	.din	(a2stg_nx_tmp1),
	.en	(a6stg_step),
	.clk	(rclk),
	.q	(a3stg_nx_tmp1),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_a3stg_nx_tmp2 (
	.din	(a2stg_nx_tmp2),
	.en	(a6stg_step),
	.clk	(rclk),
	.q	(a3stg_nx_tmp2),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_a3stg_nx_tmp3 (
	.din	(a2stg_nx_tmp3),
	.en	(a6stg_step),
	.clk	(rclk),
	.q	(a3stg_nx_tmp3),
	.se	(se),
	.si	(),
	.so	()
);
assign a3stg_nx= (a3stg_a2_expadd_11
		    && ((a3stg_nx_tmp1
				&& ((a3stg_fsdtoi_nx && a3stg_int_dst)
					|| a3stg_fsdtoix_nx))
			|| a3stg_nx_tmp2))
		|| a3stg_nx_tmp3;
assign a4stg_nv_in= ((a3stg_fadd && (!a3stg_fixtos_fxtod))
			&& a3stg_nv)
		|| ((!(a3stg_fadd && (!a3stg_fixtos_fxtod)))
			&& a4stg_nv2);
dffe_s #(1) i_a4stg_nv (
        .din    (a4stg_nv_in),
        .en     (a6stg_step),
        .clk    (rclk),
        .q      (a4stg_nv),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a4stg_nv2 (
        .din    (a3stg_nv),
        .en     (a6stg_step),
        .clk    (rclk),
 
        .q      (a4stg_nv2),
 
        .se     (se),
        .si     (),
        .so     ()
);
assign a4stg_of_mask_in= ((a3stg_fadd && (!a3stg_fixtos_fxtod))
                        && a3stg_of_mask)
		|| ((!(a3stg_fadd && (!a3stg_fixtos_fxtod)))
                        && a4stg_of_mask2);
dffe_s #(1) i_a4stg_of_mask (
        .din    (a4stg_of_mask_in),
        .en     (a6stg_step),
        .clk    (rclk),
        .q      (a4stg_of_mask),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a4stg_of_mask2 (
        .din    (a3stg_of_mask),
        .en     (a6stg_step),
        .clk    (rclk),
 
        .q      (a4stg_of_mask2),
 
        .se     (se),
        .si     (),
        .so     ()
);
assign a4stg_nx_in= ((a3stg_fadd && (!a3stg_fixtos_fxtod))
                        && a3stg_nx)
                || ((!(a3stg_fadd && (!a3stg_fixtos_fxtod)))
                        && a4stg_nx2);
dffe_s #(1) i_a4stg_nx (
        .din    (a4stg_nx_in),
        .en     (a6stg_step),
        .clk    (rclk),
        .q      (a4stg_nx),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_a4stg_nx2 (
        .din    (a3stg_nx),
        .en     (a6stg_step),
        .clk    (rclk),
 
        .q      (a4stg_nx2),
 
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_add_nv_out (
        .din    (a4stg_nv),
        .en     (a6stg_step),
        .clk    (rclk),
        .q      (add_nv_out),
        .se     (se),
        .si     (),
        .so     ()
);
assign a4stg_in_of= ((a4stg_exp[11] || (&a4stg_exp[10:0]))
			&& a4stg_faddsubd
			&& a4stg_of_mask)
		|| (((|a4stg_exp[11:8]) || (&a4stg_exp[7:0]))
			&& a4stg_faddsubs_fdtos
			&& a4stg_of_mask);
assign add_of_out_tmp1_in= ((&a4stg_exp[10:1]) && a4stg_rndup && a4stg_round
			&& a4stg_faddsubd
                        && a4stg_of_mask)
		|| ((&a4stg_exp[7:1]) && a4stg_rndup
			&& (a4stg_round || a4stg_fdtos)
			&& a4stg_faddsubs_fdtos
			&& a4stg_of_mask);
dffe_s #(1) i_add_of_out_tmp1 (
        .din    (add_of_out_tmp1_in),
        .en     (a6stg_step),
        .clk    (rclk),
        .q      (add_of_out_tmp1),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_add_of_out_tmp2 (
	.din	(a4stg_in_of),
        .en	(a6stg_step),
        .clk	(rclk),
 
        .q	(add_of_out_tmp2),
 
        .se	(se),
        .si	(),
        .so	()
);
assign add_of_out= add_of_out_tmp2
		|| (add_of_out_tmp1 && add_of_out_cout);
assign a4stg_uf= ((!(|a4stg_exp[10:0]))
			&& a4stg_frac_neq_0
			&& (a4stg_round || a4stg_fdtos)
			&& a4stg_faddsub_dtosop)
		|| (a4stg_faddsubop
			&& (!(a4stg_round || a4stg_fdtos))
			&& (!a4stg_denorm_inv)
			&& a4stg_shl_data_neq_0);
dffe_s #(1) i_add_uf_out (
        .din    (a4stg_uf),
        .en     (a6stg_step),
        .clk    (rclk),
        .q      (add_uf_out),
        .se     (se),
        .si     (),
        .so     ()
);
assign add_nx_out_in= (a4stg_of_mask
			&& a4stg_frac_dbl_nx
			&& (a4stg_faddsubd || a5stg_fxtod)
			&& ((!a4stg_faddsubd) || a4stg_round))
		|| (a4stg_of_mask
			&& a4stg_frac_sng_nx
			&& (a4stg_faddsubs_fdtos || a5stg_fixtos)
			&& ((!a4stg_faddsubs) || a4stg_round))
		|| a4stg_nx;
dffe_s #(1) i_add_nx_out (
        .din    (add_nx_out_in),
        .en     (a6stg_step),
        .clk    (rclk),
        .q      (add_nx_out),
        .se     (se),
        .si     (),
        .so     ()
);
assign add_exc_out[4:0] =
  {add_nv_out,
   add_of_out,
   add_uf_out,
   1'b0,
   (add_nx_out || add_of_out)};  
 
assign a2stg_frac1_in_frac1= a1stg_snan_in2
		|| (a1stg_qnan_in2 && (!a1stg_snan_in1));
assign a2stg_frac1_in_frac2= a1stg_faddsubop
		&& ((!a1stg_2nan_in)
			|| a1stg_snan_in2
        		|| (a1stg_qnan_in2 && (!a1stg_snan_in1)));
assign a1stg_2nan_in_inv= (!a1stg_2nan_in);
assign a1stg_faddsubop_inv= (!a1stg_faddsubop);
assign a2stg_frac1_in_qnan= (a1stg_nan_in
			|| (a1stg_2inf_in && a1stg_sub))
		&& a1stg_faddsubop;
assign a2stg_frac1_in_nv= a1stg_2inf_in && a1stg_sub && a1stg_faddsubop;
assign a2stg_frac1_in_nv_dbl= a1stg_2inf_in && a1stg_sub && a1stg_faddsubd;
assign a2stg_frac2_in_frac1= a1stg_faddsubop && (!a1stg_infnan_in);
assign a2stg_frac2_in_qnan= a1stg_snan_in2 && (!a1stg_faddsubop);
assign a1stg_exp_diff_add1= a1stg_faddsub_dtosop && (!a1stg_expadd1[11]);
assign a1stg_exp_diff_add2= a1stg_faddsubop && a1stg_expadd1[11];
assign a1stg_exp_diff_5= (!a1stg_expadd2[5]) && a1stg_fsdtox;
assign a1stg_exp_diff[10:0]= ({11{a1stg_exp_diff_add1}}
			    & a1stg_expadd1[10:0])
		| ({11{a1stg_exp_diff_add2}}
			    & (~a1stg_expadd4_inv[10:0]))
		| ({11{a1stg_fsdtoix}}
			    & {5'b0, a1stg_exp_diff_5, (~a1stg_expadd2[4:0])});
assign a1stg_clamp63[5:0]= a1stg_exp_diff[5:0] | {6{(|a1stg_exp_diff[10:6])}};
assign a2stg_shr_cnt_in[5:0]= a1stg_clamp63[5:0];
assign a2stg_shr_cnt_5_inv_in= (!a1stg_clamp63[5]);
assign a2stg_shr_frac2_shr_int= a2stg_faddsub_dtosop && a6stg_step;
assign a2stg_shr_frac2_shr_dbl= ((a2stg_fdtox && (|a2stg_exp[11:10]))
			|| (a2stg_fstox && (|a2stg_exp[11:7])))
		&& a6stg_step;
assign a2stg_shr_frac2_shr_sng= ((a2stg_fdtoi && (|a2stg_exp[11:10]))
			|| (a2stg_fstoi && (|a2stg_exp[11:7])))
		&& a6stg_step;
assign a2stg_shr_frac2_max= a2stg_fsdtoix && a6stg_step;
assign a2stg_sub_step= a2stg_sub && a6stg_step;
assign a1stg_faddsub_clamp63_0= (|(({6{a1stg_expadd1[11]}}
			    & (~{a1stg_expadd4_inv[10:6],
						a1stg_expadd4_inv[0]}))
		| ({6{(!a1stg_expadd1[11])}}
			    & {a1stg_expadd1[10:6], a1stg_expadd1[0]})));
assign a2stg_fracadd_frac2_inv_in= (a1stg_fixtosd && a1stg_in2_63)
		|| (a1stg_faddsubop && a1stg_sub
			&& (!a1stg_faddsub_clamp63_0));
assign a2stg_fracadd_frac2_inv_shr1_in= a1stg_faddsubop && a1stg_sub
			&& a1stg_faddsub_clamp63_0;
assign a2stg_fracadd_frac2_in= (a1stg_fixtosd && (!a1stg_in2_63))
		|| a1stg_fstod
		|| (a1stg_faddsubop && (!a1stg_sub));
dffe_s #(1) i_a2stg_fracadd_frac2 (
	.din	(a2stg_fracadd_frac2_in),
	.en	(a6stg_step),
	.clk	(rclk),
	.q	(a2stg_fracadd_frac2),
	.se	(se),
	.si	(),
	.so   	()
);
assign a2stg_fracadd_cin_in= (a1stg_fixtosd && a1stg_in2_63)
		|| (a1stg_faddsubop && a1stg_sub);
assign a3stg_exp_7ff= a2stg_fstod && (&a2stg_exp[7:0]);
assign a3stg_exp_ff= a2stg_fdtos && (&a2stg_exp[10:0]);
assign a3stg_exp_add= (a2stg_fstod && (!(&a2stg_exp[7:0])))
		|| (a2stg_fdtos && (!(&a2stg_exp[10:0])));
assign a2stg_expdec_neq_0= a2stg_faddsubop && (a2stg_exp[10:0]<11'h36);
assign a3stg_exp10_0_eq0= (a3stg_exp[10:0]==11'b0);
assign a3stg_exp10_1_eq0= (a3stg_exp[10:1]==10'b0);
assign a3stg_fdtos_inv= (!a3stg_fdtos);
assign a4stg_fixtos_fxtod_inv= (!a4stg_fixtos_fxtod);
assign a4stg_rnd_frac_add_inv= (!(a3stg_fsdtoix
		|| (a3stg_faddsubop && a3stg_exp10_0_eq0)));
assign a4stg_shl_cnt_in[9:0]= ({10{a3stg_denorm}}
			    & {(a3stg_exp[5:4]==2'b11),
				(a3stg_exp[5:4]==2'b10),
				(a3stg_exp[5:4]==2'b01),
				(a3stg_exp[5:4]==2'b00),
				a3stg_exp[5:0]})
		| ({10{a3stg_denorm_inv}}
			    & {(a3stg_lead0[5:4]==2'b11),
				(a3stg_lead0[5:4]==2'b10),
				(a3stg_lead0[5:4]==2'b01),
				(a3stg_lead0[5:4]==2'b00),
				a3stg_lead0[5:0]});
assign a4stg_rnd_sng= a5stg_fixtos || a4stg_faddsubs_fdtos;
assign a4stg_rnd_dbl= a5stg_fxtod || a4stg_faddsubd;
	
assign a4stg_rndup_sng= ((a4stg_rnd_mode==2'b10) && (!a4stg_sign)
			&& a4stg_frac_sng_nx)
		|| ((a4stg_rnd_mode==2'b11) && a4stg_sign
			&& a4stg_frac_sng_nx)
		|| ((a4stg_rnd_mode==2'b00) && a4stg_rnd_frac_39
			&& (a4stg_frac_38_0_nx || a4stg_rnd_frac_40));
assign a4stg_rndup_dbl= ((a4stg_rnd_mode==2'b10) && (!a4stg_sign)
                        && a4stg_frac_dbl_nx)
                || ((a4stg_rnd_mode==2'b11) && a4stg_sign
                        && a4stg_frac_dbl_nx)
                || ((a4stg_rnd_mode==2'b00) && a4stg_rnd_frac_10
			&& (a4stg_frac_9_0_nx || a4stg_rnd_frac_11));
assign a4stg_rndup= (a4stg_faddsubd && a4stg_rndup_dbl)
		|| (a4stg_faddsubs && a4stg_rndup_sng)
		|| (a4stg_fdtos && a4stg_rndup_sng && a4stg_of_mask);
assign a5stg_rndup= (a5stg_fxtod && a4stg_rndup_dbl)
		|| (a5stg_fixtos && a4stg_rndup_sng);
assign add_frac_out_rndadd= (a4stg_faddsubop && a4stg_round && a4stg_rndup
			&& (!a4stg_in_of))
		|| (a4stg_fdtos && a4stg_rndup && (!a4stg_in_of))
		|| (a5stg_fixtos_fxtod && a5stg_rndup);
assign add_frac_out_rnd_frac= (a4stg_faddsubop && a4stg_round && (!a4stg_rndup)
			&& (!a4stg_in_of))
		|| (a4stg_fdtos && (!a4stg_rndup) && (!a4stg_in_of))
		|| (a5stg_fixtos_fxtod && (!a5stg_rndup))
		|| a4stg_fsdtoix;
assign add_frac_out_shl= (a4stg_faddsubop && (!a4stg_round) && (!a4stg_in_of))
		|| a4stg_fistod;
assign a4stg_to_0= (!((a4stg_rnd_mode==2'b00)
			|| ((a4stg_rnd_mode==2'b10) && (!a4stg_sign))
			|| ((a4stg_rnd_mode==2'b11) && a4stg_sign)));
assign add_exp_out_expinc= (a4stg_faddsubop && a4stg_round && a4stg_rndup
			&& (!a4stg_in_of))
		|| (a4stg_fdtos && a4stg_rndup
			&& (!a4stg_in_of))
		|| (a5stg_fixtos_fxtod && a5stg_rndup);
assign add_exp_out_exp= (a4stg_faddsubop && a4stg_round
			&& (!a4stg_in_of))
		|| (a4stg_fdtos
			&& (!a4stg_in_of))
		|| a5stg_fixtos_fxtod;
assign add_exp_out_exp1= (a4stg_faddsubop && a4stg_round
			&& (!a4stg_rndup)
			&& (!a4stg_in_of))
		|| (a4stg_fdtos
			&& (!a4stg_rndup)
			&& (!a4stg_in_of))
		|| (a5stg_fixtos_fxtod
			&& (!a5stg_rndup));
assign add_exp_out_expadd= (a4stg_faddsubop && (!a4stg_round) && (!a4stg_in_of))
		|| a4stg_fistod;
assign a4stg_to_0_inv= (!a4stg_to_0);
endmodule
module fpu_add_exp_dp (
	inq_in1,
	inq_in2,
	inq_op,
	inq_op_7,
	a1stg_step,
	a1stg_faddsubd,
	a1stg_faddsubs,
	a1stg_fsdtoix,
	a6stg_step,
	a1stg_fstod,
	a1stg_fdtos,
	a1stg_fstoi,
	a1stg_fstox,
	a1stg_fdtoi,
	a1stg_fdtox,
	a2stg_fsdtoix_fdtos,
	a2stg_faddsubop,
	a2stg_fitos,
	a2stg_fitod,
	a2stg_fxtos,
	a2stg_fxtod,
	a3stg_exp_7ff,
	a3stg_exp_ff,
	a3stg_exp_add,
	a3stg_inc_exp_inv,
	a3stg_same_exp_inv,
	a3stg_dec_exp_inv,
	a3stg_faddsubop,
	a3stg_fdtos_inv,
	a4stg_fixtos_fxtod_inv,
	a4stg_shl_cnt,
	a4stg_denorm_inv,
	a4stg_rndadd_cout,
	add_exp_out_expinc,
	add_exp_out_exp,
	add_exp_out_exp1,
	a4stg_in_of,
	add_exp_out_expadd,
	a4stg_dblop,
	a4stg_to_0_inv,
	fadd_clken_l,
	rclk,
	
	a1stg_expadd3_11,
	a1stg_expadd1_11_0,
	a1stg_expadd4_inv,
	a1stg_expadd2_5_0,
	a2stg_exp,
	a2stg_expadd,
	a3stg_exp_10_0,
	a4stg_exp_11_0,
	add_exp_out,
	se,
	si,
	so
);
input [62:52]	inq_in1;		
input [62:52]	inq_in2;		
input [1:0]	inq_op;			
input		inq_op_7;		
input		a1stg_step;		
input		a1stg_faddsubd;		
input		a1stg_faddsubs;		
input		a1stg_fsdtoix;		
input		a6stg_step;		
input		a1stg_fstod;		
input		a1stg_fdtos;		
input		a1stg_fstoi;		
input		a1stg_fstox;		
input		a1stg_fdtoi;		
input		a1stg_fdtox;		
input		a2stg_fsdtoix_fdtos;	
input		a2stg_faddsubop;	
input		a2stg_fitos;		
input		a2stg_fitod;		
input		a2stg_fxtos;		
input		a2stg_fxtod;		
input		a3stg_exp_7ff;		
input		a3stg_exp_ff;		
input		a3stg_exp_add;		
input		a3stg_inc_exp_inv;	
input		a3stg_same_exp_inv;	
input		a3stg_dec_exp_inv;	
input		a3stg_faddsubop;	
input		a3stg_fdtos_inv;	
input		a4stg_fixtos_fxtod_inv;	
input [5:0]	a4stg_shl_cnt;		
input		a4stg_denorm_inv;	
input		a4stg_rndadd_cout;	
input		add_exp_out_expinc;	
input		add_exp_out_exp;	
input		add_exp_out_exp1;	
input		a4stg_in_of;		
input		add_exp_out_expadd;	
input		a4stg_dblop;		
input		a4stg_to_0_inv;		
input		fadd_clken_l;           
input		rclk;		
output        	a1stg_expadd3_11;	
output [11:0]	a1stg_expadd1_11_0;	
output [10:0]	a1stg_expadd4_inv;	
output [5:0]	a1stg_expadd2_5_0;	
output [11:0]	a2stg_exp;		
output [12:0]	a2stg_expadd;		
output [10:0]	a3stg_exp_10_0;		
output [11:0]	a4stg_exp_11_0;		
output [10:0]	add_exp_out;		
input           se;                     
input           si;                     
output          so;                     
wire [62:52]	a1stg_in1;
wire [62:52]	a1stg_in1a;
wire [62:52]	a1stg_in2;
wire [62:52]	a1stg_in2a;
wire [12:0]	a1stg_dp_sngop;
wire [12:0]	a1stg_dp_sngopa;
wire [12:0]	a1stg_dp_dblop;
wire [12:0]	a1stg_dp_dblopa;
wire [9:7]      a1stg_op_7;
wire            a1stg_op_7_0;
wire [10:0]	a1stg_expadd3_in1;
wire [10:0]	a1stg_expadd3_in2_in;
wire [10:0]	a1stg_expadd3_in2;
wire [12:0]	a1stg_expadd3;
wire            a1stg_expadd3_11;
wire [12:0]	a1stg_expadd1_in1;
wire [12:0]	a1stg_expadd1_in2;
wire [12:0]	a1stg_expadd1;
wire [11:0]     a1stg_expadd1_11_0;
wire [12:0]	a1stg_expadd4_in1;
wire [12:0]	a1stg_expadd4_in2;
wire [12:0]	a1stg_expadd4;
wire [10:0]	a1stg_expadd4_inv;
wire [12:0]	a1stg_expadd2_in1;
wire [12:0]	a1stg_expadd2;
wire [5:0]      a1stg_expadd2_5_0;
wire [12:0]	a2stg_exp_in;
wire [11:0]	a2stg_exp;
wire [12:0]	a2stg_expa;
wire [12:0]	a2stg_expadd_in2_in;
wire [12:0]	a2stg_expadd_in2;
wire [12:0]	a2stg_expadd;
wire [12:0]	a3stg_exp_in;
wire [12:0]	a3stg_exp;
wire [10:0]     a3stg_exp_10_0;
wire [12:0]	a3stg_exp_plus1;
wire [12:0]	a3stg_exp_minus1;
wire [12:0]	a4stg_exp_pre1_in;
wire [12:0]	a4stg_exp_pre1;
wire [12:0]	a4stg_exp_pre3_in;
wire [12:0]	a4stg_exp_pre3;
wire [12:0]	a4stg_exp_pre2_in;
wire [12:0]	a4stg_exp_pre2;
wire [12:0]	a4stg_exp_pre4_in;
wire [12:0]	a4stg_exp_pre4;
wire [12:0]	a4stg_exp;
wire [11:0]	a4stg_exp_11_0;
wire [12:0]	a4stg_exp2;
wire [12:0]	a4stg_expinc;
wire [12:0]	a4stg_expadd_in2;
wire [12:0]	a4stg_expadd;
wire [12:0]	a4stg_expshl;
wire [10:0]	add_exp_out_in1;
wire [10:0]	add_exp_out1;
wire [10:0]	add_exp_out_in2;
wire [10:0]	add_exp_out2;
wire [10:0]	add_exp_out_in3;
wire [10:0]	add_exp_out3;
wire [10:0]	add_exp_out4;
wire [10:0]	add_exp_out;
wire        clk;
wire se_l;
assign se_l = ~se;
    clken_buf  ckbuf_add_exp_dp (
      .clk(clk),
      .rclk(rclk),
      .enb_l(fadd_clken_l),
      .tmb_l(se_l)
      );
dffe_s #(11) i_a1stg_in1 (
        .din    (inq_in1[62:52]),
        .en     (a1stg_step),
        .clk    (clk),
 
        .q      (a1stg_in1[62:52]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(11) i_a1stg_in1a (
	.din	(inq_in1[62:52]),
	.en	(a1stg_step),
	.clk	(clk),
	.q	(a1stg_in1a[62:52]),
	.se	(se),
        .si	(),
        .so	()
);
dffe_s #(11) i_a1stg_in2 (
	.din	(inq_in2[62:52]),
	.en	(a1stg_step),
	.clk	(clk),
	.q	(a1stg_in2[62:52]),
	.se	(se),
	.si	(),
   	.so	()
);
dffe_s #(11) i_a1stg_in2a (
        .din	(inq_in2[62:52]),
        .en	(a1stg_step),
        .clk	(clk),
 
        .q	(a1stg_in2a[62:52]),
 
        .se	(se),
        .si	(),
        .so	()
);
dffe_s #(13) i_a1stg_dp_sngop (
	.din	({13{inq_op[0]}}),
	.en	(a1stg_step),
	.clk	(clk),
	.q	(a1stg_dp_sngop[12:0]),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(13) i_a1stg_dp_sngopa (
        .din	({13{inq_op[0]}}),
        .en	(a1stg_step),
        .clk	(clk),
 
        .q	(a1stg_dp_sngopa[12:0]),
 
        .se	(se),
        .si	(),
        .so	()
);
dffe_s #(13) i_a1stg_dp_dblop (
	.din	({13{inq_op[1]}}),
	.en	(a1stg_step),
	.clk	(clk),
	.q	(a1stg_dp_dblop[12:0]),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(13) i_a1stg_dp_dblopa (
	.din	({13{inq_op[1]}}),
	.en	(a1stg_step),
	.clk	(clk),
	.q	(a1stg_dp_dblopa[12:0]),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(4) i_a1stg_op_7 (
	.din	({4{inq_op_7}}),
	.en	(a1stg_step),
	.clk	(clk),
	.q	({a1stg_op_7[9:7], a1stg_op_7_0}),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(11) i_a1stg_expadd3_in1 (
	.din	(inq_in1[62:52]),
	.en	(a1stg_step),
	.clk	(clk),
	.q	(a1stg_expadd3_in1[10:0]),
	.se	(se),
	.si	(),
	.so	()
);
assign a1stg_expadd3_in2_in[10:0]= (~(inq_in2[62:52] 
		& {8'hff, {3{inq_op[1]}}}));
dffe_s #(11) i_a1stg_expadd3_in2 (
	.din	(a1stg_expadd3_in2_in[10:0]),
	.en	(a1stg_step),
	.clk	(clk),
	.q	(a1stg_expadd3_in2[10:0]),
	.se	(se),
	.si	(),
	.so	()
);
assign a1stg_expadd3[12:0]= ({2'b00, a1stg_expadd3_in1[10:0]}
			+ {2'b11, a1stg_expadd3_in2[10:0]}
			+ 13'h0001);
assign a1stg_expadd3_11 = a1stg_expadd3[11];
assign a1stg_expadd1_in1[12:0]= (a1stg_dp_dblopa
			    & {2'b0, a1stg_in1[62:52]})
		| (a1stg_dp_sngopa
			    & {5'b0, a1stg_in1[62:55]})
		| {3'b0, a1stg_op_7[9:7], 6'b0, a1stg_op_7_0};
assign a1stg_expadd1_in2[12:0]= (~((a1stg_dp_dblop
			    & {2'b0, a1stg_in2[62:52]})
		| (a1stg_dp_sngop
			    & {5'b0, a1stg_in2[62:55]})));
assign a1stg_expadd1[12:0]= (a1stg_expadd1_in1[12:0]
			+ a1stg_expadd1_in2[12:0]
			+ 13'h0001);
assign a1stg_expadd1_11_0[11:0] = a1stg_expadd1[11:0];
assign a1stg_expadd4_in1[12:0]= (a1stg_dp_dblopa
			    & {2'b0, a1stg_in2a[62:52]})
                | (a1stg_dp_sngopa
			    & {5'b0, a1stg_in2a[62:55]});
assign a1stg_expadd4_in2[12:0]= (~((a1stg_dp_dblop
                            & {2'b0, a1stg_in1a[62:52]})
		| (a1stg_dp_sngop
			    & {5'b0, a1stg_in1a[62:55]})));
assign a1stg_expadd4[12:0]= (a1stg_expadd4_in1[12:0]
			+ a1stg_expadd4_in2[12:0]
			+ 13'h0001);
assign a1stg_expadd4_inv[10:0]= (~a1stg_expadd4[10:0]);
assign a1stg_expadd2_in1[12:0]= (a1stg_dp_dblopa
			    & {2'b0, a1stg_in2a[62:52]})
                | (a1stg_dp_sngopa
			    & {5'b0, a1stg_in2a[62:55]});
assign a1stg_expadd2[12:0]= (a1stg_expadd2_in1[12:0]
			+ 13'h0001);
assign a1stg_expadd2_5_0[5:0] = a1stg_expadd2[5:0];
assign a2stg_exp_in[12:0]= ({13{(a1stg_faddsubd && (!a1stg_expadd1[12]))}}
			    & {2'b0, a1stg_in1a[62:52]})
		| ({13{(a1stg_faddsubs && (!a1stg_expadd1[12]))}}
			    & {5'b0, a1stg_in1a[62:55]})
		| ({13{(a1stg_faddsubd && a1stg_expadd1[12])}}
			    & {2'b0, a1stg_in2[62:52]})
		| ({13{a1stg_fdtos}}
			    & {2'b0, a1stg_in2[62:52]})
		| ({13{(a1stg_faddsubs && a1stg_expadd1[12])}}
			    & {5'b0, a1stg_in2[62:55]})
		| ({13{a1stg_fstod}}
			    & {5'b0, a1stg_in2[62:55]})
		| ({13{a1stg_fsdtoix}}
			    & a1stg_expadd2[12:0]);
dffe_s #(12) i_a2stg_exp (
	.din	(a2stg_exp_in[11:0]),
	.en     (a6stg_step),
        .clk    (clk),
 
        .q      (a2stg_exp[11:0]),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(13) i_a2stg_expa (
	.din	(a2stg_exp_in[12:0]),
	.en	(a6stg_step),
	.clk	(clk),
	.q	(a2stg_expa[12:0]),
	.se	(se),
	.si	(),
	.so	()
);
assign a2stg_expadd_in2_in[12:0]= ({13{a1stg_fstod}}
			    & 13'h0380)
		| ({13{a1stg_fdtos}}
			    & (~13'h0380))
		| ({13{a1stg_fstoi}}
			    & (~13'h009f))
		| ({13{a1stg_fstox}}
			    & (~13'h00bf))
		| ({13{a1stg_fdtoi}}
			    & (~13'h041f))
		| ({13{a1stg_fdtox}}
			    & (~13'h043f));
dffe_s #(13) i_a2stg_expadd2_in2 (
        .din	(a2stg_expadd_in2_in[12:0]),
        .en	(a6stg_step),
        .clk	(clk),
 
        .q	(a2stg_expadd_in2[12:0]),
 
        .se	(se),
        .si	(),
        .so	()
);
assign a2stg_expadd[12:0]= (a2stg_expa[12:0]
			+ a2stg_expadd_in2[12:0]
			+ {12'b0, a2stg_fsdtoix_fdtos});
assign a3stg_exp_in[12:0]= ({13{a2stg_faddsubop}}
			    & a2stg_expa[12:0])
		| ({13{a2stg_fitos}}
			    & 13'h009e)
		| ({13{a2stg_fitod}}
			    & 13'h041e)
		| ({13{a2stg_fxtos}}
			    & 13'h00be)
		| ({13{a2stg_fxtod}}
			    & 13'h043e)
		| ({13{a3stg_exp_7ff}}
			    & 13'h07ff)
		| ({13{a3stg_exp_ff}}
			    & 13'h00ff)
		| ({13{a3stg_exp_add}}
			    & (a2stg_expadd[12:0] & {13{(!a2stg_expadd[11])}}));
dffe_s #(13) i_a3stg_exp (
        .din    (a3stg_exp_in[12:0]),
        .en     (a6stg_step),
        .clk    (clk),
 
        .q      (a3stg_exp[12:0]),
 
        .se     (se),
        .si     (),
        .so     ()
);
assign a3stg_exp_10_0[10:0] = a3stg_exp[10:0];
assign a3stg_exp_plus1[12:0]= a3stg_exp[12:0] + 13'h0001;
assign a3stg_exp_minus1[12:0]= a3stg_exp[12:0] - 13'h0001;
assign a4stg_exp_pre1_in[12:0]= ({13{(a3stg_faddsubop && a6stg_step
					&& (!a3stg_inc_exp_inv))}}
			    & a3stg_exp_plus1[12:0]);
dff_s #(13) i_a4stg_exp_pre1 (
	.din	(a4stg_exp_pre1_in[12:0]),
	.clk	(clk),
	.q	(a4stg_exp_pre1[12:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign a4stg_exp_pre3_in[12:0]= ({13{(a3stg_faddsubop && a6stg_step
					&& (!a3stg_dec_exp_inv))}}
			    & a3stg_exp_minus1[12:0]);
dff_s #(13) i_a4stg_exp_pre3 (
	.din	(a4stg_exp_pre3_in[12:0]),
	.clk	(clk),
	.q	(a4stg_exp_pre3[12:0]),
	.se	(se),
	.si	(),
	.so	()
);
assign a4stg_exp_pre2_in[12:0]= ({13{((!a3stg_fdtos_inv) && a6stg_step)}}
			    & a3stg_exp[12:0])
		| ({13{((!a4stg_fixtos_fxtod_inv) && a6stg_step)}}
			    & a4stg_expshl[12:0])
		| ({13{(!a6stg_step)}}
			    & a4stg_exp[12:0]);
dff_s #(13) i_a4stg_exp_pre2 (
	.din	(a4stg_exp_pre2_in[12:0]),
        .clk    (clk),
        .q      (a4stg_exp_pre2[12:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign a4stg_exp_pre4_in[12:0]= ({13{(a3stg_faddsubop && a6stg_step
					&& (!a3stg_same_exp_inv))}}
			    & a3stg_exp[12:0]);
dff_s #(13) i_a4stg_exp_pre4 (
	.din	(a4stg_exp_pre4_in[12:0]),
	.clk	(clk),
	.q	(a4stg_exp_pre4[12:0]),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(13) i_a4stg_exp2 (
	.din	(a3stg_exp[12:0]),
	.en     (a6stg_step),
        .clk    (clk),
        .q      (a4stg_exp2[12:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign a4stg_exp[12:0]= (a4stg_exp_pre1[12:0]
		| a4stg_exp_pre2[12:0]
		| a4stg_exp_pre3[12:0]
		| a4stg_exp_pre4[12:0]);
assign a4stg_exp_11_0[11:0] = a4stg_exp[11:0];
assign a4stg_expinc[12:0]= a4stg_exp[12:0] + 13'h0001;
assign a4stg_expadd_in2[12:0]= (~{7'b0, a4stg_shl_cnt[5:0]});
assign a4stg_expadd[12:0]= (a4stg_exp2[12:0]
			+ a4stg_expadd_in2[12:0]
			+ 13'h0001);
assign a4stg_expshl[12:0]= (a4stg_expadd[12:0] & {13{a4stg_denorm_inv}});
assign add_exp_out_in1[10:0]= (~(({11{add_exp_out_exp1}}
			    & a4stg_exp[10:0])
		| ({11{a4stg_in_of}}
			    & {{3{a4stg_dblop}}, 7'h7f, a4stg_to_0_inv})
		| ({11{add_exp_out_expadd}}
			    & a4stg_expshl[10:0])));
dffe_s #(11) i_add_exp_out1 (
	.din	(add_exp_out_in1[10:0]),
	.en     (a6stg_step),
        .clk    (clk),
        .q      (add_exp_out1[10:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign add_exp_out_in2[10:0]= (~({11{(add_exp_out_expinc
					&& a4stg_rndadd_cout)}}
			    & a4stg_expinc[10:0]));
dffe_s #(11) i_add_exp_out2 (
	.din	(add_exp_out_in2[10:0]),
	.en	(a6stg_step),
	.clk	(clk),
	.q	(add_exp_out2[10:0]),
	.se  	(se),
	.si	(),
	.so	()
);
assign add_exp_out_in3[10:0]= (~({11{add_exp_out_exp}}
			    & a4stg_exp[10:0]));
dffe_s #(11) i_add_exp_out3 (
	.din	(add_exp_out_in3[10:0]),
	.en	(a6stg_step),
	.clk	(clk),
	.q	(add_exp_out3[10:0]),
	.se  	(se),
	.si	(),
	.so	()
);
dffe_s #(11) i_add_exp_out4 (
	.din	({11{a4stg_rndadd_cout}}),
	.en	(a6stg_step),
	.clk	(clk),
	.q	(add_exp_out4[10:0]),
	.se  	(se),
	.si	(),
	.so	()
);
assign add_exp_out[10:0]= (~(add_exp_out1[10:0]
		& add_exp_out2[10:0]
		& (add_exp_out3[10:0] | add_exp_out4[10:0])));
endmodule
module fpu_add_frac_dp (
	inq_in1,
	inq_in2,
	a1stg_step,
	a1stg_sngop,
	a1stg_expadd3_11,
	a1stg_norm_dbl_in1,
	a1stg_denorm_dbl_in1,
	a1stg_norm_sng_in1,
	a1stg_denorm_sng_in1,
	a1stg_norm_dbl_in2,
	a1stg_denorm_dbl_in2,
	a1stg_norm_sng_in2,
	a1stg_denorm_sng_in2,
	a1stg_intlngop,
	a2stg_frac1_in_frac1,
	a2stg_frac1_in_frac2,
	a1stg_2nan_in_inv,
	a1stg_faddsubop_inv,
	a2stg_frac1_in_qnan,
	a2stg_frac1_in_nv,
	a2stg_frac1_in_nv_dbl,
	a6stg_step,
	a2stg_frac2_in_frac1,
	a2stg_frac2_in_qnan,
	a2stg_shr_cnt_in,
	a2stg_shr_cnt_5_inv_in,
	a2stg_shr_frac2_shr_int,
	a2stg_shr_frac2_shr_dbl,
	a2stg_shr_frac2_shr_sng,
	a2stg_shr_frac2_max,
	a2stg_expadd_11,
	a2stg_sub_step,
	a2stg_fracadd_frac2_inv_in,
	a2stg_fracadd_frac2_inv_shr1_in,
	a2stg_fracadd_frac2,
	a2stg_fracadd_cin_in,
	a2stg_exp,
	a2stg_expdec_neq_0,
	a3stg_faddsubopa,
	a3stg_sub_in,
	a3stg_exp10_0_eq0,
	a3stg_exp10_1_eq0,
	a3stg_exp_0,
	a4stg_rnd_frac_add_inv,
	a3stg_fdtos_inv,
	a4stg_fixtos_fxtod_inv,
	a4stg_rnd_sng,
	a4stg_rnd_dbl,
	a4stg_shl_cnt_in,
	add_frac_out_rndadd,
	add_frac_out_rnd_frac,
	a4stg_in_of,
	add_frac_out_shl,
	a4stg_to_0,
	fadd_clken_l,
	rclk,
	
	a1stg_in2_neq_in1_frac,
	a1stg_in2_gt_in1_frac,
	a1stg_in2_eq_in1_exp,
	a2stg_frac2_63,
	a2stg_frac2hi_neq_0,
	a2stg_frac2lo_neq_0,
	a3stg_fsdtoix_nx,
	a3stg_fsdtoi_nx,
	a3stg_denorm,
	a3stg_denorm_inv,
	a3stg_lead0,
	a4stg_round,
	a4stg_shl_cnt,
	a4stg_denorm_inv,
	a3stg_inc_exp_inv,
	a3stg_same_exp_inv,
	a3stg_dec_exp_inv,
	a4stg_rnd_frac_40,
	a4stg_rnd_frac_39,
	a4stg_rnd_frac_11,
	a4stg_rnd_frac_10,
	a4stg_rndadd_cout,
	a4stg_frac_9_0_nx,
	a4stg_frac_dbl_nx,
	a4stg_frac_38_0_nx,
	a4stg_frac_sng_nx,
	a4stg_frac_neq_0,
	a4stg_shl_data_neq_0,
	add_of_out_cout,
	add_frac_out,
	se,
        si,
        so
);
input [62:0]	inq_in1;		
input [63:0]	inq_in2;		
input		a1stg_step;		
input		a1stg_sngop;		
input		a1stg_expadd3_11;	
input		a1stg_norm_dbl_in1;	
input		a1stg_denorm_dbl_in1;	
input		a1stg_norm_sng_in1;	
input		a1stg_denorm_sng_in1;	
input		a1stg_norm_dbl_in2;	
input		a1stg_denorm_dbl_in2;	
input		a1stg_norm_sng_in2;	
input		a1stg_denorm_sng_in2;	
input		a1stg_intlngop;		
input		a2stg_frac1_in_frac1;	
input		a2stg_frac1_in_frac2;	
input		a1stg_2nan_in_inv;	
input		a1stg_faddsubop_inv;	
input		a2stg_frac1_in_qnan;	
input		a2stg_frac1_in_nv;	
input		a2stg_frac1_in_nv_dbl;	
input		a6stg_step;		
input		a2stg_frac2_in_frac1;	
input		a2stg_frac2_in_qnan;	
input [5:0]	a2stg_shr_cnt_in;	
input		a2stg_shr_cnt_5_inv_in;	
input		a2stg_shr_frac2_shr_int; 
input		a2stg_shr_frac2_shr_dbl; 
input		a2stg_shr_frac2_shr_sng; 
input		a2stg_shr_frac2_max;	
input		a2stg_expadd_11;	
input		a2stg_sub_step;		
input		a2stg_fracadd_frac2_inv_in; 
input		a2stg_fracadd_frac2_inv_shr1_in; 
input		a2stg_fracadd_frac2;	
input		a2stg_fracadd_cin_in;	
input [5:0]	a2stg_exp;		
input		a2stg_expdec_neq_0;	
input [1:0]	a3stg_faddsubopa;	
input		a3stg_sub_in;		
input		a3stg_exp10_0_eq0;	
input		a3stg_exp10_1_eq0;	
input		a3stg_exp_0;		
input		a4stg_rnd_frac_add_inv;	
input		a3stg_fdtos_inv;	
input		a4stg_fixtos_fxtod_inv;	
input		a4stg_rnd_sng;		
input		a4stg_rnd_dbl;		
input [9:0]	a4stg_shl_cnt_in;	
input		add_frac_out_rndadd;	
input		add_frac_out_rnd_frac;	
input		a4stg_in_of;		
input		add_frac_out_shl;	
input		a4stg_to_0;		
input		fadd_clken_l;           
input		rclk;		
output		a1stg_in2_neq_in1_frac;	
output		a1stg_in2_gt_in1_frac;	
output		a1stg_in2_eq_in1_exp;	
output		a2stg_frac2_63;		
output		a2stg_frac2hi_neq_0;	
output		a2stg_frac2lo_neq_0;	
output		a3stg_fsdtoix_nx;	
output		a3stg_fsdtoi_nx;	
output		a3stg_denorm;		
output		a3stg_denorm_inv;	
output [5:0]	a3stg_lead0;		
output		a4stg_round;		
output [5:0]	a4stg_shl_cnt;		
output		a4stg_denorm_inv;	
output		a3stg_inc_exp_inv;	
output		a3stg_same_exp_inv;	
output		a3stg_dec_exp_inv;	
output		a4stg_rnd_frac_40;	
output		a4stg_rnd_frac_39;	
output		a4stg_rnd_frac_11;	
output		a4stg_rnd_frac_10;	
output		a4stg_rndadd_cout;	
output		a4stg_frac_9_0_nx;	
output		a4stg_frac_dbl_nx;	
output		a4stg_frac_38_0_nx;	
output		a4stg_frac_sng_nx;	
output		a4stg_frac_neq_0;	
output		a4stg_shl_data_neq_0;	
output		add_of_out_cout;	
output [63:0]	add_frac_out;		
input           se;                     
input           si;                     
output          so;                     
wire [62:0]	a1stg_in1;
wire [54:0]	a1stg_in1a;
wire		a1stg_in1_31_0_neq_0;
wire		a1stg_in1_50_32_neq_0;
wire		a1stg_in1_50_0_neq_0;
wire		a1stg_in1_53_32_neq_0;
wire		a1stg_in1_51;
wire		a1stg_in1_54;
wire [63:0]	a1stg_in2;
wire [54:0]	a1stg_in2a;
wire		a1stg_in2_31_0_neq_0;
wire		a1stg_in2_50_32_neq_0;
wire		a1stg_in2_50_0_neq_0;
wire		a1stg_in2_53_32_neq_0;
wire		a1stg_in2_51;
wire		a1stg_in2_54;
wire		a1stg_in2_neq_in1_frac;
wire		a1stg_in2_gt_in1_frac;
wire		a1stg_in2_gt_in1;
wire		a1stg_in2_eq_in1_exp;
wire [63:0]	a1stg_norm_frac1;
wire [63:0]	a1stg_norm_frac2;
wire [63:0]	a2stg_frac1_in;
wire [63:0]	a2stg_frac1;
wire [63:0]	a2stg_frac2_in;
wire [63:0]	a2stg_frac2;
wire [63:0]	a2stg_frac2a;
wire		a2stg_frac2_63;
wire		a2stg_frac2hi_neq_0;
wire		a2stg_frac2lo_neq_0;
wire [115:52]	a2stg_shr;
wire		a2stg_fsdtoix_nx;
wire		a2stg_fsdtoi_nx;
wire		a2stg_shr_60_0_neq_0;
wire [63:0]	a2stg_shr_frac2_inv;
wire [63:0]	a3stg_frac2_in;
wire [63:0]	a3stg_frac2;
wire [63:0]	a3stg_frac1;
wire [63:0]	a2stg_fracadd_in2;
wire [63:0]	a2stg_fracadd;
wire [63:0]	a3stg_ld0_frac;
wire [53:0]	a2stg_expdec_tmp;
wire [53:0]	a2stg_expdec;
wire [53:0]	a3stg_expdec;
wire		a3stg_ld0_dnrm_10;
wire		a3stg_denorm;
wire		a3stg_denorm_inv;
wire		a3stg_denorma;
wire		a3stg_denorm_inva;
wire [5:0]	a3stg_lead0;
wire [63:0]	a3stg_fracadd;
wire		a4stg_round_in;
wire		a4stg_round;
wire [5:0]	a2stg_shr_cnt;
wire [5:3]	a2stg_shr_cnta;
wire [2:0]	a2stg_shr_cnta_5;
wire [3:0]	a2stg_shr_cnt_5_inv;
wire [3:0]	a2stg_shr_cnt_5;
wire [4:0]	a2stg_shr_cnt_4;
wire [4:0]	a2stg_shr_cnt_3;
wire [1:0]	a2stg_shr_cnt_2;
wire [1:0]	a2stg_shr_cnt_1;
wire [1:0]	a2stg_shr_cnt_0;
wire		a3stg_sub;
wire		a3stg_suba;
wire [2:0]	a4stg_shl_cnt_dec54_0;
wire [2:0]	a4stg_shl_cnt_dec54_1;
wire [2:0]	a4stg_shl_cnt_dec54_2;
wire [2:0]	a4stg_shl_cnt_dec54_3;
wire [5:0]	a4stg_shl_cnt;
wire		a2stg_fracadd_frac2_inv;
wire		a2stg_fracadd_frac2_inv_shr1;
wire		a4stg_denorm_inv;
wire		a3stg_fsdtoix_nx;
wire		a3stg_fsdtoi_nx;
wire		a2stg_fracadd_cin;
wire [63:0]	astg_xtra_regs;
wire		a3stg_inc_exp_inv;
wire		a3stg_same_exp_inv;
wire		a3stg_dec_exp_inv;
wire		a3stg_inc_exp_inva;
wire		a3stg_fsame_exp_inv;
wire		a3stg_fdec_exp_inv;
wire [63:0]	a4stg_rnd_frac_pre1_in;
wire [63:0]	a4stg_rnd_frac_pre1;
wire [63:0]	a4stg_rnd_frac_pre2_in;
wire [63:0]	a4stg_rnd_frac_pre2;
wire [63:0]	a4stg_rnd_frac_pre3_in;
wire [63:0]	a4stg_rnd_frac_pre3;
wire [63:0]	a4stg_rnd_frac;
wire [63:0]	a4stg_rnd_fraca;
wire		a4stg_rnd_frac_40;
wire		a4stg_rnd_frac_39;
wire		a4stg_rnd_frac_11;
wire		a4stg_rnd_frac_10;
wire [63:0]	a4stg_shl_data_in;
wire [63:0]	a4stg_shl_data;
wire [52:0]	a4stg_rndadd_tmp;
wire		a4stg_rndadd_cout;
wire [51:0]	a4stg_rndadd;
wire		a4stg_frac_9_0_nx;
wire		a4stg_frac_dbl_nx;
wire		a4stg_frac_38_0_nx;
wire		a4stg_frac_sng_nx;
wire		a4stg_frac_neq_0;
wire		a4stg_shl_data_neq_0;
wire [126:0]	a4stg_shl_tmp;
wire [63:0]	a4stg_shl;
wire		add_of_out_cout;
wire		a5stg_frac_out_rndadd;
wire		a5stg_frac_out_rnd_frac;
wire		a5stg_in_of;
wire		a5stg_frac_out_shl;
wire		a5stg_to_0;
wire [51:0]	a5stg_rndadd;
wire [63:0]	a5stg_rnd_frac;
wire [63:0]	a5stg_shl;
wire [63:0]	add_frac_out;
wire [63:0] a2stg_shr_tmp2;
wire [63:0] a2stg_shr_tmp4;
wire [63:0] a2stg_shr_tmp6;
wire [63:0] a2stg_shr_tmp8;
wire [63:0] a2stg_shr_tmp10;
wire [63:0] a2stg_shr_tmp13;
wire [63:0] a2stg_shr_tmp18;
wire [63:20] a2stg_nx_neq0_84_tmp_1;
wire [63:36] a2stg_nx_neq0_84_tmp_2;
wire [63:44] a2stg_nx_neq0_84_tmp_3;
wire [63:48] a2stg_nx_neq0_84_tmp_4;
wire [61:50] a2stg_nx_neq0_84_tmp_5;
wire [60:59] a2stg_nx_neq0_84_tmp_6;
wire a2stg_nx_neq0_84_tmp_6_51;
wire [63:0] a4stg_shl_tmp4;
wire se_l;
wire        clk;
assign se_l = ~se;
    clken_buf  ckbuf_add_frac_dp (
      .clk(clk),
      .rclk(rclk),
      .enb_l(fadd_clken_l),
      .tmb_l(se_l)
      );
dffe_s #(63) i_a1stg_in1 (
        .din    (inq_in1[62:0]),
        .en     (a1stg_step),
        .clk    (clk),
 
        .q      (a1stg_in1[62:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(55) i_a1stg_in1a (
        .din	(inq_in1[54:0]),
        .en	(a1stg_step),
        .clk	(clk),
 
        .q	(a1stg_in1a[54:0]),
 
        .se	(se),
        .si	(),
        .so	()
);
dffe_s #(64) i_a1stg_in2 (
        .din    (inq_in2[63:0]),
        .en     (a1stg_step),
        .clk    (clk),
 
        .q      (a1stg_in2[63:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(55) i_a1stg_in2a (
        .din	(inq_in2[54:0]),
        .en	(a1stg_step),
        .clk	(clk),
 
        .q	(a1stg_in2a[54:0]),
 
        .se	(se),
        .si	(),
        .so	()
);
fpu_in2_gt_in1_frac i_a1stg_in2_gt_in1_frac (
	.din1			(a1stg_in1a[54:0]),
	.din2			(a1stg_in2a[54:0]),
	.sngop			(a1stg_sngop),
	.expadd11		(a1stg_expadd3_11),
	.expeq			(a1stg_in2_eq_in1_exp),
	.din2_neq_din1		(a1stg_in2_neq_in1_frac),
	.din2_gt_din1		(a1stg_in2_gt_in1_frac),
	.din2_gt1_din1		(a1stg_in2_gt_in1)
);
assign a1stg_in2_eq_in1_exp= (&{(~(a1stg_in1[62:55] ^ a1stg_in2[62:55])),
				((~(a1stg_in1[54:52] ^ a1stg_in2[54:52]))
					| {3{a1stg_sngop}})});
assign a1stg_norm_frac1[63:0]= ({64{a1stg_norm_dbl_in1}}
			    & {1'b1, a1stg_in1[51:0], 11'b0})
		| ({64{a1stg_denorm_dbl_in1}}
			    & {a1stg_in1[51:0], 12'b0})
		| ({64{a1stg_norm_sng_in1}}
			    & {1'b1, a1stg_in1[54:32], 40'b0})
		| ({64{a1stg_denorm_sng_in1}}
			    & {a1stg_in1[54:32], 41'b0});
assign a1stg_norm_frac2[63:0]= ({64{a1stg_norm_dbl_in2}}
			    & {1'b1, a1stg_in2[51:0], 11'b0})
                | ({64{a1stg_denorm_dbl_in2}}
                            & {a1stg_in2[51:0], 12'b0})
                | ({64{a1stg_norm_sng_in2}} 
                            & {1'b1, a1stg_in2[54:32], 40'b0})
                | ({64{a1stg_denorm_sng_in2}}
                            & {a1stg_in2[54:32], 41'b0})
		| ({64{a1stg_intlngop}}
			    & a1stg_in2[63:0]);
assign a2stg_frac1_in[63:0]= ({64{(a1stg_faddsubop_inv
				|| (!((a1stg_in2_gt_in1 && a1stg_2nan_in_inv)
						|| a2stg_frac1_in_frac1)))}}
			    & {a1stg_norm_frac1[63],
				(a1stg_norm_frac1[62] || a2stg_frac1_in_qnan),
				(a1stg_norm_frac1[61:40]
						| {22{a2stg_frac1_in_nv}}),
				(a1stg_norm_frac1[39:11]
						| {29{a2stg_frac1_in_nv_dbl}}),
				a1stg_norm_frac1[10:0]})
		| ({64{(a2stg_frac1_in_frac2
				    && (a1stg_in2_gt_in1 || a2stg_frac1_in_frac1))}}
			    & {a1stg_norm_frac2[63],
				(a1stg_norm_frac2[62] || a2stg_frac1_in_qnan),
				(a1stg_norm_frac2[61:40]
						| {22{a2stg_frac1_in_nv}}),
				(a1stg_norm_frac2[39:11]
						| {29{a2stg_frac1_in_nv_dbl}}),
				a1stg_norm_frac2[10:0]});
dffe_s #(64) i_a2stg_frac1 (
	.din	(a2stg_frac1_in[63:0]),
	.en	(a6stg_step),
	.clk    (clk),
        .q      (a2stg_frac1[63:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign a2stg_frac2_in[63:0]= ({64{a1stg_faddsubop_inv}}
			    & {a1stg_norm_frac2[63],
				(a1stg_norm_frac2[62] || a2stg_frac2_in_qnan),
                                a1stg_norm_frac2[61:0]})
		| ({64{(a2stg_frac2_in_frac1 && (!a1stg_in2_gt_in1))}}
			    & {a1stg_norm_frac2[63],
        			(a1stg_norm_frac2[62] || a2stg_frac2_in_qnan),
        			a1stg_norm_frac2[61:0]})
		| ({64{(a2stg_frac2_in_frac1 && a1stg_in2_gt_in1)}}
			    & a1stg_norm_frac1[63:0]);
dffe_s #(64) i_a2stg_frac2 (
	.din	(a2stg_frac2_in[63:0]),
	.en	(a6stg_step),
	.clk    (clk),
        .q      (a2stg_frac2[63:0]),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(64) i_a2stg_frac2a (
	.din	(a2stg_frac2_in[63:0]),
	.en	(a6stg_step),
	.clk	(clk),
	.q	(a2stg_frac2a[63:0]),
	.se	(se),
	.si	(),
	.so	()
);
assign a2stg_frac2_63= a2stg_frac2[63];
assign a2stg_frac2hi_neq_0= (|a2stg_frac2[62:32]);
assign a2stg_frac2lo_neq_0= (|a2stg_frac2[31:11]);
assign a2stg_shr_tmp2[63:0] = ({{24{a2stg_shr_cnt_5[0]}}, {16{a2stg_shr_cnt_5[1]}}, {13{a2stg_shr_cnt_5[2]}}, {11{a2stg_shr_cnt_5[3]}}} & {32'h00000000, a2stg_frac2a[63:32]})
	| ({{24{a2stg_shr_cnt_5_inv[0]}}, {16{a2stg_shr_cnt_5_inv[1]}}, {13{a2stg_shr_cnt_5_inv[2]}}, {11{a2stg_shr_cnt_5_inv[3]}}} & a2stg_frac2a[63:0]);
assign a2stg_shr_tmp4[63:0] = ({{24{a2stg_shr_cnt_4[0]}}, {16{a2stg_shr_cnt_4[1]}}, {13{a2stg_shr_cnt_4[2]}}, {11{a2stg_shr_cnt_4[3]}}} & {16'h0000, a2stg_shr_tmp2[63:16]})
	| ({{43{~a2stg_shr_cnt_4[4]}}, {21{~a2stg_shr_cnt_4[4]}}} & a2stg_shr_tmp2[63:0]);
assign a2stg_shr_tmp6[63:0] = ~(({{24{a2stg_shr_cnt_3[0]}}, {16{a2stg_shr_cnt_3[1]}}, {13{a2stg_shr_cnt_3[2]}}, {11{a2stg_shr_cnt_3[3]}}} & {8'h00, a2stg_shr_tmp4[63:8]})
	| ({64{~a2stg_shr_cnt_3[4]}} & a2stg_shr_tmp4[63:0]));
assign a2stg_shr_tmp8[63:0] = ~(({{43{a2stg_shr_cnt_2[0]}}, {21{a2stg_shr_cnt_2[0]}}} | a2stg_shr_tmp6[63:0])
	& ({64{~a2stg_shr_cnt_2[1]}} | {4'hf, a2stg_shr_tmp6[63:4]}));
assign a2stg_shr_tmp10[63:0] = ~(({{43{a2stg_shr_cnt_1[0]}}, {21{a2stg_shr_cnt_1[0]}}} & {2'b00, a2stg_shr_tmp8[63:2]})
	| ({64{~a2stg_shr_cnt_1[1]}} & a2stg_shr_tmp8[63:0]));
assign a2stg_shr[115:52] = ~(({{43{a2stg_shr_cnt_0[0]}}, {21{a2stg_shr_cnt_0[0]}}} | a2stg_shr_tmp10[63:0])
	 & ({64{~a2stg_shr_cnt_0[1]}} | {1'b1, a2stg_shr_tmp10[63:1]}));
assign a2stg_shr_tmp18[63:0] = ~a2stg_shr_tmp2[63:0];
assign a2stg_shr_tmp13[63:0] = a2stg_shr_tmp4[63:0];
assign a2stg_fsdtoi_nx = (| a2stg_shr_tmp13[31:0])
	| (~(& a2stg_shr_tmp6[31:24]))
	| (| a2stg_shr_tmp8[31:28])
	| (~(& a2stg_shr_tmp10[31:30]))
	| a2stg_shr[83];
assign a2stg_nx_neq0_84_tmp_1[63:20] = ~((a2stg_frac2a[43:0] & {44{a2stg_shr_cnt[5]}})
	| ({a2stg_frac2a[11:0], 32'h00000000} & {44{~a2stg_shr_cnt[5]}}));
assign a2stg_nx_neq0_84_tmp_2[63:36] = ~(({a2stg_shr_tmp18[27:12], a2stg_nx_neq0_84_tmp_1[63:52]} | {28{~a2stg_shr_cnt[4]}})
	& (a2stg_nx_neq0_84_tmp_1[63:36] | {28{a2stg_shr_cnt[4]}}));
assign a2stg_nx_neq0_84_tmp_3[63:44] = ~(({a2stg_shr_tmp13[19:12], a2stg_nx_neq0_84_tmp_2[63:52]} & {20{a2stg_shr_cnt[3]}})
	| (a2stg_nx_neq0_84_tmp_2[63:44] & {20{~a2stg_shr_cnt[3]}}));
assign a2stg_nx_neq0_84_tmp_4[63:48] = ~(({a2stg_shr_tmp6[15:12], a2stg_nx_neq0_84_tmp_3[63:52]} | {16{~a2stg_shr_cnt[2]}})
	& (a2stg_nx_neq0_84_tmp_3[63:48] | {16{a2stg_shr_cnt[2]}}));
assign a2stg_nx_neq0_84_tmp_5[61:50] = ~((a2stg_nx_neq0_84_tmp_4[63:52] & {12{a2stg_shr_cnt[1]}})
	| (a2stg_nx_neq0_84_tmp_4[61:50] & {12{~a2stg_shr_cnt[1]}}));
assign a2stg_nx_neq0_84_tmp_6[59] = ~(a2stg_shr_cnt[0] | a2stg_nx_neq0_84_tmp_5[60]);
assign a2stg_nx_neq0_84_tmp_6[60] = ~(~a2stg_shr_cnt[0] | a2stg_nx_neq0_84_tmp_5[61]);
assign a2stg_nx_neq0_84_tmp_6_51 = ~((a2stg_nx_neq0_84_tmp_5[52] | ~a2stg_shr_cnt[0])
	& (a2stg_nx_neq0_84_tmp_5[51] | a2stg_shr_cnt[0]));
assign a2stg_fsdtoix_nx = (~(& a2stg_nx_neq0_84_tmp_1[51:20])
	| (| a2stg_nx_neq0_84_tmp_2[51:36])
	| ~(& a2stg_nx_neq0_84_tmp_3[51:44])
	| (| a2stg_nx_neq0_84_tmp_4[51:48])
	| ~(& a2stg_nx_neq0_84_tmp_5[51:50])
	| a2stg_nx_neq0_84_tmp_6_51);
assign a2stg_shr_60_0_neq_0 = (~(& a2stg_nx_neq0_84_tmp_1[60:20])
	| (| a2stg_nx_neq0_84_tmp_2[60:45])
	| ~(& a2stg_nx_neq0_84_tmp_3[60:53])
	| (| a2stg_nx_neq0_84_tmp_4[60:57])
	| ~(& a2stg_nx_neq0_84_tmp_5[60:59])
	| (| a2stg_nx_neq0_84_tmp_6[60:59]));
assign a2stg_shr_frac2_inv[63:0]= (~(({64{a2stg_shr_frac2_shr_int}}
			    & {1'b0, a2stg_shr[115:61], a2stg_shr_60_0_neq_0,
					7'b0})
		| ({64{(a2stg_shr_frac2_shr_dbl && a2stg_expadd_11)}}
			    & a2stg_shr[115:52])
		| ({64{(a2stg_shr_frac2_shr_sng && a2stg_expadd_11)}}
			    & {a2stg_shr[115:84], 32'b0})
		| ({64{(a2stg_shr_frac2_max && (!a2stg_expadd_11))}}
			    & 64'h7fffffffffffffff)
		| ({64{(!a6stg_step)}}
			    & a3stg_frac2[63:0])));
assign a3stg_frac2_in[63:0]= (~(a2stg_shr_frac2_inv[63:0]
		^ {64{a2stg_sub_step}}));
dff_s #(64) i_a3stg_frac2 (
	.din	(a3stg_frac2_in[63:0]),
        .clk    (clk),
        .q      (a3stg_frac2[63:0]),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(64) i_a3stg_frac1 (
	.din    ({1'b0, a2stg_frac1[63:1]}),
	.en     (a6stg_step),
        .clk    (clk),
        .q      (a3stg_frac1[63:0]),
         
        .se     (se),
        .si     (),
        .so     ()
);
assign a2stg_fracadd_in2[63:0]= ({64{a2stg_fracadd_frac2_inv}}
			    & (~a2stg_frac2[63:0]))
		| ({64{a2stg_fracadd_frac2_inv_shr1}}
			    & (~{1'b0, a2stg_frac2[63:1]}))
		| ({64{a2stg_fracadd_frac2}}
			    & a2stg_frac2[63:0]);
assign a2stg_fracadd[63:0]= (a2stg_frac1[63:0]
			+ a2stg_fracadd_in2[63:0]
			+ {63'b0, a2stg_fracadd_cin});
dffe_s #(64) i_a3stg_ld0_frac (
	.din	(a2stg_fracadd[63:0]),
	.en     (a6stg_step),
        .clk    (clk),
        .q      (a3stg_ld0_frac[63:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign a2stg_expdec_tmp[53:0] =          54'h20000000000000  >> a2stg_exp[5:0] ;
assign a2stg_expdec[53:0]= a2stg_expdec_tmp[53:0] & {54{a2stg_expdec_neq_0}};
dffe_s #(54) i_a3stg_expdec (
	.din	(a2stg_expdec[53:0]),
	.en     (a6stg_step),
        .clk    (clk),
        .q      (a3stg_expdec[53:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign a3stg_ld0_dnrm_10= (a3stg_faddsubopa[0] && a3stg_ld0_frac[10])
		|| ((!a3stg_faddsubopa[0]) && (|a3stg_ld0_frac[10:0]));
fpu_denorm_frac i_a3stg_denorm (
	.din1			({a3stg_ld0_frac[63:11], a3stg_ld0_dnrm_10}),
	.din2			(a3stg_expdec[53:0]),
	.din2_din1_denorm	(a3stg_denorm),
	.din2_din1_denorm_inv	(a3stg_denorm_inv),
	.din2_din1_denorma	(a3stg_denorma),
	.din2_din1_denorm_inva	(a3stg_denorm_inva)
);
fpu_cnt_lead0_64b i_a3stg_lead0 (
	.din	(a3stg_ld0_frac[63:0]),
	.lead0	(a3stg_lead0[5:0])
);
assign a3stg_fracadd[63:0]= (a3stg_frac1[63:0]
			+ a3stg_frac2[63:0]
			+ {63'b0, a3stg_suba});
dffe_s #(64) i_astg_xtra_regs (
	.din	({{4{a2stg_shr_cnt_5_inv_in}}, {4{a2stg_shr_cnt_in[5]}},
			a2stg_shr_cnt_in[5:3],
			{5{a2stg_shr_cnt_in[4]}}, {5{a2stg_shr_cnt_in[3]}},
			a2stg_shr_cnt_in[5:0], a4stg_round_in,
			{2{a2stg_shr_cnt_in[2]}}, {2{a2stg_shr_cnt_in[1]}},
			{2{a2stg_shr_cnt_in[0]}},
			{3{a4stg_shl_cnt_in[6]}},
			{3{a4stg_shl_cnt_in[7]}},
			{3{a4stg_shl_cnt_in[8]}},
			{3{a4stg_shl_cnt_in[9]}},
			a4stg_shl_cnt_in[5:0],
			{3{a2stg_shr_cnt_in[5]}},
			a2stg_fracadd_frac2_inv_in,
			a2stg_fracadd_frac2_inv_shr1_in,
			a3stg_denorm_inva,
			a2stg_fsdtoix_nx, a2stg_fsdtoi_nx,
			1'b0, a2stg_fracadd_cin_in, {2{a3stg_sub_in}}}),
	.en	(a6stg_step),
	.clk	(clk),
	.q	({a2stg_shr_cnt_5_inv[3:0], a2stg_shr_cnt_5[3:0],
			a2stg_shr_cnta[5:3],
			a2stg_shr_cnt_4[4:0], a2stg_shr_cnt_3[4:0],
			a2stg_shr_cnt[5:0], a4stg_round,
			a2stg_shr_cnt_2[1:0], a2stg_shr_cnt_1[1:0],
			a2stg_shr_cnt_0[1:0],
			a4stg_shl_cnt_dec54_0[2:0],
			a4stg_shl_cnt_dec54_1[2:0],
			a4stg_shl_cnt_dec54_2[2:0],
			a4stg_shl_cnt_dec54_3[2:0],
			a4stg_shl_cnt[5:0],
			a2stg_shr_cnta_5[2:0],
			a2stg_fracadd_frac2_inv,
			a2stg_fracadd_frac2_inv_shr1,
			a4stg_denorm_inv,
			a3stg_fsdtoix_nx, a3stg_fsdtoi_nx,
			astg_xtra_regs[3], a2stg_fracadd_cin,
			a3stg_sub, a3stg_suba}),
	.se     (se),
        .si     (),
        .so     ()
);
assign a4stg_round_in= a3stg_fracadd[61]
		|| a3stg_fracadd[62]
		|| a3stg_fracadd[63];
assign a3stg_inc_exp_inv= (!a3stg_fracadd[63]);
assign a3stg_same_exp_inv= (!(((!a3stg_fracadd[63]) && a3stg_fracadd[62])
		|| ((!a3stg_fracadd[63]) && a3stg_exp10_0_eq0)));
assign a3stg_dec_exp_inv= (!((!a3stg_fracadd[63])
		&& (!a3stg_fracadd[62])
		&& a3stg_fracadd[61]
		&& (!a3stg_exp10_0_eq0)));
assign a3stg_inc_exp_inva= (!a3stg_fracadd[63]);
assign a3stg_fsame_exp_inv= (!(((!a3stg_fracadd[63])
			&& (!a3stg_fracadd[62])
			&& a3stg_fracadd[61]
			&& a3stg_exp10_1_eq0
			&& a3stg_exp_0)
		|| ((!a3stg_fracadd[63])
			&& a3stg_fracadd[62]
			&& (!a3stg_exp10_0_eq0))));
assign a3stg_fdec_exp_inv= (!((!a3stg_fracadd[63])
		&& (!a3stg_fracadd[62])
		&& a3stg_fracadd[61]
		&& (!a3stg_exp10_1_eq0)));
assign a4stg_rnd_frac_pre1_in[63:0]= ({64{(a3stg_faddsubopa[1] && a6stg_step
					&& (!a3stg_fdec_exp_inv))}}
			    & {a3stg_fracadd[61:0], 2'b00});
dff_s #(64) i_a4stg_rnd_frac_pre1 (
	.din	(a4stg_rnd_frac_pre1_in[63:0]),
        .clk    (clk),
        .q      (a4stg_rnd_frac_pre1[63:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign a4stg_rnd_frac_pre3_in[63:0]= ({64{(a3stg_faddsubopa[1] && a6stg_step
					&& (!a3stg_fsame_exp_inv))}}
			    & {a3stg_fracadd[62:0], 1'b0});
dff_s #(64) i_a4stg_rnd_frac_pre3 (
	.din	(a4stg_rnd_frac_pre3_in[63:0]),
        .clk    (clk),
        .q      (a4stg_rnd_frac_pre3[63:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign a4stg_rnd_frac_pre2_in[63:0]= ({64{(a3stg_faddsubopa[1] && a6stg_step
					&& (!a3stg_inc_exp_inva))}}
			    & a3stg_fracadd[63:0])
		| ({64{((!a4stg_rnd_frac_add_inv) && a6stg_step)}}
			    & a3stg_fracadd[63:0])
		| ({64{((!a3stg_fdtos_inv) && a6stg_step)}}
			    & {a3stg_fracadd[62:0], 1'b0})
		| ({64{((!a4stg_fixtos_fxtod_inv) && a6stg_step)}}
			    & a4stg_shl[63:0])
		| ({64{(!a6stg_step)}}
			    & a4stg_rnd_frac[63:0]);
dff_s #(64) i_a4stg_rnd_frac_pre2 (
	.din	(a4stg_rnd_frac_pre2_in[63:0]),
        .clk    (clk),
        .q      (a4stg_rnd_frac_pre2[63:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign a4stg_shl_data_in[63:0]= ({64{a3stg_denorm_inva}}
			    & a3stg_ld0_frac[63:0])
		| ({64{a3stg_denorma}}
			    & {1'b0, a3stg_ld0_frac[63:1]});
dffe_s #(64) i_a4stg_shl_data (
	.din	(a4stg_shl_data_in[63:0]),
	.en     (a6stg_step),
        .clk    (clk),
        .q      (a4stg_shl_data[63:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign a4stg_rnd_frac[63:0]= (a4stg_rnd_frac_pre1[63:0]
				| a4stg_rnd_frac_pre2[63:0]
				| a4stg_rnd_frac_pre3[63:0]);
assign a4stg_rnd_frac_40= a4stg_rnd_frac[40];
assign a4stg_rnd_frac_39= a4stg_rnd_frac[39];
assign a4stg_rnd_frac_11= a4stg_rnd_frac[11];
assign a4stg_rnd_frac_10= a4stg_rnd_frac[10];
assign a4stg_frac_9_0_nx= (|a4stg_rnd_frac[9:0]);
assign a4stg_frac_dbl_nx= a4stg_frac_9_0_nx || a4stg_rnd_frac[10];
assign a4stg_frac_38_0_nx= a4stg_frac_dbl_nx || (|a4stg_rnd_frac[38:11]);
assign a4stg_frac_sng_nx= a4stg_frac_38_0_nx || a4stg_rnd_frac[39];
assign a4stg_frac_neq_0= a4stg_frac_sng_nx || (|a4stg_rnd_frac[63:40]);
assign a4stg_rndadd_tmp[52:0]= {1'b0, a4stg_rnd_frac[62:11]}
			+ {23'b0, a4stg_rnd_sng, 28'b0, a4stg_rnd_dbl};
assign a4stg_rndadd_cout= a4stg_rndadd_tmp[52];
assign a4stg_rndadd[51:0]= a4stg_rndadd_tmp[51:0];
assign a4stg_shl_data_neq_0= (|a4stg_shl_data[63:0]);
assign a4stg_shl_tmp4[63:0] = ({{32{a4stg_shl_cnt_dec54_0[0]}}, {21{a4stg_shl_cnt_dec54_0[1]}}, {11{a4stg_shl_cnt_dec54_0[2]}}} & a4stg_shl_data[63:0])
	| ({{32{a4stg_shl_cnt_dec54_1[0]}}, {21{a4stg_shl_cnt_dec54_1[1]}}, {11{a4stg_shl_cnt_dec54_1[2]}}} & {a4stg_shl_data[47:0], 16'h0000})
	| ({{32{a4stg_shl_cnt_dec54_2[0]}}, {21{a4stg_shl_cnt_dec54_2[1]}}, {11{a4stg_shl_cnt_dec54_2[2]}}} & {a4stg_shl_data[31:0], 32'h00000000})
	| ({{32{a4stg_shl_cnt_dec54_3[0]}}, {21{a4stg_shl_cnt_dec54_3[1]}}, {11{a4stg_shl_cnt_dec54_3[2]}}} & {a4stg_shl_data[15:0], 32'h00000000, 16'h0000});
assign a4stg_shl[63:0] = a4stg_shl_tmp4[63:0] << a4stg_shl_cnt[3:0];
dffe_s #(58) i_a5stg_rndadd (
	.din	({a4stg_rndadd_cout, add_frac_out_rndadd, add_frac_out_rnd_frac,
			a4stg_in_of, add_frac_out_shl, a4stg_to_0,
			a4stg_rndadd[51:0]}),
	.en	(a6stg_step),
        .clk    (clk),
	.q	({add_of_out_cout, a5stg_frac_out_rndadd,
			a5stg_frac_out_rnd_frac, a5stg_in_of,
			a5stg_frac_out_shl, a5stg_to_0,
			a5stg_rndadd[51:0]}),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(64) i_a5stg_rnd_frac (
	.din	(a4stg_rnd_frac[63:0]),
	.en	(a6stg_step),
	.clk	(clk),
	.q	(a5stg_rnd_frac[63:0]),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(64) i_a5stg_shl (
	.din	(a4stg_shl[63:0]),
	.en	(a6stg_step),
	.clk	(clk),
	.q	(a5stg_shl[63:0]),
	.se	(se),
	.si	(),
	.so	()
);
assign add_frac_out[63:0]= ({64{a5stg_frac_out_rndadd}}
			    & {1'b0, a5stg_rndadd[51:0], 11'b0})
		| ({64{a5stg_frac_out_rnd_frac}}
			    & a5stg_rnd_frac[63:0])
		| ({64{a5stg_in_of}}
			    & {64{a5stg_to_0}})
		| ({64{a5stg_frac_out_shl}}
			    & a5stg_shl[63:0]);
endmodule
module fpu_arb (
	arst_l,
	grst_l,
	gclk,
	cluster_cken,
    
	pcx_fpio_data_rdy_px1,
    pcx_fpio_data_rdy_squashed,
	pcx_fpio_data_px2,
    l15_fp_rdy,
    
	fpu_arb_data_rdy,
	fpu_arb_data,
	fpu_arb_grant,
	ctu_tst_pre_grst_l,
	global_shift_enable,
	ctu_tst_scan_disable,
	ctu_tst_scanmode,
	ctu_tst_macrotest,
	ctu_tst_short_chain,
	si,
	so
);
input		    arst_l;			
input		    grst_l;			
input		    gclk;			
input		    cluster_cken;			
input		    pcx_fpio_data_rdy_px1;	
input           pcx_fpio_data_rdy_squashed;  
input [123:0]	pcx_fpio_data_px2;	
input           l15_fp_rdy;
input			ctu_tst_pre_grst_l;
input			global_shift_enable;
input			ctu_tst_scan_disable;
input			ctu_tst_scanmode;
input 			ctu_tst_macrotest;
input 			ctu_tst_short_chain;
input           si;                     
output      	fpu_arb_data_rdy;		
output [144:0]	fpu_arb_data;		
output reg      fpu_arb_grant;
output          so;                     
wire [7:0]   fp_cpx_req_cq;
wire [144:0] fp_cpx_data_ca;
reg pcx_fpio_data_rdy_px2;
reg is_fp;
always @*
begin
    is_fp = pcx_fpio_data_px2[122:119] == 4'b0101;
    pcx_fpio_data_rdy_px2 = pcx_fpio_data_px2[123] && is_fp;
    
    
    
    fpu_arb_grant = 1'b0;
    
end
always @(posedge gclk)
begin
    if (~grst_l)
    begin
        
        
        
    end
    else
    begin
        
        
        
        
        
    end
end
fpu fpu (
    .pcx_fpio_data_rdy_px2 (pcx_fpio_data_rdy_px2),
    .pcx_fpio_data_px2 (pcx_fpio_data_px2[123:0]),
    .arst_l (arst_l),
    .grst_l (grst_l),
    .gclk (gclk),
    .cluster_cken (cluster_cken),
    .fp_cpx_req_cq (fp_cpx_req_cq[7:0]),
    .fp_cpx_data_ca (fp_cpx_data_ca[144:0]),
    .ctu_tst_pre_grst_l (ctu_tst_pre_grst_l),
    .global_shift_enable (global_shift_enable),
    .ctu_tst_scan_disable (ctu_tst_scan_disable),
    .ctu_tst_scanmode (ctu_tst_scanmode),
    .ctu_tst_macrotest (ctu_tst_macrotest),
    .ctu_tst_short_chain (ctu_tst_short_chain),
    .si (si),
    .so (so)
);
fpu_buf fpu_buf (
    .rst_n (grst_l),
    .clk (gclk),
    .fp_cpx_req_cq (fp_cpx_req_cq[7:0]),
    .fp_cpx_data_ca (fp_cpx_data_ca[144:0]),
    .l15_fp_rdy (l15_fp_rdy),
    .fpu_arb_data_rdy (fpu_arb_data_rdy),
    .fpu_arb_data (fpu_arb_data[144:0])
);
endmodule
module fpu_arb_wrap
(
    input           clk,
    input           rst_n,
    
    input [67:0]    pcx_fpio_data_px2_67_0,
    input [79:72]   pcx_fpio_data_px2_79_72,
    input [116:112] pcx_fpio_data_px2_116_112,
    input [123:118] pcx_fpio_data_px2_123_118,
    input           l15_fp_rdy,
    
    output          fpu_arb_data_rdy,
    output [144:0]  fpu_arb_data,
    output          fpu_arb_grant
);
    wire[123:0]  pcx_fpio_data_px2 = {pcx_fpio_data_px2_123_118, 
                                                           1'bx, 
                                      pcx_fpio_data_px2_116_112, 
                                                          32'bx,
                                        pcx_fpio_data_px2_79_72,
                                                           4'bx,
                                         pcx_fpio_data_px2_67_0};
    fpu_arb fpu_arb
    (
        .arst_l (rst_n),
        .grst_l (rst_n),
        .gclk (clk),
        .cluster_cken (1'b1),
        .pcx_fpio_data_rdy_px1 (1'bx),
        .pcx_fpio_data_rdy_squashed (1'bx),
        .pcx_fpio_data_px2 (pcx_fpio_data_px2),
        .l15_fp_rdy (l15_fp_rdy),
        .fpu_arb_data_rdy (fpu_arb_data_rdy),
        .fpu_arb_data (fpu_arb_data),
        .fpu_arb_grant (fpu_arb_grant),
        .ctu_tst_pre_grst_l(1'b1),
        .global_shift_enable(1'b0),
        .ctu_tst_scan_disable(1'b1),
        .ctu_tst_scanmode(),
        .ctu_tst_macrotest(1'b0),
        .ctu_tst_short_chain(),
        .si(),
        .so()
    );
endmodule
module fpu_buf (
    input wire rst_n,
    input wire clk,
    input wire [7:0] fp_cpx_req_cq,
    input wire [144:0] fp_cpx_data_ca,
    input wire l15_fp_rdy,
    output reg fpu_arb_data_rdy,
    output reg [144:0] fpu_arb_data
);
reg fp_cpx_req;
reg fp_cpx_req_d1;
reg output_rdy;
reg output_val;
reg [144:0] output_data;
reg buffer_val_next;
reg buffer_val;
reg [144:0] buffer_next;
reg [144:0] buffer;
reg buffer_wr_en;
always @*
begin
    
    fp_cpx_req = fp_cpx_req_cq[0];
    output_rdy = !l15_fp_rdy;
    
    
    output_val = (buffer_val || fp_cpx_req_d1) && output_rdy;
    output_data = buffer_val ? buffer : fp_cpx_data_ca;
    
    
    
    buffer_val_next = (buffer_val || fp_cpx_req_d1) && !output_val;
    
    buffer_wr_en = fp_cpx_req_d1 && !output_val;
    buffer_next = buffer_wr_en ? fp_cpx_data_ca : buffer;
    
    fpu_arb_data_rdy = output_val;
    fpu_arb_data = output_data;
end
always @(posedge clk)
begin
    if (~rst_n)
    begin
        fp_cpx_req_d1 <= 1'b0;
        buffer_val <= 1'b0;
        buffer <= 145'b0;
    end
    else
    begin 
        fp_cpx_req_d1 <= fp_cpx_req;
        buffer_val <= buffer_val_next;
        buffer <= buffer_next;
    end
end
endmodule
module fpu_cnt_lead0_53b (
	din,
	lead0
);
input [52:0]	din;			
output [5:0]	lead0;			
wire		din_52_49_eq_0;
wire		din_52_51_eq_0;
wire		lead0_52_49_0;
wire		din_48_45_eq_0;
wire		din_48_47_eq_0;
wire		lead0_48_45_0;
wire		din_44_41_eq_0;
wire		din_44_43_eq_0;
wire		lead0_44_41_0;
wire		din_40_37_eq_0;
wire		din_40_39_eq_0;
wire		lead0_40_37_0;
wire		din_36_33_eq_0;
wire		din_36_35_eq_0;
wire		lead0_36_33_0;
wire		din_32_29_eq_0;
wire		din_32_31_eq_0;
wire		lead0_32_29_0;
wire		din_28_25_eq_0;
wire		din_28_27_eq_0;
wire		lead0_28_25_0;
wire		din_24_21_eq_0;
wire		din_24_23_eq_0;
wire		lead0_24_21_0;
wire		din_20_17_eq_0;
wire		din_20_19_eq_0;
wire		lead0_20_17_0;
wire		din_16_13_eq_0;
wire		din_16_15_eq_0;
wire		lead0_16_13_0;
wire		din_12_9_eq_0;
wire		din_12_11_eq_0;
wire		lead0_12_9_0;
wire		din_8_5_eq_0;
wire		din_8_7_eq_0;
wire		lead0_8_5_0;
wire		din_4_1_eq_0;
wire		din_4_3_eq_0;
wire		lead0_4_1_0;
wire		lead0_0_0;
wire		din_52_45_eq_0;
wire		lead0_52_45_1;
wire		lead0_52_45_0;
wire		din_44_37_eq_0;
wire		lead0_44_37_1;
wire		lead0_44_37_0;
wire		din_36_29_eq_0;
wire		lead0_36_29_1;
wire		lead0_36_29_0;
wire		din_28_21_eq_0;
wire		lead0_28_21_1;
wire		lead0_28_21_0;
wire		din_20_13_eq_0;
wire		lead0_20_13_1;
wire		lead0_20_13_0;
wire		din_12_5_eq_0;
wire		lead0_12_5_1;
wire		lead0_12_5_0;
wire		lead0_4_0_1;
wire		lead0_4_0_0;
wire		din_52_37_eq_0;
wire		lead0_52_37_2;
wire		lead0_52_37_1;
wire		lead0_52_37_0;
wire		din_36_21_eq_0;
wire		lead0_36_21_2;
wire		lead0_36_21_1;
wire		lead0_36_21_0;
wire		din_20_5_eq_0;
wire		lead0_20_5_2;
wire		lead0_20_5_1;
wire		lead0_20_5_0;
wire		lead0_4_0_2;
wire		din_52_21_eq_0;
wire		lead0_52_21_3;
wire		lead0_52_21_2;
wire		lead0_52_21_1;
wire		lead0_52_21_0;
wire		lead0_20_0_3;
wire		lead0_20_0_2;
wire		lead0_20_0_1;
wire		lead0_20_0_0;
wire		lead0_5;
wire		lead0_4;
wire		lead0_3;
wire		lead0_2;
wire		lead0_1;
wire		lead0_0;
wire [5:0]	lead0;
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_52_49 (
	.din			(din[52:49]),
	.din_3_0_eq_0		(din_52_49_eq_0),
	.din_3_2_eq_0		(din_52_51_eq_0),
	.lead0_4b_0		(lead0_52_49_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_48_45 (
        .din                    (din[48:45]),
        .din_3_0_eq_0           (din_48_45_eq_0),
        .din_3_2_eq_0           (din_48_47_eq_0),
        .lead0_4b_0             (lead0_48_45_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_44_41 (
        .din                    (din[44:41]),
        .din_3_0_eq_0           (din_44_41_eq_0),
        .din_3_2_eq_0           (din_44_43_eq_0),
        .lead0_4b_0             (lead0_44_41_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_40_37 (
        .din                    (din[40:37]),
        .din_3_0_eq_0           (din_40_37_eq_0),
        .din_3_2_eq_0           (din_40_39_eq_0),
        .lead0_4b_0             (lead0_40_37_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_36_33 (
        .din                    (din[36:33]),
        .din_3_0_eq_0           (din_36_33_eq_0),
        .din_3_2_eq_0           (din_36_35_eq_0),
        .lead0_4b_0             (lead0_36_33_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_32_29 (
        .din                    (din[32:29]),
        .din_3_0_eq_0           (din_32_29_eq_0),
        .din_3_2_eq_0           (din_32_31_eq_0),
        .lead0_4b_0             (lead0_32_29_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_28_25 (
        .din                    (din[28:25]),
        .din_3_0_eq_0           (din_28_25_eq_0),
        .din_3_2_eq_0           (din_28_27_eq_0),
        .lead0_4b_0             (lead0_28_25_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_24_21 (
        .din                    (din[24:21]),
        .din_3_0_eq_0           (din_24_21_eq_0),
        .din_3_2_eq_0           (din_24_23_eq_0),
        .lead0_4b_0             (lead0_24_21_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_20_17 (
        .din                    (din[20:17]),
        .din_3_0_eq_0           (din_20_17_eq_0),
        .din_3_2_eq_0           (din_20_19_eq_0),
        .lead0_4b_0             (lead0_20_17_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_16_13 (
        .din                    (din[16:13]),
        .din_3_0_eq_0           (din_16_13_eq_0),
        .din_3_2_eq_0           (din_16_15_eq_0),
        .lead0_4b_0             (lead0_16_13_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_12_9 (
        .din                    (din[12:9]),
        .din_3_0_eq_0           (din_12_9_eq_0),
        .din_3_2_eq_0           (din_12_11_eq_0),
        .lead0_4b_0             (lead0_12_9_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_8_5 (
        .din                    (din[8:5]),
        .din_3_0_eq_0           (din_8_5_eq_0),
        .din_3_2_eq_0           (din_8_7_eq_0),
        .lead0_4b_0             (lead0_8_5_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_4_1 (
        .din                    (din[4:1]),
        .din_3_0_eq_0           (din_4_1_eq_0),
        .din_3_2_eq_0           (din_4_3_eq_0),
        .lead0_4b_0             (lead0_4_1_0)
);
assign lead0_0_0= (!din[0]);
fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_52_45 (
	.din_7_4_eq_0		(din_52_49_eq_0),
	.din_7_6_eq_0		(din_52_51_eq_0),
	.lead0_4b_0_hi		(lead0_52_49_0),
	.din_3_0_eq_0		(din_48_45_eq_0),
	.din_3_2_eq_0		(din_48_47_eq_0),
	.lead0_4b_0_lo		(lead0_48_45_0),
	.din_7_0_eq_0		(din_52_45_eq_0),
	.lead0_8b_1		(lead0_52_45_1),
	.lead0_8b_0		(lead0_52_45_0)
);
fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_44_37 (
        .din_7_4_eq_0           (din_44_41_eq_0),
        .din_7_6_eq_0           (din_44_43_eq_0),
        .lead0_4b_0_hi          (lead0_44_41_0),
        .din_3_0_eq_0           (din_40_37_eq_0),
        .din_3_2_eq_0           (din_40_39_eq_0),
        .lead0_4b_0_lo          (lead0_40_37_0),
        .din_7_0_eq_0           (din_44_37_eq_0),
        .lead0_8b_1             (lead0_44_37_1),
        .lead0_8b_0             (lead0_44_37_0)
);
fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_36_29 (
        .din_7_4_eq_0           (din_36_33_eq_0),
        .din_7_6_eq_0           (din_36_35_eq_0),
        .lead0_4b_0_hi          (lead0_36_33_0),
        .din_3_0_eq_0           (din_32_29_eq_0),
        .din_3_2_eq_0           (din_32_31_eq_0),
        .lead0_4b_0_lo          (lead0_32_29_0),
        .din_7_0_eq_0           (din_36_29_eq_0),
        .lead0_8b_1             (lead0_36_29_1),
        .lead0_8b_0             (lead0_36_29_0)
);
fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_28_21 (
        .din_7_4_eq_0           (din_28_25_eq_0),
        .din_7_6_eq_0           (din_28_27_eq_0),
        .lead0_4b_0_hi          (lead0_28_25_0),
        .din_3_0_eq_0           (din_24_21_eq_0),
        .din_3_2_eq_0           (din_24_23_eq_0),
        .lead0_4b_0_lo          (lead0_24_21_0),
        .din_7_0_eq_0           (din_28_21_eq_0),
        .lead0_8b_1             (lead0_28_21_1),
        .lead0_8b_0             (lead0_28_21_0)
);
fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_20_13 (
        .din_7_4_eq_0           (din_20_17_eq_0),
        .din_7_6_eq_0           (din_20_19_eq_0),
        .lead0_4b_0_hi          (lead0_20_17_0),
        .din_3_0_eq_0           (din_16_13_eq_0),
        .din_3_2_eq_0           (din_16_15_eq_0),
        .lead0_4b_0_lo          (lead0_16_13_0),
        .din_7_0_eq_0           (din_20_13_eq_0),
        .lead0_8b_1             (lead0_20_13_1),
        .lead0_8b_0             (lead0_20_13_0)
);
fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_12_5 (
        .din_7_4_eq_0           (din_12_9_eq_0),
        .din_7_6_eq_0           (din_12_11_eq_0),
        .lead0_4b_0_hi          (lead0_12_9_0),
        .din_3_0_eq_0           (din_8_5_eq_0),
        .din_3_2_eq_0           (din_8_7_eq_0),
        .lead0_4b_0_lo          (lead0_8_5_0),
        .din_7_0_eq_0           (din_12_5_eq_0),
        .lead0_8b_1             (lead0_12_5_1),
        .lead0_8b_0             (lead0_12_5_0)
);
assign lead0_4_0_1= (!din_4_1_eq_0) && din_4_3_eq_0;
assign lead0_4_0_0= ((!din_4_1_eq_0) && lead0_4_1_0)
		|| (din_4_1_eq_0 && lead0_0_0);
fpu_cnt_lead0_lvl3 i_fpu_cnt_lead0_lvl3_52_37 (
	.din_15_8_eq_0		(din_52_45_eq_0),
	.din_15_12_eq_0		(din_52_49_eq_0),
	.lead0_8b_1_hi		(lead0_52_45_1),
	.lead0_8b_0_hi		(lead0_52_45_0),
	.din_7_0_eq_0		(din_44_37_eq_0),
	.din_7_4_eq_0		(din_44_41_eq_0),
	.lead0_8b_1_lo		(lead0_44_37_1),
	.lead0_8b_0_lo		(lead0_44_37_0),
	.din_15_0_eq_0		(din_52_37_eq_0),
	.lead0_16b_2		(lead0_52_37_2),
	.lead0_16b_1		(lead0_52_37_1),
	.lead0_16b_0		(lead0_52_37_0)
);
fpu_cnt_lead0_lvl3 i_fpu_cnt_lead0_lvl3_36_21 (
        .din_15_8_eq_0          (din_36_29_eq_0),
        .din_15_12_eq_0         (din_36_33_eq_0),           
        .lead0_8b_1_hi          (lead0_36_29_1),
        .lead0_8b_0_hi          (lead0_36_29_0),
        .din_7_0_eq_0           (din_28_21_eq_0),
        .din_7_4_eq_0           (din_28_25_eq_0),
        .lead0_8b_1_lo          (lead0_28_21_1),
        .lead0_8b_0_lo          (lead0_28_21_0),
        .din_15_0_eq_0          (din_36_21_eq_0),
        .lead0_16b_2            (lead0_36_21_2),
        .lead0_16b_1            (lead0_36_21_1),
        .lead0_16b_0            (lead0_36_21_0)
);
fpu_cnt_lead0_lvl3 i_fpu_cnt_lead0_lvl3_20_5 (
        .din_15_8_eq_0          (din_20_13_eq_0),
        .din_15_12_eq_0         (din_20_17_eq_0),           
        .lead0_8b_1_hi          (lead0_20_13_1),
        .lead0_8b_0_hi          (lead0_20_13_0),
        .din_7_0_eq_0           (din_12_5_eq_0),
        .din_7_4_eq_0           (din_12_9_eq_0),
        .lead0_8b_1_lo          (lead0_12_5_1),
        .lead0_8b_0_lo          (lead0_12_5_0),
        .din_15_0_eq_0          (din_20_5_eq_0),
        .lead0_16b_2            (lead0_20_5_2),
        .lead0_16b_1            (lead0_20_5_1),
        .lead0_16b_0            (lead0_20_5_0)
);
assign lead0_4_0_2= din_4_1_eq_0;
fpu_cnt_lead0_lvl4 i_fpu_cnt_lead0_lvl4_52_21 (
	.din_31_16_eq_0		(din_52_37_eq_0),
	.din_31_24_eq_0		(din_52_45_eq_0),
	.lead0_16b_2_hi		(lead0_52_37_2),
	.lead0_16b_1_hi		(lead0_52_37_1),
	.lead0_16b_0_hi		(lead0_52_37_0),
	.din_15_0_eq_0		(din_36_21_eq_0),
	.din_15_8_eq_0		(din_36_29_eq_0),
	.lead0_16b_2_lo		(lead0_36_21_2),
	.lead0_16b_1_lo		(lead0_36_21_1),
	.lead0_16b_0_lo		(lead0_36_21_0),
	.din_31_0_eq_0		(din_52_21_eq_0),
	.lead0_32b_3		(lead0_52_21_3),
	.lead0_32b_2		(lead0_52_21_2),
	.lead0_32b_1		(lead0_52_21_1),
	.lead0_32b_0		(lead0_52_21_0)
);
fpu_cnt_lead0_lvl4 i_fpu_cnt_lead0_lvl4_20_0 (
        .din_31_16_eq_0         (din_20_5_eq_0),
        .din_31_24_eq_0         (din_20_13_eq_0),
        .lead0_16b_2_hi         (lead0_20_5_2),
        .lead0_16b_1_hi         (lead0_20_5_1),
        .lead0_16b_0_hi         (lead0_20_5_0),
        .din_15_0_eq_0          (1'b0),     
        .din_15_8_eq_0          (1'b0),
        .lead0_16b_2_lo         (lead0_4_0_2),
        .lead0_16b_1_lo         (lead0_4_0_1),
        .lead0_16b_0_lo         (lead0_4_0_0),
        .din_31_0_eq_0          (            ),
        .lead0_32b_3            (lead0_20_0_3),
        .lead0_32b_2            (lead0_20_0_2),
        .lead0_32b_1            (lead0_20_0_1),
        .lead0_32b_0            (lead0_20_0_0)
);
assign lead0_5= din_52_21_eq_0;
assign lead0_4= ((!din_52_21_eq_0) && din_52_37_eq_0)
		|| (din_52_21_eq_0 && din_20_5_eq_0);
assign lead0_3= ((!din_52_21_eq_0) && lead0_52_21_3)
		|| (din_52_21_eq_0 && lead0_20_0_3);
assign lead0_2= ((!din_52_21_eq_0) && lead0_52_21_2)
		|| (din_52_21_eq_0 && lead0_20_0_2);
assign lead0_1= ((!din_52_21_eq_0) && lead0_52_21_1)
		|| (din_52_21_eq_0 && lead0_20_0_1);
assign lead0_0= ((!din_52_21_eq_0) && lead0_52_21_0)
		|| (din_52_21_eq_0 && lead0_20_0_0);
assign lead0[5:0]= {lead0_5, lead0_4, lead0_3, lead0_2, lead0_1, lead0_0};
endmodule
module fpu_cnt_lead0_64b (
        din,
        lead0
);
input [63:0]    din;                    
output [5:0]    lead0;                  
wire		din_63_60_eq_0;
wire		din_63_62_eq_0;
wire		lead0_63_60_0;
wire		din_59_56_eq_0;
wire		din_59_58_eq_0;
wire		lead0_59_56_0;
wire		din_55_52_eq_0;
wire		din_55_54_eq_0;
wire		lead0_55_52_0;
wire		din_51_48_eq_0;
wire		din_51_50_eq_0;
wire		lead0_51_48_0;
wire		din_47_44_eq_0;
wire		din_47_46_eq_0;
wire		lead0_47_44_0;
wire		din_43_40_eq_0;
wire		din_43_42_eq_0;
wire		lead0_43_40_0;
wire		din_39_36_eq_0;
wire		din_39_38_eq_0;
wire		lead0_39_36_0;
wire		din_35_32_eq_0;
wire		din_35_34_eq_0;
wire		lead0_35_32_0;
wire		din_31_28_eq_0;
wire		din_31_30_eq_0;
wire		lead0_31_28_0;
wire		din_27_24_eq_0;
wire		din_27_26_eq_0;
wire		lead0_27_24_0;
wire		din_23_20_eq_0;
wire		din_23_22_eq_0;
wire		lead0_23_20_0;
wire		din_19_16_eq_0;
wire		din_19_18_eq_0;
wire		lead0_19_16_0;
wire		din_15_12_eq_0;
wire		din_15_14_eq_0;
wire		lead0_15_12_0;
wire		din_11_8_eq_0;
wire		din_11_10_eq_0;
wire		lead0_11_8_0;
wire		din_7_4_eq_0;
wire		din_7_6_eq_0;
wire		lead0_7_4_0;
wire		din_3_0_eq_0;
wire		din_3_2_eq_0;
wire		lead0_3_0_0;
wire		din_63_56_eq_0;
wire		lead0_63_56_1;
wire		lead0_63_56_0;
wire		din_55_48_eq_0;
wire		lead0_55_48_1;
wire		lead0_55_48_0;
wire		din_47_40_eq_0;
wire		lead0_47_40_1;
wire		lead0_47_40_0;
wire		din_39_32_eq_0;
wire		lead0_39_32_1;
wire		lead0_39_32_0;
wire		din_31_24_eq_0;
wire		lead0_31_24_1;
wire		lead0_31_24_0;
wire		din_23_16_eq_0;
wire		lead0_23_16_1;
wire		lead0_23_16_0;
wire		din_15_8_eq_0;
wire		lead0_15_8_1;
wire		lead0_15_8_0;
wire		din_7_0_eq_0;
wire		lead0_7_0_1;
wire		lead0_7_0_0;
wire		din_63_48_eq_0;
wire		lead0_63_48_2;
wire		lead0_63_48_1;
wire		lead0_63_48_0;
wire		din_47_32_eq_0;
wire		lead0_47_32_2;
wire		lead0_47_32_1;
wire		lead0_47_32_0;
wire		din_31_16_eq_0;
wire		lead0_31_16_2;
wire		lead0_31_16_1;
wire		lead0_31_16_0;
wire		din_15_0_eq_0;
wire		lead0_15_0_2;
wire		lead0_15_0_1;
wire		lead0_15_0_0;
wire		din_63_32_eq_0;
wire		lead0_63_32_3;
wire		lead0_63_32_2;
wire		lead0_63_32_1;
wire		din_31_0_eq_0;
wire		lead0_31_0_3;
wire		lead0_31_0_2;
wire		lead0_31_0_1;
wire		lead0_31_0_0;
wire		lead0_6;
wire		lead0_5;
wire		lead0_4;
wire		lead0_3;
wire		lead0_2;
wire		lead0_1;
wire		lead0_0;
wire [5:0]	lead0;
wire        lead0_63_32_0;
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_63_60 (
	.din			(din[63:60]),
	.din_3_0_eq_0		(din_63_60_eq_0),
	.din_3_2_eq_0		(din_63_62_eq_0),
	.lead0_4b_0		(lead0_63_60_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_59_56 (
        .din                    (din[59:56]),
        .din_3_0_eq_0           (din_59_56_eq_0),
        .din_3_2_eq_0           (din_59_58_eq_0),
        .lead0_4b_0             (lead0_59_56_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_55_52 (
        .din                    (din[55:52]),
        .din_3_0_eq_0           (din_55_52_eq_0),
        .din_3_2_eq_0           (din_55_54_eq_0),
        .lead0_4b_0             (lead0_55_52_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_51_48 (
        .din                    (din[51:48]),
        .din_3_0_eq_0           (din_51_48_eq_0),
        .din_3_2_eq_0           (din_51_50_eq_0),
        .lead0_4b_0             (lead0_51_48_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_47_44 (
        .din                    (din[47:44]),
        .din_3_0_eq_0           (din_47_44_eq_0),
        .din_3_2_eq_0           (din_47_46_eq_0),
        .lead0_4b_0             (lead0_47_44_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_43_40 (
        .din                    (din[43:40]),
        .din_3_0_eq_0           (din_43_40_eq_0),
        .din_3_2_eq_0           (din_43_42_eq_0),
        .lead0_4b_0             (lead0_43_40_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_39_36 (
        .din                    (din[39:36]),
        .din_3_0_eq_0           (din_39_36_eq_0),
        .din_3_2_eq_0           (din_39_38_eq_0),
        .lead0_4b_0             (lead0_39_36_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_35_32 (
        .din                    (din[35:32]),
        .din_3_0_eq_0           (din_35_32_eq_0),
        .din_3_2_eq_0           (din_35_34_eq_0),
        .lead0_4b_0             (lead0_35_32_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_31_28 (
        .din                    (din[31:28]),
        .din_3_0_eq_0           (din_31_28_eq_0),
        .din_3_2_eq_0           (din_31_30_eq_0),
        .lead0_4b_0             (lead0_31_28_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_27_24 (
        .din                    (din[27:24]),
        .din_3_0_eq_0           (din_27_24_eq_0),
        .din_3_2_eq_0           (din_27_26_eq_0),
        .lead0_4b_0             (lead0_27_24_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_23_20 (
        .din                    (din[23:20]),
        .din_3_0_eq_0           (din_23_20_eq_0),
        .din_3_2_eq_0           (din_23_22_eq_0),
        .lead0_4b_0             (lead0_23_20_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_19_16 (
        .din                    (din[19:16]),
        .din_3_0_eq_0           (din_19_16_eq_0),
        .din_3_2_eq_0           (din_19_18_eq_0),
        .lead0_4b_0             (lead0_19_16_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_15_12 (
        .din                    (din[15:12]),
        .din_3_0_eq_0           (din_15_12_eq_0),
        .din_3_2_eq_0           (din_15_14_eq_0),
        .lead0_4b_0             (lead0_15_12_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_11_8 (
        .din                    (din[11:8]),
        .din_3_0_eq_0           (din_11_8_eq_0),
        .din_3_2_eq_0           (din_11_10_eq_0),
        .lead0_4b_0             (lead0_11_8_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_7_4 (
        .din                    (din[7:4]),
        .din_3_0_eq_0           (din_7_4_eq_0),
        .din_3_2_eq_0           (din_7_6_eq_0),
        .lead0_4b_0             (lead0_7_4_0)
);
fpu_cnt_lead0_lvl1 i_fpu_cnt_lead0_lvl1_3_0 (
        .din                    (din[3:0]),
        .din_3_0_eq_0           (din_3_0_eq_0),
        .din_3_2_eq_0           (din_3_2_eq_0),
        .lead0_4b_0             (lead0_3_0_0)
);
fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_63_56 (
	.din_7_4_eq_0		(din_63_60_eq_0),
	.din_7_6_eq_0		(din_63_62_eq_0),
	.lead0_4b_0_hi		(lead0_63_60_0),
	.din_3_0_eq_0		(din_59_56_eq_0),
	.din_3_2_eq_0		(din_59_58_eq_0),
	.lead0_4b_0_lo		(lead0_59_56_0),
	.din_7_0_eq_0		(din_63_56_eq_0),
	.lead0_8b_1		(lead0_63_56_1),
	.lead0_8b_0		(lead0_63_56_0)
);
fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_55_48 (
        .din_7_4_eq_0           (din_55_52_eq_0),
        .din_7_6_eq_0           (din_55_54_eq_0),
        .lead0_4b_0_hi          (lead0_55_52_0),
        .din_3_0_eq_0           (din_51_48_eq_0),
        .din_3_2_eq_0           (din_51_50_eq_0),
        .lead0_4b_0_lo          (lead0_51_48_0),
        .din_7_0_eq_0           (din_55_48_eq_0),
        .lead0_8b_1             (lead0_55_48_1),
        .lead0_8b_0             (lead0_55_48_0)
);
fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_47_40 (
        .din_7_4_eq_0           (din_47_44_eq_0),
        .din_7_6_eq_0           (din_47_46_eq_0),
        .lead0_4b_0_hi          (lead0_47_44_0),
        .din_3_0_eq_0           (din_43_40_eq_0),
        .din_3_2_eq_0           (din_43_42_eq_0),
        .lead0_4b_0_lo          (lead0_43_40_0),
        .din_7_0_eq_0           (din_47_40_eq_0),
        .lead0_8b_1             (lead0_47_40_1),
        .lead0_8b_0             (lead0_47_40_0)
);
fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_39_32 (
        .din_7_4_eq_0           (din_39_36_eq_0),
        .din_7_6_eq_0           (din_39_38_eq_0),
        .lead0_4b_0_hi          (lead0_39_36_0),
        .din_3_0_eq_0           (din_35_32_eq_0),
        .din_3_2_eq_0           (din_35_34_eq_0),
        .lead0_4b_0_lo          (lead0_35_32_0),
        .din_7_0_eq_0           (din_39_32_eq_0),
        .lead0_8b_1             (lead0_39_32_1),
        .lead0_8b_0             (lead0_39_32_0)
);
fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_31_24 (
        .din_7_4_eq_0           (din_31_28_eq_0),
        .din_7_6_eq_0           (din_31_30_eq_0),
        .lead0_4b_0_hi          (lead0_31_28_0),
        .din_3_0_eq_0           (din_27_24_eq_0),
        .din_3_2_eq_0           (din_27_26_eq_0),
        .lead0_4b_0_lo          (lead0_27_24_0),
        .din_7_0_eq_0           (din_31_24_eq_0),
        .lead0_8b_1             (lead0_31_24_1),
        .lead0_8b_0             (lead0_31_24_0)
);
fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_23_16 (
        .din_7_4_eq_0           (din_23_20_eq_0),
        .din_7_6_eq_0           (din_23_22_eq_0),
        .lead0_4b_0_hi          (lead0_23_20_0),
        .din_3_0_eq_0           (din_19_16_eq_0),
        .din_3_2_eq_0           (din_19_18_eq_0),
        .lead0_4b_0_lo          (lead0_19_16_0),
        .din_7_0_eq_0           (din_23_16_eq_0),
        .lead0_8b_1             (lead0_23_16_1),
        .lead0_8b_0             (lead0_23_16_0)
);
fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_15_8 (
        .din_7_4_eq_0           (din_15_12_eq_0),
        .din_7_6_eq_0           (din_15_14_eq_0),
        .lead0_4b_0_hi          (lead0_15_12_0),
        .din_3_0_eq_0           (din_11_8_eq_0),
        .din_3_2_eq_0           (din_11_10_eq_0),
        .lead0_4b_0_lo          (lead0_11_8_0),
        .din_7_0_eq_0           (din_15_8_eq_0),
        .lead0_8b_1             (lead0_15_8_1),
        .lead0_8b_0             (lead0_15_8_0)
);
fpu_cnt_lead0_lvl2 i_fpu_cnt_lead0_lvl2_7_0 (
        .din_7_4_eq_0           (din_7_4_eq_0),
        .din_7_6_eq_0           (din_7_6_eq_0),
        .lead0_4b_0_hi          (lead0_7_4_0),
        .din_3_0_eq_0           (din_3_0_eq_0),
        .din_3_2_eq_0           (din_3_2_eq_0),
        .lead0_4b_0_lo          (lead0_3_0_0),
        .din_7_0_eq_0           (din_7_0_eq_0),
        .lead0_8b_1             (lead0_7_0_1),
        .lead0_8b_0             (lead0_7_0_0)
);
fpu_cnt_lead0_lvl3 i_fpu_cnt_lead0_lvl3_63_48 (
	.din_15_8_eq_0		(din_63_56_eq_0),
	.din_15_12_eq_0		(din_63_60_eq_0),
	.lead0_8b_1_hi		(lead0_63_56_1),
	.lead0_8b_0_hi		(lead0_63_56_0),
	.din_7_0_eq_0		(din_55_48_eq_0),
	.din_7_4_eq_0		(din_55_52_eq_0),
	.lead0_8b_1_lo		(lead0_55_48_1),
	.lead0_8b_0_lo		(lead0_55_48_0),
	.din_15_0_eq_0		(din_63_48_eq_0),
	.lead0_16b_2		(lead0_63_48_2),
	.lead0_16b_1		(lead0_63_48_1),
	.lead0_16b_0		(lead0_63_48_0)
);
fpu_cnt_lead0_lvl3 i_fpu_cnt_lead0_lvl3_47_32 (
        .din_15_8_eq_0          (din_47_40_eq_0),
        .din_15_12_eq_0         (din_47_44_eq_0),
        .lead0_8b_1_hi          (lead0_47_40_1),
        .lead0_8b_0_hi          (lead0_47_40_0),
        .din_7_0_eq_0           (din_39_32_eq_0),
        .din_7_4_eq_0           (din_39_36_eq_0),
        .lead0_8b_1_lo          (lead0_39_32_1),
        .lead0_8b_0_lo          (lead0_39_32_0),
        .din_15_0_eq_0          (din_47_32_eq_0),
        .lead0_16b_2            (lead0_47_32_2),
        .lead0_16b_1            (lead0_47_32_1),
        .lead0_16b_0            (lead0_47_32_0)
);
fpu_cnt_lead0_lvl3 i_fpu_cnt_lead0_lvl3_31_16 (
        .din_15_8_eq_0          (din_31_24_eq_0),
        .din_15_12_eq_0         (din_31_28_eq_0),
        .lead0_8b_1_hi          (lead0_31_24_1),
        .lead0_8b_0_hi          (lead0_31_24_0),
        .din_7_0_eq_0           (din_23_16_eq_0),
        .din_7_4_eq_0           (din_23_20_eq_0),
        .lead0_8b_1_lo          (lead0_23_16_1),
        .lead0_8b_0_lo          (lead0_23_16_0),
        .din_15_0_eq_0          (din_31_16_eq_0),
        .lead0_16b_2            (lead0_31_16_2),
        .lead0_16b_1            (lead0_31_16_1),
        .lead0_16b_0            (lead0_31_16_0)
);
fpu_cnt_lead0_lvl3 i_fpu_cnt_lead0_lvl3_15_0 (
        .din_15_8_eq_0          (din_15_8_eq_0),
        .din_15_12_eq_0         (din_15_12_eq_0),
        .lead0_8b_1_hi          (lead0_15_8_1),
        .lead0_8b_0_hi          (lead0_15_8_0),
        .din_7_0_eq_0           (din_7_0_eq_0),
        .din_7_4_eq_0           (din_7_4_eq_0),
        .lead0_8b_1_lo          (lead0_7_0_1),
        .lead0_8b_0_lo          (lead0_7_0_0),
        .din_15_0_eq_0          (din_15_0_eq_0),
        .lead0_16b_2            (lead0_15_0_2),
        .lead0_16b_1            (lead0_15_0_1),
        .lead0_16b_0            (lead0_15_0_0)
);
fpu_cnt_lead0_lvl4 i_fpu_cnt_lead0_lvl4_63_32 (
	.din_31_16_eq_0		(din_63_48_eq_0),
	.din_31_24_eq_0		(din_63_56_eq_0),
	.lead0_16b_2_hi		(lead0_63_48_2),
	.lead0_16b_1_hi		(lead0_63_48_1),
	.lead0_16b_0_hi		(lead0_63_48_0),
	.din_15_0_eq_0		(din_47_32_eq_0),
	.din_15_8_eq_0		(din_47_40_eq_0),
	.lead0_16b_2_lo		(lead0_47_32_2),
	.lead0_16b_1_lo		(lead0_47_32_1),
	.lead0_16b_0_lo		(lead0_47_32_0),
	.din_31_0_eq_0		(din_63_32_eq_0),
	.lead0_32b_3		(lead0_63_32_3),
	.lead0_32b_2		(lead0_63_32_2),
	.lead0_32b_1		(lead0_63_32_1),
	.lead0_32b_0		(lead0_63_32_0)
);
fpu_cnt_lead0_lvl4 i_fpu_cnt_lead0_lvl4_31_0 (
        .din_31_16_eq_0         (din_31_16_eq_0),
        .din_31_24_eq_0         (din_31_24_eq_0),
        .lead0_16b_2_hi         (lead0_31_16_2),
        .lead0_16b_1_hi         (lead0_31_16_1),
        .lead0_16b_0_hi         (lead0_31_16_0),
        .din_15_0_eq_0          (din_15_0_eq_0),
        .din_15_8_eq_0          (din_15_8_eq_0),
        .lead0_16b_2_lo         (lead0_15_0_2),
        .lead0_16b_1_lo         (lead0_15_0_1),
        .lead0_16b_0_lo         (lead0_15_0_0),
        .din_31_0_eq_0          (din_31_0_eq_0),
        .lead0_32b_3            (lead0_31_0_3),
        .lead0_32b_2            (lead0_31_0_2),
        .lead0_32b_1            (lead0_31_0_1),
        .lead0_32b_0            (lead0_31_0_0)
);
assign lead0_6= din_63_32_eq_0 && din_31_0_eq_0;
assign lead0_5= (!lead0_6) && din_63_32_eq_0;
assign lead0_4= ((!din_63_32_eq_0) && din_63_48_eq_0)
		|| (din_63_32_eq_0 && din_31_16_eq_0 && (!lead0_6));
assign lead0_3= ((!din_63_32_eq_0) && lead0_63_32_3)
		|| (din_63_32_eq_0 && lead0_31_0_3 && (!lead0_6));
assign lead0_2= ((!din_63_32_eq_0) && lead0_63_32_2)
		|| (din_63_32_eq_0 && lead0_31_0_2 && (!lead0_6));
 
assign lead0_1= ((!din_63_32_eq_0) && lead0_63_32_1)
		|| (din_63_32_eq_0 && lead0_31_0_1 && (!lead0_6));
 
assign lead0_0= ((!din_63_32_eq_0) && lead0_63_32_0)
		|| (din_63_32_eq_0 && lead0_31_0_0 && (!lead0_6));
assign lead0[5:0]= {lead0_5, lead0_4, lead0_3, lead0_2, lead0_1,
		lead0_0};
endmodule
module fpu_cnt_lead0_lvl1 (
	din,
	din_3_0_eq_0,
	din_3_2_eq_0,
	lead0_4b_0
);
input [3:0]	din;			
output		din_3_0_eq_0;		
output		din_3_2_eq_0;		
output		lead0_4b_0;		
wire		din_3_0_eq_0;
wire		din_3_2_eq_0;
wire		lead0_4b_0;
assign din_3_0_eq_0= (!(|din[3:0]));
assign din_3_2_eq_0= (!(|din[3:2]));
assign lead0_4b_0= ((!din_3_2_eq_0) && (!din[3]))
		|| (din_3_2_eq_0 && (!din[1]));
endmodule
module fpu_cnt_lead0_lvl2 (
	din_7_4_eq_0,
	din_7_6_eq_0,
	lead0_4b_0_hi,
	din_3_0_eq_0,
	din_3_2_eq_0,
	lead0_4b_0_lo,
	din_7_0_eq_0,
	lead0_8b_1,
	lead0_8b_0
);
input		din_7_4_eq_0;		
input		din_7_6_eq_0;		
input		lead0_4b_0_hi;		
input		din_3_0_eq_0;		
input		din_3_2_eq_0;		
input		lead0_4b_0_lo;		
output		din_7_0_eq_0;		
output		lead0_8b_1;		
output		lead0_8b_0;		
wire		din_7_0_eq_0;
wire		lead0_8b_1;
wire		lead0_8b_0;
assign din_7_0_eq_0= din_3_0_eq_0 && din_7_4_eq_0;
assign lead0_8b_1= ((!din_7_4_eq_0) && din_7_6_eq_0)
		|| (din_7_4_eq_0 && din_3_2_eq_0);
assign lead0_8b_0= ((!din_7_4_eq_0) && lead0_4b_0_hi)
		|| (din_7_4_eq_0 && lead0_4b_0_lo);
endmodule
module fpu_cnt_lead0_lvl3 (
	din_15_8_eq_0,
	din_15_12_eq_0,
	lead0_8b_1_hi,
	lead0_8b_0_hi,
	din_7_0_eq_0,
	din_7_4_eq_0,
	lead0_8b_1_lo,
	lead0_8b_0_lo,
	din_15_0_eq_0,
	lead0_16b_2,
	lead0_16b_1,
	lead0_16b_0
);
input		din_15_8_eq_0;		
input		din_15_12_eq_0;		
input		lead0_8b_1_hi;		
input		lead0_8b_0_hi;		
input		din_7_0_eq_0;		
input		din_7_4_eq_0;		
input		lead0_8b_1_lo;		
input		lead0_8b_0_lo;		
output		din_15_0_eq_0;		
output		lead0_16b_2;		
output		lead0_16b_1;		
output		lead0_16b_0;		
wire		din_15_0_eq_0;
wire		lead0_16b_2;
wire		lead0_16b_1;
wire		lead0_16b_0;
assign din_15_0_eq_0= din_7_0_eq_0 && din_15_8_eq_0;
assign lead0_16b_2= ((!din_15_8_eq_0) && din_15_12_eq_0)
		|| (din_15_8_eq_0 && din_7_4_eq_0);
assign lead0_16b_1= ((!din_15_8_eq_0) && lead0_8b_1_hi)
		|| (din_15_8_eq_0 && lead0_8b_1_lo);
assign lead0_16b_0= ((!din_15_8_eq_0) && lead0_8b_0_hi)
		|| (din_15_8_eq_0 && lead0_8b_0_lo);
endmodule
module fpu_cnt_lead0_lvl4 (
	din_31_16_eq_0,
	din_31_24_eq_0,
	lead0_16b_2_hi,
	lead0_16b_1_hi,
	lead0_16b_0_hi,
	din_15_0_eq_0,
	din_15_8_eq_0,
	lead0_16b_2_lo,
	lead0_16b_1_lo,
	lead0_16b_0_lo,
	din_31_0_eq_0,
	lead0_32b_3,
	lead0_32b_2,
	lead0_32b_1,
	lead0_32b_0
);
input		din_31_16_eq_0;		
input		din_31_24_eq_0;		
input		lead0_16b_2_hi;		
input		lead0_16b_1_hi;		
input		lead0_16b_0_hi;		
input		din_15_0_eq_0;		
input		din_15_8_eq_0;		
input		lead0_16b_2_lo;		
input		lead0_16b_1_lo;		
input		lead0_16b_0_lo;		
output		din_31_0_eq_0;		
output		lead0_32b_3;		
output		lead0_32b_2;		
output		lead0_32b_1;		
output		lead0_32b_0;		
wire		din_31_0_eq_0;
wire		lead0_32b_3;
wire		lead0_32b_2;
wire		lead0_32b_1;
wire		lead0_32b_0;
assign din_31_0_eq_0= din_15_0_eq_0 && din_31_16_eq_0;
assign lead0_32b_3= ((!din_31_16_eq_0) && din_31_24_eq_0)
		|| (din_31_16_eq_0 && din_15_8_eq_0);
assign lead0_32b_2= ((!din_31_16_eq_0) && lead0_16b_2_hi)
		|| (din_31_16_eq_0 && lead0_16b_2_lo);
assign lead0_32b_1= ((!din_31_16_eq_0) && lead0_16b_1_hi)
		|| (din_31_16_eq_0 && lead0_16b_1_lo);
assign lead0_32b_0= ((!din_31_16_eq_0) && lead0_16b_0_hi)
		|| (din_31_16_eq_0 && lead0_16b_0_lo);
endmodule
module fpu_denorm_3b (
	din1,
	din2,
	din2_din1_nz,
	din2_din1_denorm
);
input [2:0]     din1;                   
input [2:0]     din2;                   
output		din2_din1_nz;		
output		din2_din1_denorm;	
wire [2:0]	din2_din1_zero;
wire		din2_din1_nz;
wire		din2_din1_denorm;
assign din2_din1_zero[2:0]= (~(din1 | din2));
assign din2_din1_nz= (!(&din2_din1_zero[2:0]));
assign din2_din1_denorm= din2[2]
		|| (din2_din1_zero[2] && din2[1])
		|| ((&din2_din1_zero[2:1]) && din2[0]);
endmodule
module fpu_denorm_3to1 (
	din2_din1_nz_hi,
	din2_din1_denorm_hi,
	din2_din1_nz_mid,
	din2_din1_denorm_mid,
	din2_din1_nz_lo,
	din2_din1_denorm_lo,
	din2_din1_nz,
	din2_din1_denorm
);
input		din2_din1_nz_hi;	
input		din2_din1_denorm_hi;	
input		din2_din1_nz_mid;	
input		din2_din1_denorm_mid;	
input		din2_din1_nz_lo;	
input		din2_din1_denorm_lo;	
output		din2_din1_nz;		
output		din2_din1_denorm;	
wire		din2_din1_nz;
wire		din2_din1_denorm;
assign din2_din1_nz= din2_din1_nz_hi || din2_din1_nz_mid
		|| din2_din1_nz_lo;
assign din2_din1_denorm= (din2_din1_nz_hi && din2_din1_denorm_hi)
		|| ((!din2_din1_nz_hi) && din2_din1_nz_mid
			&& din2_din1_denorm_mid)
		|| ((!din2_din1_nz_hi) && (!din2_din1_nz_mid)
			&& din2_din1_denorm_lo);
endmodule
module fpu_denorm_frac (
	din1,
	din2,
	din2_din1_denorm,
	din2_din1_denorm_inv,
	din2_din1_denorma,
	din2_din1_denorm_inva
);
input [53:0]	din1;                   
input [53:0]    din2;                   
output		din2_din1_denorm;	
output		din2_din1_denorm_inv;	
output		din2_din1_denorma;	
output		din2_din1_denorm_inva;	
wire		din2_din1_nz_53_51;
wire		din2_din1_denorm_53_51;
wire		din2_din1_nz_50_48;
wire		din2_din1_denorm_50_48;
wire		din2_din1_nz_47_45;
wire		din2_din1_denorm_47_45;
wire		din2_din1_nz_44_42;
wire		din2_din1_denorm_44_42;
wire		din2_din1_nz_41_39;
wire		din2_din1_denorm_41_39;
wire		din2_din1_nz_38_36;
wire		din2_din1_denorm_38_36;
wire		din2_din1_nz_35_33;
wire		din2_din1_denorm_35_33;
wire		din2_din1_nz_32_30;
wire		din2_din1_denorm_32_30;
wire		din2_din1_nz_29_27;
wire		din2_din1_denorm_29_27;
wire		din2_din1_nz_26_24;
wire		din2_din1_denorm_26_24;
wire		din2_din1_nz_23_21;
wire		din2_din1_denorm_23_21;
wire		din2_din1_nz_20_18;
wire		din2_din1_denorm_20_18;
wire		din2_din1_nz_17_15;
wire		din2_din1_denorm_17_15;
wire		din2_din1_nz_14_12;
wire		din2_din1_denorm_14_12;
wire		din2_din1_nz_11_9;
wire		din2_din1_denorm_11_9;
wire		din2_din1_nz_8_6;
wire		din2_din1_denorm_8_6;
wire		din2_din1_nz_5_3;
wire		din2_din1_denorm_5_3;
wire		din2_din1_nz_2_0;
wire		din2_din1_denorm_2_0;
wire		din2_din1_nz_53_45;
wire		din2_din1_denorm_53_45;
wire		din2_din1_nz_44_36;
wire		din2_din1_denorm_44_36;
wire		din2_din1_nz_35_27;
wire		din2_din1_denorm_35_27;
wire		din2_din1_nz_26_18;
wire		din2_din1_denorm_26_18;
wire		din2_din1_nz_17_9;
wire		din2_din1_denorm_17_9;
wire		din2_din1_nz_8_0;
wire		din2_din1_denorm_8_0;
wire		din2_din1_nz_53_27;
wire		din2_din1_denorm_53_27;
wire		din2_din1_nz_26_0;
wire		din2_din1_denorm_26_0;
wire		din2_din1_denorm;
wire		din2_din1_denorm_inv;
wire		din2_din1_denorma;
wire		din2_din1_denorm_inva;
fpu_denorm_3b i_fpu_denorm_53_51 (
	.din1			(din1[53:51]),
	.din2			(din2[53:51]),
	.din2_din1_nz		(din2_din1_nz_53_51),
	.din2_din1_denorm	(din2_din1_denorm_53_51)
);
fpu_denorm_3b i_fpu_denorm_50_48 (
        .din1                   (din1[50:48]),
        .din2                   (din2[50:48]),
        .din2_din1_nz           (din2_din1_nz_50_48),
        .din2_din1_denorm       (din2_din1_denorm_50_48)
);
fpu_denorm_3b i_fpu_denorm_47_45 (
        .din1                   (din1[47:45]),
        .din2                   (din2[47:45]),
        .din2_din1_nz           (din2_din1_nz_47_45),
        .din2_din1_denorm       (din2_din1_denorm_47_45)
);
fpu_denorm_3b i_fpu_denorm_44_42 (
        .din1                   (din1[44:42]),
        .din2                   (din2[44:42]),
        .din2_din1_nz           (din2_din1_nz_44_42),
        .din2_din1_denorm       (din2_din1_denorm_44_42)
);
fpu_denorm_3b i_fpu_denorm_41_39 (
        .din1                   (din1[41:39]),
        .din2                   (din2[41:39]),
        .din2_din1_nz           (din2_din1_nz_41_39),
        .din2_din1_denorm       (din2_din1_denorm_41_39)
);
fpu_denorm_3b i_fpu_denorm_38_36 (
        .din1                   (din1[38:36]),
        .din2                   (din2[38:36]),
        .din2_din1_nz           (din2_din1_nz_38_36),
        .din2_din1_denorm       (din2_din1_denorm_38_36)
);
fpu_denorm_3b i_fpu_denorm_35_33 (
        .din1                   (din1[35:33]),
        .din2                   (din2[35:33]),
        .din2_din1_nz           (din2_din1_nz_35_33),
        .din2_din1_denorm       (din2_din1_denorm_35_33)
);
fpu_denorm_3b i_fpu_denorm_32_30 (
        .din1                   (din1[32:30]),
        .din2                   (din2[32:30]),
        .din2_din1_nz           (din2_din1_nz_32_30),
        .din2_din1_denorm       (din2_din1_denorm_32_30)
);
fpu_denorm_3b i_fpu_denorm_29_27 (
        .din1                   (din1[29:27]),
        .din2                   (din2[29:27]),
        .din2_din1_nz           (din2_din1_nz_29_27),
        .din2_din1_denorm       (din2_din1_denorm_29_27)
);
fpu_denorm_3b i_fpu_denorm_26_24 (
        .din1                   (din1[26:24]),
        .din2                   (din2[26:24]),
        .din2_din1_nz           (din2_din1_nz_26_24),
        .din2_din1_denorm       (din2_din1_denorm_26_24)
);
fpu_denorm_3b i_fpu_denorm_23_21 (
        .din1                   (din1[23:21]),
        .din2                   (din2[23:21]),
        .din2_din1_nz           (din2_din1_nz_23_21),
        .din2_din1_denorm       (din2_din1_denorm_23_21)
);
fpu_denorm_3b i_fpu_denorm_20_18 (
        .din1                   (din1[20:18]),
        .din2                   (din2[20:18]),
        .din2_din1_nz           (din2_din1_nz_20_18),
        .din2_din1_denorm       (din2_din1_denorm_20_18)
);
fpu_denorm_3b i_fpu_denorm_17_15 (
        .din1                   (din1[17:15]),
        .din2                   (din2[17:15]),
        .din2_din1_nz           (din2_din1_nz_17_15),
        .din2_din1_denorm       (din2_din1_denorm_17_15)
);
fpu_denorm_3b i_fpu_denorm_14_12 (
        .din1                   (din1[14:12]),
        .din2                   (din2[14:12]),
        .din2_din1_nz           (din2_din1_nz_14_12),
        .din2_din1_denorm       (din2_din1_denorm_14_12)
);
fpu_denorm_3b i_fpu_denorm_11_9 (
        .din1                   (din1[11:9]),
        .din2                   (din2[11:9]),
        .din2_din1_nz           (din2_din1_nz_11_9),
        .din2_din1_denorm       (din2_din1_denorm_11_9)
);
fpu_denorm_3b i_fpu_denorm_8_6 (
        .din1                   (din1[8:6]),
        .din2                   (din2[8:6]),
        .din2_din1_nz           (din2_din1_nz_8_6),
        .din2_din1_denorm       (din2_din1_denorm_8_6)
);
fpu_denorm_3b i_fpu_denorm_5_3 (
        .din1                   (din1[5:3]),
        .din2                   (din2[5:3]),
        .din2_din1_nz           (din2_din1_nz_5_3),
        .din2_din1_denorm       (din2_din1_denorm_5_3)
);
fpu_denorm_3b i_fpu_denorm_2_0 (
        .din1                   (din1[2:0]),
        .din2                   (din2[2:0]),
        .din2_din1_nz           (din2_din1_nz_2_0),
        .din2_din1_denorm       (din2_din1_denorm_2_0)
);
fpu_denorm_3to1 i_fpu_denorm_53_45 (
	.din2_din1_nz_hi	(din2_din1_nz_53_51),
	.din2_din1_denorm_hi	(din2_din1_denorm_53_51),
	.din2_din1_nz_mid	(din2_din1_nz_50_48),
	.din2_din1_denorm_mid	(din2_din1_denorm_50_48),
	.din2_din1_nz_lo	(din2_din1_nz_47_45),
	.din2_din1_denorm_lo	(din2_din1_denorm_47_45),
	.din2_din1_nz		(din2_din1_nz_53_45),
	.din2_din1_denorm	(din2_din1_denorm_53_45)
);
fpu_denorm_3to1 i_fpu_denorm_44_36 (
        .din2_din1_nz_hi        (din2_din1_nz_44_42),
        .din2_din1_denorm_hi    (din2_din1_denorm_44_42),
        .din2_din1_nz_mid       (din2_din1_nz_41_39),
        .din2_din1_denorm_mid   (din2_din1_denorm_41_39),
        .din2_din1_nz_lo        (din2_din1_nz_38_36),
        .din2_din1_denorm_lo    (din2_din1_denorm_38_36),
        .din2_din1_nz           (din2_din1_nz_44_36),
        .din2_din1_denorm       (din2_din1_denorm_44_36)
);
fpu_denorm_3to1 i_fpu_denorm_35_27 (
        .din2_din1_nz_hi        (din2_din1_nz_35_33),
        .din2_din1_denorm_hi    (din2_din1_denorm_35_33),
        .din2_din1_nz_mid       (din2_din1_nz_32_30),
        .din2_din1_denorm_mid   (din2_din1_denorm_32_30),
        .din2_din1_nz_lo        (din2_din1_nz_29_27),
        .din2_din1_denorm_lo    (din2_din1_denorm_29_27),
        .din2_din1_nz           (din2_din1_nz_35_27),
        .din2_din1_denorm       (din2_din1_denorm_35_27)
);
fpu_denorm_3to1 i_fpu_denorm_26_18 (
        .din2_din1_nz_hi        (din2_din1_nz_26_24),
        .din2_din1_denorm_hi    (din2_din1_denorm_26_24),
        .din2_din1_nz_mid       (din2_din1_nz_23_21),
        .din2_din1_denorm_mid   (din2_din1_denorm_23_21),
        .din2_din1_nz_lo        (din2_din1_nz_20_18),
        .din2_din1_denorm_lo    (din2_din1_denorm_20_18),
        .din2_din1_nz           (din2_din1_nz_26_18),
        .din2_din1_denorm       (din2_din1_denorm_26_18)
);
fpu_denorm_3to1 i_fpu_denorm_17_9 (
        .din2_din1_nz_hi        (din2_din1_nz_17_15),
        .din2_din1_denorm_hi    (din2_din1_denorm_17_15),
        .din2_din1_nz_mid       (din2_din1_nz_14_12),
        .din2_din1_denorm_mid   (din2_din1_denorm_14_12),
        .din2_din1_nz_lo        (din2_din1_nz_11_9),
        .din2_din1_denorm_lo    (din2_din1_denorm_11_9),
        .din2_din1_nz           (din2_din1_nz_17_9),
        .din2_din1_denorm       (din2_din1_denorm_17_9)
);
fpu_denorm_3to1 i_fpu_denorm_8_0 (
        .din2_din1_nz_hi        (din2_din1_nz_8_6),
        .din2_din1_denorm_hi    (din2_din1_denorm_8_6),
        .din2_din1_nz_mid       (din2_din1_nz_5_3),
        .din2_din1_denorm_mid   (din2_din1_denorm_5_3),
        .din2_din1_nz_lo        (din2_din1_nz_2_0),
        .din2_din1_denorm_lo    (din2_din1_denorm_2_0),
        .din2_din1_nz           (din2_din1_nz_8_0),
        .din2_din1_denorm       (din2_din1_denorm_8_0)
);
fpu_denorm_3to1 i_fpu_denorm_53_27 (
	.din2_din1_nz_hi	(din2_din1_nz_53_45),
	.din2_din1_denorm_hi	(din2_din1_denorm_53_45),
	.din2_din1_nz_mid	(din2_din1_nz_44_36),
	.din2_din1_denorm_mid	(din2_din1_denorm_44_36),
	.din2_din1_nz_lo	(din2_din1_nz_35_27),
	.din2_din1_denorm_lo	(din2_din1_denorm_35_27),
	.din2_din1_nz		(din2_din1_nz_53_27),
	.din2_din1_denorm	(din2_din1_denorm_53_27)
);
fpu_denorm_3to1 i_fpu_denorm_26_0 (
        .din2_din1_nz_hi        (din2_din1_nz_26_18),
        .din2_din1_denorm_hi    (din2_din1_denorm_26_18),
        .din2_din1_nz_mid       (din2_din1_nz_17_9),
        .din2_din1_denorm_mid   (din2_din1_denorm_17_9),
        .din2_din1_nz_lo        (din2_din1_nz_8_0),
        .din2_din1_denorm_lo    (din2_din1_denorm_8_0),
        .din2_din1_nz           (din2_din1_nz_26_0),
        .din2_din1_denorm       (din2_din1_denorm_26_0)
);
assign din2_din1_denorm= (din2_din1_nz_53_27 && din2_din1_denorm_53_27)
		|| ((!din2_din1_nz_53_27) && (!din2_din1_nz_26_0))
		|| ((!din2_din1_nz_53_27) && din2_din1_denorm_26_0);
assign din2_din1_denorm_inv= (!din2_din1_denorm);
assign din2_din1_denorma= din2_din1_denorm;
assign din2_din1_denorm_inva= din2_din1_denorm_inv;
endmodule
module fpu_div (
	inq_op,
	inq_rnd_mode,
	inq_id,
	inq_in1,
	inq_in1_53_0_neq_0,
	inq_in1_50_0_neq_0,
	inq_in1_53_32_neq_0,
	inq_in1_exp_eq_0,
	inq_in1_exp_neq_ffs,
	inq_in2,
	inq_in2_53_0_neq_0,
	inq_in2_50_0_neq_0,
	inq_in2_53_32_neq_0,
	inq_in2_exp_eq_0,
	inq_in2_exp_neq_ffs,
	inq_div,
	div_dest_rdy,
	fdiv_clken_l,
	fdiv_clken_l_div_exp_buf1,
	arst_l,
	grst_l,
	rclk,
	
	div_pipe_active,
	d1stg_step,
	d8stg_fdiv_in,
	div_id_out_in,
	div_exc_out,
	d8stg_fdivd,
	d8stg_fdivs,
	div_sign_out,
	div_exp_outa,
	div_frac_outa,
	se,
	si,
	so
);
input [7:0]	inq_op;			
input [1:0]	inq_rnd_mode;		
input [4:0]	inq_id;			
input [63:0]	inq_in1;		
input		inq_in1_53_0_neq_0;	
input		inq_in1_50_0_neq_0;	
input		inq_in1_53_32_neq_0;	
input		inq_in1_exp_eq_0;	
input		inq_in1_exp_neq_ffs;	
input [63:0]	inq_in2;		
input		inq_in2_53_0_neq_0;	
input		inq_in2_50_0_neq_0;	
input		inq_in2_53_32_neq_0;	
input		inq_in2_exp_eq_0;	
input		inq_in2_exp_neq_ffs;	
input		inq_div;		
input		div_dest_rdy;		
input		fdiv_clken_l;           
input		fdiv_clken_l_div_exp_buf1;           
input		arst_l;			
input		grst_l;			
input		rclk;			
output		div_pipe_active;        
output		d1stg_step;		
output		d8stg_fdiv_in;		
output [9:0]	div_id_out_in;		
output [4:0]	div_exc_out;		
output		d8stg_fdivd;		
output		d8stg_fdivs;		
output		div_sign_out;		
output [10:0]	div_exp_outa;		
output [51:0]	div_frac_outa;		
input           se;                     
input           si;                     
output          so;                     
wire		d1stg_snan_sng_in1;	
wire		d1stg_snan_dbl_in1;	
wire		d1stg_snan_sng_in2;	
wire		d1stg_snan_dbl_in2;	
wire		d1stg_step;		
wire		d1stg_dblop;		
wire		d234stg_fdiv;		
wire		d3stg_fdiv;		
wire		d4stg_fdiv;		
wire		d5stg_fdiva;		
wire		d5stg_fdivb;		
wire		d5stg_fdivs;		
wire		d5stg_fdivd;		
wire		d6stg_fdiv;		
wire		d6stg_fdivs;		
wire		d6stg_fdivd;		
wire		d7stg_fdiv;		
wire		d7stg_fdivd;		
wire		d8stg_fdiv_in;		
wire		d8stg_fdivs;		
wire		d8stg_fdivd;		
wire [9:0]	div_id_out_in;		
wire		div_sign_out;		
wire [4:0]	div_exc_out;		
wire		div_norm_frac_in1_dbl_norm; 
wire		div_norm_frac_in1_dbl_dnrm; 
wire		div_norm_frac_in1_sng_norm; 
wire		div_norm_frac_in1_sng_dnrm; 
wire		div_norm_frac_in2_dbl_norm; 
wire		div_norm_frac_in2_dbl_dnrm; 
wire		div_norm_frac_in2_sng_norm; 
wire		div_norm_frac_in2_sng_dnrm; 
wire		div_norm_inf;		
wire		div_norm_qnan;		
wire		div_norm_zero;		
wire		div_frac_add_in2_load;	
wire		d6stg_frac_out_shl1;	
wire		d6stg_frac_out_nosh;	
wire		div_frac_add_in1_add;	
wire		div_frac_add_in1_load;	
wire		d7stg_rndup_inv;	
wire		d7stg_to_0;		
wire		d7stg_to_0_inv;		
wire		div_frac_out_add_in1;	
wire		div_frac_out_add;	
wire		div_frac_out_shl1_dbl;	
wire		div_frac_out_shl1_sng;	
wire		div_frac_out_of;	
wire		div_frac_out_load;	
wire		div_expadd1_in1_dbl;	
wire		div_expadd1_in1_sng;	
wire		div_expadd1_in2_exp_in2_dbl; 
wire		div_expadd1_in2_exp_in2_sng; 
wire		div_exp1_expadd1;	
wire		div_exp1_0835;		
wire		div_exp1_0118;		
wire		div_exp1_zero;		
wire		div_exp1_load;		
wire		div_expadd2_in1_exp_out; 
wire		div_expadd2_no_decr_inv; 
wire		div_expadd2_cin;	
wire		div_exp_out_expadd22_inv; 
wire		div_exp_out_expadd2;	
wire		div_exp_out_of;		
wire		div_exp_out_exp_out;	
wire		div_exp_out_load;	
wire		div_pipe_active;        
wire [12:0]	div_exp1;		
wire [12:12]	div_expadd2;		
wire [12:0]	div_exp_out;		
wire [10:0]	div_exp_outa;		
wire [5:0]	div_shl_cnt;		
wire		d6stg_frac_0;		
wire		d6stg_frac_1;		
wire		d6stg_frac_2;		
wire		d6stg_frac_29;		
wire		d6stg_frac_30;		
wire		d6stg_frac_31;		
wire		div_frac_add_in1_neq_0;	
wire		div_frac_add_52_inv;	
wire		div_frac_add_52_inva;	
wire [54:53]	div_frac_out;		
wire [51:0]	div_frac_outa;		
wire        scan_out_fpu_div_ctl;
wire        scan_out_fpu_div_exp_dp;
fpu_div_ctl fpu_div_ctl (
	.inq_in1_51			(inq_in1[51]),
	.inq_in1_54			(inq_in1[54]),
	.inq_in1_53_0_neq_0		(inq_in1_53_0_neq_0),
	.inq_in1_50_0_neq_0		(inq_in1_50_0_neq_0),
	.inq_in1_53_32_neq_0		(inq_in1_53_32_neq_0),
	.inq_in1_exp_eq_0		(inq_in1_exp_eq_0),
	.inq_in1_exp_neq_ffs		(inq_in1_exp_neq_ffs),
	.inq_in2_51			(inq_in2[51]),
	.inq_in2_54			(inq_in2[54]),
	.inq_in2_53_0_neq_0		(inq_in2_53_0_neq_0),
	.inq_in2_50_0_neq_0		(inq_in2_50_0_neq_0),
	.inq_in2_53_32_neq_0		(inq_in2_53_32_neq_0),
	.inq_in2_exp_eq_0		(inq_in2_exp_eq_0),
	.inq_in2_exp_neq_ffs		(inq_in2_exp_neq_ffs),
	.inq_op				(inq_op[7:0]),
	.div_exp1			(div_exp1[12:0]),
	.div_dest_rdy			(div_dest_rdy),
	.inq_rnd_mode			(inq_rnd_mode[1:0]),
	.inq_id				(inq_id[4:0]),
	.inq_in1_63			(inq_in1[63]),
	.inq_in2_63			(inq_in2[63]),
	.inq_div			(inq_div),
	.div_exp_out			(div_exp_out[12:0]),
	.div_frac_add_52_inva		(div_frac_add_52_inva),
	.div_frac_add_in1_neq_0		(div_frac_add_in1_neq_0),
	.div_frac_out_54		(div_frac_out[54]),
	.d6stg_frac_0			(d6stg_frac_0),
	.d6stg_frac_1			(d6stg_frac_1),
	.d6stg_frac_2			(d6stg_frac_2),
	.d6stg_frac_29			(d6stg_frac_29),
	.d6stg_frac_30			(d6stg_frac_30),
	.d6stg_frac_31			(d6stg_frac_31),
	.div_frac_out_53		(div_frac_out[53]),
	.div_expadd2_12			(div_expadd2[12]),
	.arst_l				(arst_l),
	.grst_l				(grst_l),
	.rclk			(rclk),
	.div_pipe_active		(div_pipe_active),
	.d1stg_snan_sng_in1		(d1stg_snan_sng_in1),
	.d1stg_snan_dbl_in1		(d1stg_snan_dbl_in1),
	.d1stg_snan_sng_in2		(d1stg_snan_sng_in2),
	.d1stg_snan_dbl_in2		(d1stg_snan_dbl_in2),
	.d1stg_step			(d1stg_step),
	.d1stg_dblop			(d1stg_dblop),
	.d234stg_fdiv			(d234stg_fdiv),
	.d3stg_fdiv			(d3stg_fdiv),
	.d4stg_fdiv			(d4stg_fdiv),
	.d5stg_fdiva			(d5stg_fdiva),
	.d5stg_fdivb			(d5stg_fdivb),
	.d5stg_fdivs			(d5stg_fdivs),
	.d5stg_fdivd			(d5stg_fdivd),
	.d6stg_fdiv			(d6stg_fdiv),
	.d6stg_fdivs			(d6stg_fdivs),
	.d6stg_fdivd			(d6stg_fdivd),
	.d7stg_fdiv			(d7stg_fdiv),
	.d7stg_fdivd			(d7stg_fdivd),
	.d8stg_fdiv_in			(d8stg_fdiv_in),
	.d8stg_fdivs			(d8stg_fdivs),
	.d8stg_fdivd			(d8stg_fdivd),
	.div_id_out_in			(div_id_out_in[9:0]),
	.div_sign_out			(div_sign_out),
	.div_exc_out			(div_exc_out[4:0]),
	.div_norm_frac_in1_dbl_norm	(div_norm_frac_in1_dbl_norm),
	.div_norm_frac_in1_dbl_dnrm	(div_norm_frac_in1_dbl_dnrm),
	.div_norm_frac_in1_sng_norm	(div_norm_frac_in1_sng_norm),
	.div_norm_frac_in1_sng_dnrm	(div_norm_frac_in1_sng_dnrm),
	.div_norm_frac_in2_dbl_norm	(div_norm_frac_in2_dbl_norm),
	.div_norm_frac_in2_dbl_dnrm	(div_norm_frac_in2_dbl_dnrm),
	.div_norm_frac_in2_sng_norm	(div_norm_frac_in2_sng_norm),
	.div_norm_frac_in2_sng_dnrm	(div_norm_frac_in2_sng_dnrm),
	.div_norm_inf			(div_norm_inf),
	.div_norm_qnan			(div_norm_qnan),
	.div_norm_zero			(div_norm_zero),
	.div_frac_add_in2_load		(div_frac_add_in2_load),
	.d6stg_frac_out_shl1		(d6stg_frac_out_shl1),
	.d6stg_frac_out_nosh		(d6stg_frac_out_nosh),
	.div_frac_add_in1_add		(div_frac_add_in1_add),
	.div_frac_add_in1_load		(div_frac_add_in1_load),
	.d7stg_rndup_inv		(d7stg_rndup_inv),
	.d7stg_to_0			(d7stg_to_0),
	.d7stg_to_0_inv			(d7stg_to_0_inv),
	.div_frac_out_add_in1		(div_frac_out_add_in1),
	.div_frac_out_add		(div_frac_out_add),
	.div_frac_out_shl1_dbl		(div_frac_out_shl1_dbl),
	.div_frac_out_shl1_sng		(div_frac_out_shl1_sng),
	.div_frac_out_of		(div_frac_out_of),
	.div_frac_out_load		(div_frac_out_load),
	.div_expadd1_in1_dbl		(div_expadd1_in1_dbl),
	.div_expadd1_in1_sng		(div_expadd1_in1_sng),
	.div_expadd1_in2_exp_in2_dbl	(div_expadd1_in2_exp_in2_dbl),
	.div_expadd1_in2_exp_in2_sng	(div_expadd1_in2_exp_in2_sng),
	.div_exp1_expadd1		(div_exp1_expadd1),
	.div_exp1_0835			(div_exp1_0835),
	.div_exp1_0118			(div_exp1_0118),
	.div_exp1_zero			(div_exp1_zero),
	.div_exp1_load			(div_exp1_load),
	.div_expadd2_in1_exp_out	(div_expadd2_in1_exp_out),
	.div_expadd2_no_decr_inv	(div_expadd2_no_decr_inv),
	.div_expadd2_cin		(div_expadd2_cin),
	.div_exp_out_expadd22_inv	(div_exp_out_expadd22_inv),
	.div_exp_out_expadd2		(div_exp_out_expadd2),
	.div_exp_out_of			(div_exp_out_of),
	.div_exp_out_exp_out		(div_exp_out_exp_out),
	.div_exp_out_load		(div_exp_out_load),
	.se                             (se),
        .si                             (si),
        .so                             (scan_out_fpu_div_ctl)
);
fpu_div_exp_dp fpu_div_exp_dp (
	.inq_in1			(inq_in1[62:52]),
	.inq_in2			(inq_in2[62:52]),
	.d1stg_step			(d1stg_step),
	.d234stg_fdiv			(d234stg_fdiv),
	.div_expadd1_in1_dbl		(div_expadd1_in1_dbl),
	.div_expadd1_in1_sng		(div_expadd1_in1_sng),
	.div_expadd1_in2_exp_in2_dbl	(div_expadd1_in2_exp_in2_dbl),
	.div_expadd1_in2_exp_in2_sng	(div_expadd1_in2_exp_in2_sng),
	.d3stg_fdiv			(d3stg_fdiv),
	.d4stg_fdiv			(d4stg_fdiv),
	.div_shl_cnt			(div_shl_cnt[5:0]),
	.div_exp1_expadd1		(div_exp1_expadd1),
	.div_exp1_0835			(div_exp1_0835),
	.div_exp1_0118			(div_exp1_0118),
	.div_exp1_zero			(div_exp1_zero),
	.div_exp1_load			(div_exp1_load),
	.div_expadd2_in1_exp_out	(div_expadd2_in1_exp_out),
	.d5stg_fdiva			(d5stg_fdiva),
	.d5stg_fdivd			(d5stg_fdivd),
	.d5stg_fdivs			(d5stg_fdivs),
	.d6stg_fdiv			(d6stg_fdiv),
	.d7stg_fdiv			(d7stg_fdiv),
	.div_expadd2_no_decr_inv	(div_expadd2_no_decr_inv),
	.div_expadd2_cin		(div_expadd2_cin),
	.div_exp_out_expadd2		(div_exp_out_expadd2),
	.div_exp_out_expadd22_inv	(div_exp_out_expadd22_inv),
	.div_exp_out_of			(div_exp_out_of),
	.d7stg_to_0_inv			(d7stg_to_0_inv),
	.d7stg_fdivd			(d7stg_fdivd),
	.div_exp_out_exp_out		(div_exp_out_exp_out),
	.d7stg_rndup_inv		(d7stg_rndup_inv),
	.div_frac_add_52_inv		(div_frac_add_52_inv),
	.div_exp_out_load		(div_exp_out_load),
	.fdiv_clken_l			(fdiv_clken_l_div_exp_buf1),
	.rclk			(rclk),
	.div_exp1			(div_exp1[12:0]),
	.div_expadd2_12			(div_expadd2[12]),
	.div_exp_out			(div_exp_out[12:0]),
	.div_exp_outa			(div_exp_outa[10:0]),
	.se                             (se),
        .si                             (scan_out_fpu_div_ctl),
        .so                             (scan_out_fpu_div_exp_dp)
);
fpu_div_frac_dp fpu_div_frac_dp (
	.inq_in1			(inq_in1[54:0]),
	.inq_in2			(inq_in2[54:0]),
	.d1stg_step			(d1stg_step),
	.div_norm_frac_in1_dbl_norm	(div_norm_frac_in1_dbl_norm),
	.div_norm_frac_in1_dbl_dnrm	(div_norm_frac_in1_dbl_dnrm),
	.div_norm_frac_in1_sng_norm	(div_norm_frac_in1_sng_norm),
	.div_norm_frac_in1_sng_dnrm	(div_norm_frac_in1_sng_dnrm),
	.div_norm_frac_in2_dbl_norm	(div_norm_frac_in2_dbl_norm),
	.div_norm_frac_in2_dbl_dnrm	(div_norm_frac_in2_dbl_dnrm),
	.div_norm_frac_in2_sng_norm	(div_norm_frac_in2_sng_norm),
	.div_norm_frac_in2_sng_dnrm	(div_norm_frac_in2_sng_dnrm),
	.div_norm_inf			(div_norm_inf),
	.div_norm_qnan			(div_norm_qnan),
	.d1stg_dblop			(d1stg_dblop),
	.div_norm_zero			(div_norm_zero),
	.d1stg_snan_dbl_in1		(d1stg_snan_dbl_in1),
	.d1stg_snan_sng_in1		(d1stg_snan_sng_in1),
	.d1stg_snan_dbl_in2		(d1stg_snan_dbl_in2),
	.d1stg_snan_sng_in2		(d1stg_snan_sng_in2),
	.d3stg_fdiv			(d3stg_fdiv),
	.d6stg_fdiv			(d6stg_fdiv),
	.d6stg_fdivd			(d6stg_fdivd),
	.d6stg_fdivs			(d6stg_fdivs),
	.div_frac_add_in2_load		(div_frac_add_in2_load),
	.d6stg_frac_out_shl1		(d6stg_frac_out_shl1),
	.d6stg_frac_out_nosh		(d6stg_frac_out_nosh),
	.d4stg_fdiv			(d4stg_fdiv),
	.div_frac_add_in1_add		(div_frac_add_in1_add),
	.div_frac_add_in1_load		(div_frac_add_in1_load),
	.d5stg_fdivb			(d5stg_fdivb),
	.div_frac_out_add_in1		(div_frac_out_add_in1),
	.div_frac_out_add		(div_frac_out_add),
	.div_frac_out_shl1_dbl		(div_frac_out_shl1_dbl),
	.div_frac_out_shl1_sng		(div_frac_out_shl1_sng),
	.div_frac_out_of		(div_frac_out_of),
	.d7stg_to_0			(d7stg_to_0),
	.div_frac_out_load		(div_frac_out_load),
	.fdiv_clken_l			(fdiv_clken_l),
	.rclk			(rclk),
	.div_shl_cnt			(div_shl_cnt[5:0]),
	.d6stg_frac_0			(d6stg_frac_0),
	.d6stg_frac_1			(d6stg_frac_1),
	.d6stg_frac_2			(d6stg_frac_2),
	.d6stg_frac_29			(d6stg_frac_29),
	.d6stg_frac_30			(d6stg_frac_30),
	.d6stg_frac_31			(d6stg_frac_31),
	.div_frac_add_in1_neq_0		(div_frac_add_in1_neq_0),
	.div_frac_add_52_inv		(div_frac_add_52_inv),
	.div_frac_add_52_inva		(div_frac_add_52_inva),
	.div_frac_out_54_53      	(div_frac_out[54:53]),
	.div_frac_outa			(div_frac_outa[51:0]),
	.se                             (se),
        .si                             (scan_out_fpu_div_exp_dp),
        .so                             (so)
);
endmodule
module fpu_div_ctl (
	inq_in1_51,
	inq_in1_54,
	inq_in1_53_0_neq_0,
	inq_in1_50_0_neq_0,
	inq_in1_53_32_neq_0,
	inq_in1_exp_eq_0,
	inq_in1_exp_neq_ffs,
	inq_in2_51,
	inq_in2_54,
	inq_in2_53_0_neq_0,
	inq_in2_50_0_neq_0,
	inq_in2_53_32_neq_0,
	inq_in2_exp_eq_0,
	inq_in2_exp_neq_ffs,
	inq_op,
	div_exp1,
	div_dest_rdy,
	inq_rnd_mode,
	inq_id,
	inq_in1_63,
	inq_in2_63,
	inq_div,
	div_exp_out,
	div_frac_add_52_inva,
	div_frac_add_in1_neq_0,
	div_frac_out_54,
	d6stg_frac_0,
	d6stg_frac_1,
	d6stg_frac_2,
	d6stg_frac_29,
	d6stg_frac_30,
	d6stg_frac_31,
	div_frac_out_53,
	div_expadd2_12,
	arst_l,
	grst_l,
	rclk,
	div_pipe_active,	
	d1stg_snan_sng_in1,
	d1stg_snan_dbl_in1,
	d1stg_snan_sng_in2,
	d1stg_snan_dbl_in2,
	d1stg_step,
	d1stg_dblop,
	d234stg_fdiv,
	d3stg_fdiv,
	d4stg_fdiv,
	d5stg_fdiva,
	d5stg_fdivb,
	d5stg_fdivs,
	d5stg_fdivd,
	d6stg_fdiv,
	d6stg_fdivs,
	d6stg_fdivd,
	d7stg_fdiv,
	d7stg_fdivd,
	d8stg_fdiv_in,
	d8stg_fdivs,
	d8stg_fdivd,
	div_id_out_in,
	div_sign_out,
	div_exc_out,
	div_norm_frac_in1_dbl_norm,
	div_norm_frac_in1_dbl_dnrm,
	div_norm_frac_in1_sng_norm,
	div_norm_frac_in1_sng_dnrm,
	div_norm_frac_in2_dbl_norm,
	div_norm_frac_in2_dbl_dnrm,
	div_norm_frac_in2_sng_norm,
	div_norm_frac_in2_sng_dnrm,
	div_norm_inf,
	div_norm_qnan,
	div_norm_zero,
	div_frac_add_in2_load,
	d6stg_frac_out_shl1,
	d6stg_frac_out_nosh,
	div_frac_add_in1_add,
	div_frac_add_in1_load,
	d7stg_rndup_inv,
	d7stg_to_0,
	d7stg_to_0_inv,
	div_frac_out_add_in1,
	div_frac_out_add,
	div_frac_out_shl1_dbl,
	div_frac_out_shl1_sng,
	div_frac_out_of,
	div_frac_out_load,
	div_expadd1_in1_dbl,
	div_expadd1_in1_sng,
	div_expadd1_in2_exp_in2_dbl,
	div_expadd1_in2_exp_in2_sng,
	div_exp1_expadd1,
	div_exp1_0835,
	div_exp1_0118,
	div_exp1_zero,
	div_exp1_load,
	div_expadd2_in1_exp_out,
	div_expadd2_no_decr_inv,
	div_expadd2_cin,
	div_exp_out_expadd22_inv,
	div_exp_out_expadd2,
	div_exp_out_of,
	div_exp_out_exp_out,
	div_exp_out_load,
	se,
	si,
	so
);
parameter
		FDIVS=  8'h4d,
		FDIVD=	8'h4e;
input		inq_in1_51;		
input		inq_in1_54;		
input		inq_in1_53_0_neq_0;	
input		inq_in1_50_0_neq_0;	
input		inq_in1_53_32_neq_0;	
input		inq_in1_exp_eq_0;	
input		inq_in1_exp_neq_ffs;	
input		inq_in2_51;		
input		inq_in2_54;		
input		inq_in2_53_0_neq_0;	
input		inq_in2_50_0_neq_0;	
input		inq_in2_53_32_neq_0;	
input		inq_in2_exp_eq_0;	
input		inq_in2_exp_neq_ffs;	
input [7:0]	inq_op;			
input [12:0]	div_exp1;		
input		div_dest_rdy;		
input [1:0]	inq_rnd_mode;		
input [4:0]	inq_id;			
input		inq_in1_63;		
input		inq_in2_63;		
input		inq_div;		
input [12:0]	div_exp_out;		
input		div_frac_add_52_inva;	
input		div_frac_add_in1_neq_0;	
input		div_frac_out_54;	
input		d6stg_frac_0;		
input		d6stg_frac_1;		
input		d6stg_frac_2;		
input		d6stg_frac_29;		
input		d6stg_frac_30;		
input		d6stg_frac_31;		
input		div_frac_out_53;	
input		div_expadd2_12;		
input		arst_l;			
input		grst_l;			
input		rclk;		
output		div_pipe_active;        
output		d1stg_snan_sng_in1;	
output		d1stg_snan_dbl_in1;	
output		d1stg_snan_sng_in2;	
output		d1stg_snan_dbl_in2;	
output		d1stg_step;		
output		d1stg_dblop;		
output		d234stg_fdiv;		
output		d3stg_fdiv;		
output		d4stg_fdiv;		
output		d5stg_fdiva;		
output		d5stg_fdivb;		
output		d5stg_fdivs;		
output		d5stg_fdivd;		
output		d6stg_fdiv;		
output		d6stg_fdivs;		
output		d6stg_fdivd;		
output		d7stg_fdiv;		
output		d7stg_fdivd;		
output		d8stg_fdiv_in;		
output		d8stg_fdivs;		
output		d8stg_fdivd;		
output [9:0]	div_id_out_in;		
output		div_sign_out;		
output [4:0]	div_exc_out;		
output		div_norm_frac_in1_dbl_norm; 
output		div_norm_frac_in1_dbl_dnrm; 
output		div_norm_frac_in1_sng_norm; 
output		div_norm_frac_in1_sng_dnrm; 
output		div_norm_frac_in2_dbl_norm; 
output		div_norm_frac_in2_dbl_dnrm; 
output		div_norm_frac_in2_sng_norm; 
output		div_norm_frac_in2_sng_dnrm; 
output		div_norm_inf;		
output		div_norm_qnan;		
output		div_norm_zero;		
output		div_frac_add_in2_load;	
output		d6stg_frac_out_shl1;	
output		d6stg_frac_out_nosh;	
output		div_frac_add_in1_add;	
output		div_frac_add_in1_load;	
output		d7stg_rndup_inv;	
output		d7stg_to_0;		
output		d7stg_to_0_inv;		
output		div_frac_out_add_in1;	
output		div_frac_out_add;	
output		div_frac_out_shl1_dbl;	
output		div_frac_out_shl1_sng;	
output		div_frac_out_of;	
output		div_frac_out_load;	
output		div_expadd1_in1_dbl;	
output		div_expadd1_in1_sng;	
output		div_expadd1_in2_exp_in2_dbl; 
output		div_expadd1_in2_exp_in2_sng; 
output		div_exp1_expadd1;	
output		div_exp1_0835;		
output		div_exp1_0118;		
output		div_exp1_zero;		
output		div_exp1_load;		
output		div_expadd2_in1_exp_out; 
output		div_expadd2_no_decr_inv; 
output		div_expadd2_cin;	
output		div_exp_out_expadd22_inv; 
output		div_exp_out_expadd2;	
output		div_exp_out_of;		
output		div_exp_out_exp_out;	
output		div_exp_out_load;	
input           se;                     
input           si;                     
output          so;                     
wire		reset;
wire		div_frac_in1_51;
wire		div_frac_in1_54;
wire		div_frac_in1_53_0_neq_0;
wire		div_frac_in1_50_0_neq_0;
wire		div_frac_in1_53_32_neq_0;
wire		div_exp_in1_exp_eq_0;
wire		div_exp_in1_exp_neq_ffs;
wire		div_frac_in2_51;
wire		div_frac_in2_54;
wire		div_frac_in2_53_0_neq_0;
wire		div_frac_in2_50_0_neq_0;
wire		div_frac_in2_53_32_neq_0;
wire		div_exp_in2_exp_eq_0;
wire		div_exp_in2_exp_neq_ffs;
wire		d1stg_denorm_sng_in1;
wire		d1stg_denorm_dbl_in1;
wire		d1stg_denorm_sng_in2;
wire		d1stg_denorm_dbl_in2;
wire		d2stg_denorm_sng_in2;
wire		d2stg_denorm_dbl_in2;
wire		d1stg_norm_sng_in1;
wire		d1stg_norm_dbl_in1;
wire		d1stg_norm_sng_in2;
wire		d1stg_norm_dbl_in2;
wire		d2stg_norm_sng_in2;
wire		d2stg_norm_dbl_in2;
wire		d1stg_snan_sng_in1;
wire		d1stg_snan_dbl_in1;
wire		d1stg_snan_sng_in2;
wire		d1stg_snan_dbl_in2;
wire		d1stg_qnan_sng_in1;
wire		d1stg_qnan_dbl_in1;
wire		d1stg_qnan_sng_in2;
wire		d1stg_qnan_dbl_in2;
wire		d1stg_snan_in1;
wire		d1stg_snan_in2;
wire		d1stg_qnan_in1;
wire		d1stg_qnan_in2;
wire		d1stg_nan_sng_in1;
wire		d1stg_nan_dbl_in1;
wire		d1stg_nan_sng_in2;
wire		d1stg_nan_dbl_in2;
wire		d1stg_nan_in1;
wire		d1stg_nan_in2;
wire		d1stg_nan_in;
wire		d2stg_snan_in1;
wire		d2stg_snan_in2;
wire		d2stg_qnan_in1;
wire		d2stg_qnan_in2;
wire		d2stg_nan_in2;
wire		d2stg_nan_in;
wire		d1stg_inf_sng_in1;
wire		d1stg_inf_dbl_in1;
wire		d1stg_inf_sng_in2;
wire		d1stg_inf_dbl_in2;
wire		d1stg_inf_in1;
wire		d1stg_inf_in2;
wire		d1stg_inf_in;
wire		d1stg_2inf_in;
wire		d2stg_inf_in1;
wire		d2stg_inf_in2;
wire		d2stg_2inf_in;
wire		d1stg_infnan_sng_in1;
wire		d1stg_infnan_dbl_in1;
wire		d1stg_infnan_sng_in2;
wire		d1stg_infnan_dbl_in2;
wire		d1stg_infnan_in1;
wire		d1stg_infnan_in2;
wire		d1stg_infnan_in;
wire		d2stg_infnan_in1;
wire		d2stg_infnan_in2;
wire		d2stg_infnan_in;
wire		d1stg_zero_in1;
wire		d1stg_zero_in2;
wire		d1stg_zero_in;
wire		d1stg_2zero_in;
wire		d2stg_zero_in1;
wire		d2stg_zero_in2;
wire		d2stg_zero_in;
wire		d2stg_2zero_in;
wire		d1stg_hold;
wire		d1stg_holda;
wire		d1stg_step;
wire		d1stg_stepa;
wire [7:0]	d1stg_op_in;
wire [7:0]	d1stg_op;
wire		d1stg_div_in;
wire		d1stg_div;
wire [4:0]	d1stg_sngopa;
wire		d1stg_dblop;
wire [4:0]	d1stg_dblopa;
wire		d1stg_fdiv;
wire		d1stg_fdivs;
wire		d1stg_fdivd;
wire [2:0]	d1stg_opdec;
wire		d234stg_fdiv_in;
wire [2:0]	d2stg_opdec;
wire		d234stg_fdiv;
wire		d2stg_fdiv;
wire		d2stg_fdivs;
wire		d2stg_fdivd;
wire [2:0]	d3stg_opdec;
wire		d3stg_fdiv;
wire [2:0]	d4stg_opdec;
wire		d4stg_fdiv;
wire		d4stg_fdivs;
wire		d4stg_fdivd;
wire		d5stg_step;
wire [2:0]	d5stg_opdec;
wire		d5stg_fdiva;
wire		d5stg_fdivb_in;
wire		d5stg_fdivb;
wire		d5stg_fdiv;
wire		d5stg_fdivs;
wire		d5stg_fdivd;
wire		d6stg_step;
wire [2:0]	d6stg_opdec_in;
wire [2:0]	d6stg_opdec;
wire		d6stg_fdiv;
wire		d6stg_fdivs;
wire		d6stg_fdivd;
wire [2:0]	d7stg_opdec;
wire		d7stg_fdiv;
wire		d7stg_fdivs;
wire		d7stg_fdivd;
wire		d8stg_fdiv_in;
wire [2:0]	d8stg_opdec;
wire		d8stg_fdiv;
wire		d8stg_fdivs;
wire		d8stg_fdivd;
wire		d8stg_hold;
wire		d8stg_step;
wire [1:0]	d1stg_rnd_mode;
wire [4:0]	d1stg_id;
wire		d1stg_sign1;
wire		d1stg_sign2;
wire		d1stg_sign;
wire		div_bkend_step;
wire [1:0]	div_rnd_mode;
wire [9:0]	div_id_out_in;
wire [9:0]	div_id_out;
wire		div_sign_out;
wire [5:0]	div_cnt_plus1;
wire [5:0]	div_cnt_in;
wire		div_cnt_step;
wire [5:0]	div_cnt;
wire		div_cnt_lt_step;
wire		divs_cnt_lt_23_in;
wire		divs_cnt_lt_23;
wire		divs_cnt_lt_23a;
wire		divd_cnt_lt_52_in;
wire		divd_cnt_lt_52;
wire		divd_cnt_lt_52a;
wire		div_exc_step;
wire		div_of_mask_in;
wire		div_of_mask;
wire		div_nv_out_in;
wire		div_nv_out;
wire		div_dz_out_in;
wire		div_dz_out;
wire		d7stg_in_of;
wire		div_of_out_tmp1_in;
wire		div_of_out_tmp1;
wire		div_of_out_tmp2;
wire		div_out_52_inv;
wire		div_of_out;
wire		div_uf_out_in;
wire		div_uf_out;
wire		div_nx_out_in;
wire		div_nx_out;
wire [4:0]	div_exc_out;
wire		d1stg_spc_rslt;
wire		div_norm_frac_in1_dbl_norm;
wire		div_norm_frac_in1_dbl_dnrm;
wire		div_norm_frac_in1_sng_norm;
wire		div_norm_frac_in1_sng_dnrm;
wire		div_norm_frac_in2_dbl_norm;
wire		div_norm_frac_in2_dbl_dnrm;
wire		div_norm_frac_in2_sng_norm;
wire		div_norm_frac_in2_sng_dnrm;
wire		div_norm_inf;
wire		div_norm_qnan;
wire		div_norm_zero;
wire		div_frac_add_in2_load;
wire		d6stg_frac_out_shl1;
wire		d6stg_frac_out_nosh;
wire		div_frac_add_in1_add;
wire		div_frac_add_in1_load;
wire		d7stg_lsb_in;
wire		d7stg_grd_in;
wire		d7stg_stk_in;
wire		d7stg_lsb;
wire		d7stg_grd;
wire		d7stg_stk;
wire		d7stg_rndup;
wire		d7stg_rndup_inv;
wire		d7stg_to_0;
wire		d7stg_to_0_inv;
wire		div_frac_out_add_in1;
wire		div_frac_out_add;
wire		div_frac_out_shl1_dbl;
wire		div_frac_out_shl1_sng;
wire		div_frac_out_of;
wire		div_frac_out_load;
wire		div_expadd1_in1_dbl_in;
wire		div_expadd1_in1_dbl;
wire		div_expadd1_in1_sng_in;
wire		div_expadd1_in1_sng;
wire		div_expadd1_in2_exp_in2_dbl;
wire		div_expadd1_in2_exp_in2_sng;
wire		div_exp1_expadd1;
wire		div_exp1_0835;
wire		div_exp1_0118;
wire		div_exp1_zero;
wire		d2stg_max_exp;
wire		d2stg_zero_exp;
wire		div_exp1_load;
wire		div_expadd2_in1_exp_out_in;
wire		div_expadd2_in1_exp_out;
wire		div_expadd2_no_decr_inv_in;
wire		div_expadd2_no_decr_load;
wire		div_expadd2_no_decr_inv;
wire		div_expadd2_cin;
wire		div_exp_out_zero;
wire		div_exp_out_expadd22_inv;
wire		div_exp_out_expadd2;
wire		div_exp_out_of;
wire		div_exp_out_exp_out;
wire		div_exp_out_load;
wire		div_pipe_active_in;
wire		div_pipe_active;
wire        div_ctl_rst_l;
dffrl_async #(1)  dffrl_div_ctl (
  .din  (grst_l),
  .clk  (rclk),
  .rst_l(arst_l),
  .q    (div_ctl_rst_l),
	.se (se),
	.si (),
	.so ()
  );
assign reset= (!div_ctl_rst_l);
dffe_s #(1) i_div_frac_in1_51 (
	.din	(inq_in1_51),
	.en     (d1stg_step),
        .clk    (rclk),
 
        .q      (div_frac_in1_51),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_div_frac_in1_54 (
	.din	(inq_in1_54),
	.en     (d1stg_step),
        .clk    (rclk),
 
        .q      (div_frac_in1_54),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_div_frac_in1_53_0_neq_0 (
	.din	(inq_in1_53_0_neq_0),
	.en     (d1stg_step),
        .clk    (rclk),
 
        .q      (div_frac_in1_53_0_neq_0),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_div_frac_in1_50_0_neq_0 (
	.din	(inq_in1_50_0_neq_0),
	.en	(d1stg_step),
	.clk	(rclk),
	.q	(div_frac_in1_50_0_neq_0),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_div_frac_in1_53_32_neq_0 (
	.din	(inq_in1_53_32_neq_0),
	.en	(d1stg_step),
	.clk	(rclk),
	.q	(div_frac_in1_53_32_neq_0),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_div_exp_in1_exp_eq_0 (
        .din	(inq_in1_exp_eq_0),
        .en	(d1stg_step),
        .clk	(rclk),
 
        .q	(div_exp_in1_exp_eq_0),
 
        .se	(se),
        .si	(),
        .so	()
);
dffe_s #(1) i_div_exp_in1_exp_neq_ffs (
	.din	(inq_in1_exp_neq_ffs),
	.en	(d1stg_step),
	.clk	(rclk),
	.q	(div_exp_in1_exp_neq_ffs),
   	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_div_frac_in2_51 (
	.din	(inq_in2_51),
	.en	(d1stg_step),
	.clk	(rclk),
	.q	(div_frac_in2_51),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_div_frac_in2_54 (
	.din	(inq_in2_54),
	.en	(d1stg_step),
	.clk	(rclk),
	.q	(div_frac_in2_54),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_div_frac_in2_53_0_neq_0 (
	.din	(inq_in2_53_0_neq_0),
	.en  	(d1stg_step),
	.clk	(rclk),
	.q	(div_frac_in2_53_0_neq_0),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_div_frac_in2_50_0_neq_0 (
	.din	(inq_in2_50_0_neq_0),
	.en	(d1stg_step),
	.clk	(rclk),
	.q	(div_frac_in2_50_0_neq_0),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_div_frac_in2_53_32_neq_0 (
	.din	(inq_in2_53_32_neq_0),
	.en	(d1stg_step),
	.clk	(rclk),
	.q	(div_frac_in2_53_32_neq_0),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_div_exp_in2_exp_eq_0 (
	.din	(inq_in2_exp_eq_0),
	 .en	(d1stg_step),
	.clk	(rclk),
	.q	(div_exp_in2_exp_eq_0),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_div_exp_in2_exp_neq_ffs (
        .din	(inq_in2_exp_neq_ffs),
        .en	(d1stg_step),
        .clk	(rclk),
 
        .q	(div_exp_in2_exp_neq_ffs),
 
        .se	(se),
        .si	(),
        .so	()
);
assign d1stg_denorm_sng_in1= div_exp_in1_exp_eq_0 && d1stg_sngopa[0];
assign d1stg_denorm_dbl_in1= div_exp_in1_exp_eq_0 && d1stg_dblopa[0];
assign d1stg_denorm_sng_in2= div_exp_in2_exp_eq_0 && d1stg_sngopa[0];
assign d1stg_denorm_dbl_in2= div_exp_in2_exp_eq_0 && d1stg_dblopa[0];
dff_s #(1) i_d2stg_denorm_sng_in2 (
	.din	(d1stg_denorm_sng_in2),
	.clk	(rclk),
	.q	(d2stg_denorm_sng_in2),
	.se	(se),
	.si	(),
	.so	()
);
dff_s #(1) i_d2stg_denorm_dbl_in2 (
	.din	(d1stg_denorm_dbl_in2),
	.clk	(rclk),
	.q	(d2stg_denorm_dbl_in2),
	.se	(se),
	.si	(),
	.so	()
);
assign d1stg_norm_sng_in1= (!div_exp_in1_exp_eq_0) && d1stg_sngopa[0];
assign d1stg_norm_dbl_in1= (!div_exp_in1_exp_eq_0) && d1stg_dblopa[0];
assign d1stg_norm_sng_in2= (!div_exp_in2_exp_eq_0) && d1stg_sngopa[0];
assign d1stg_norm_dbl_in2= (!div_exp_in2_exp_eq_0) && d1stg_dblopa[0];
dff_s #(1) i_d2stg_norm_sng_in2 (
	.din	(d1stg_norm_sng_in2),
	.clk	(rclk),
	.q	(d2stg_norm_sng_in2),
	.se	(se),
	.si	(),
	.so	()
);
dff_s #(1) i_d2stg_norm_dbl_in2 (
	.din	(d1stg_norm_dbl_in2),
	.clk	(rclk),
	.q	(d2stg_norm_dbl_in2),
	.se	(se),
	.si	(),
	.so	()
);
assign d1stg_snan_sng_in1= (!div_exp_in1_exp_neq_ffs) && (!div_frac_in1_54)
		&& div_frac_in1_53_32_neq_0 && d1stg_sngopa[1];
assign d1stg_snan_dbl_in1= (!div_exp_in1_exp_neq_ffs) && (!div_frac_in1_51)
		&& div_frac_in1_50_0_neq_0 && d1stg_dblopa[1];
assign d1stg_snan_sng_in2= (!div_exp_in2_exp_neq_ffs) && (!div_frac_in2_54)
                && div_frac_in2_53_32_neq_0 && d1stg_sngopa[1];
assign d1stg_snan_dbl_in2= (!div_exp_in2_exp_neq_ffs) && (!div_frac_in2_51)
                && div_frac_in2_50_0_neq_0 && d1stg_dblopa[1];
assign d1stg_qnan_sng_in1= (!div_exp_in1_exp_neq_ffs) && div_frac_in1_54
		&& d1stg_sngopa[1];
assign d1stg_qnan_dbl_in1= (!div_exp_in1_exp_neq_ffs) && div_frac_in1_51
		&& d1stg_dblopa[1];
assign d1stg_qnan_sng_in2= (!div_exp_in2_exp_neq_ffs) && div_frac_in2_54
                && d1stg_sngopa[1];
assign d1stg_qnan_dbl_in2= (!div_exp_in2_exp_neq_ffs) && div_frac_in2_51
                && d1stg_dblopa[1];
assign d1stg_snan_in1= d1stg_snan_sng_in1 || d1stg_snan_dbl_in1;
assign d1stg_snan_in2= d1stg_snan_sng_in2 || d1stg_snan_dbl_in2;
assign d1stg_qnan_in1= d1stg_qnan_sng_in1 || d1stg_qnan_dbl_in1;
 
assign d1stg_qnan_in2= d1stg_qnan_sng_in2 || d1stg_qnan_dbl_in2;
assign d1stg_nan_sng_in1= (!div_exp_in1_exp_neq_ffs)
		&& (div_frac_in1_54 || div_frac_in1_53_32_neq_0)
		&& d1stg_sngopa[2];
assign d1stg_nan_dbl_in1= (!div_exp_in1_exp_neq_ffs)
		&& (div_frac_in1_51 || div_frac_in1_50_0_neq_0)
		&& d1stg_dblopa[2];
assign d1stg_nan_sng_in2= (!div_exp_in2_exp_neq_ffs)
		&& (div_frac_in2_54 || div_frac_in2_53_32_neq_0)
		&& d1stg_sngopa[2];
assign d1stg_nan_dbl_in2= (!div_exp_in2_exp_neq_ffs)
		&& (div_frac_in2_51 || div_frac_in2_50_0_neq_0)
		&& d1stg_dblopa[2];
assign d1stg_nan_in1= d1stg_nan_sng_in1 || d1stg_nan_dbl_in1;
assign d1stg_nan_in2= d1stg_nan_sng_in2 || d1stg_nan_dbl_in2;
assign d1stg_nan_in= d1stg_nan_in1 || d1stg_nan_in2;
dff_s #(1) i_d2stg_snan_in1 (
	.din	(d1stg_snan_in1),
	.clk	(rclk),
	.q	(d2stg_snan_in1),
	.se	(se),
	.si	(),
	.so	()
);
dff_s #(1) i_d2stg_snan_in2 (
	.din	(d1stg_snan_in2),
	.clk	(rclk),
	.q	(d2stg_snan_in2),
	.se	(se),
	.si	(),
	.so	()
);
dff_s #(1) i_d2stg_qnan_in1 (
	.din	(d1stg_qnan_in1),
	.clk	(rclk),
	.q	(d2stg_qnan_in1),
	.se	(se),
	.si	(),
	.so	()
);
dff_s #(1) i_d2stg_qnan_in2 (
	.din	(d1stg_qnan_in2),
	.clk	(rclk),
	.q	(d2stg_qnan_in2),
	.se	(se),
	.si	(),
	.so	()
);
dff_s #(1) i_d2stg_nan_in2 (
	.din	(d1stg_nan_in2),
	.clk	(rclk),
	.q	(d2stg_nan_in2),
	.se	(se),
	.si	(),
	.so	()
);
dff_s #(1) i_d2stg_nan_in (
	.din	(d1stg_nan_in),
	.clk	(rclk),
	.q	(d2stg_nan_in),
	.se	(se),
	.si	(),
	.so	()
);
assign d1stg_inf_sng_in1= (!div_exp_in1_exp_neq_ffs)
		&& (!div_frac_in1_54) && (!div_frac_in1_53_32_neq_0)
		&& d1stg_sngopa[2];
assign d1stg_inf_dbl_in1= (!div_exp_in1_exp_neq_ffs)
		&& (!div_frac_in1_51) && (!div_frac_in1_50_0_neq_0)
		&& d1stg_dblopa[2];
assign d1stg_inf_sng_in2= (!div_exp_in2_exp_neq_ffs)
		&& (!div_frac_in2_54) && (!div_frac_in2_53_32_neq_0)
		&& d1stg_sngopa[2];
assign d1stg_inf_dbl_in2= (!div_exp_in2_exp_neq_ffs)
		&& (!div_frac_in2_51) && (!div_frac_in2_50_0_neq_0)
		&& d1stg_dblopa[2];
assign d1stg_inf_in1= d1stg_inf_sng_in1 || d1stg_inf_dbl_in1;
assign d1stg_inf_in2= d1stg_inf_sng_in2 || d1stg_inf_dbl_in2;
assign d1stg_inf_in= d1stg_inf_in1 || d1stg_inf_in2;
assign d1stg_2inf_in= d1stg_inf_in1 && d1stg_inf_in2;
dff_s #(1) i_d2stg_inf_in1 (
	.din	(d1stg_inf_in1),
	.clk	(rclk),
	.q	(d2stg_inf_in1),
	.se	(se),
	.si	(),
	.so	()
);
dff_s #(1) i_d2stg_inf_in2 (
	.din	(d1stg_inf_in2),
	.clk	(rclk),
	.q	(d2stg_inf_in2),
	.se	(se),
	.si	(),
	.so	()
);
dff_s #(1) i_d2stg_2inf_in (
	.din	(d1stg_2inf_in),
	.clk	(rclk),
	.q	(d2stg_2inf_in),
	.se	(se),
	.si	(),
	.so	()
);
assign d1stg_infnan_sng_in1= (!div_exp_in1_exp_neq_ffs) && d1stg_sngopa[3];
assign d1stg_infnan_dbl_in1= (!div_exp_in1_exp_neq_ffs) && d1stg_dblopa[3];
assign d1stg_infnan_sng_in2= (!div_exp_in2_exp_neq_ffs) && d1stg_sngopa[3];
assign d1stg_infnan_dbl_in2= (!div_exp_in2_exp_neq_ffs) && d1stg_dblopa[3];
assign d1stg_infnan_in1= d1stg_infnan_sng_in1 || d1stg_infnan_dbl_in1;
assign d1stg_infnan_in2= d1stg_infnan_sng_in2 || d1stg_infnan_dbl_in2;
assign d1stg_infnan_in= d1stg_infnan_in1 || d1stg_infnan_in2;
dff_s #(1) i_d2stg_infnan_in1 (
	.din	(d1stg_infnan_in1),
	.clk	(rclk),
	.q	(d2stg_infnan_in1),
	.se	(se),
	.si	(),
	.so	()
);
dff_s #(1) i_d2stg_infnan_in2 (
	.din	(d1stg_infnan_in2),
	.clk	(rclk),
	.q	(d2stg_infnan_in2),
	.se	(se),
	.si	(),
	.so	()
);
dff_s #(1) i_d2stg_infnan_in (
	.din	(d1stg_infnan_in),
	.clk	(rclk),
	.q	(d2stg_infnan_in),
	.se	(se),
	.si	(),
	.so	()
);
assign d1stg_zero_in1= div_exp_in1_exp_eq_0
		&& (!div_frac_in1_53_0_neq_0) && (!div_frac_in1_54);
assign d1stg_zero_in2= div_exp_in2_exp_eq_0
		&& (!div_frac_in2_53_0_neq_0) && (!div_frac_in2_54);
assign d1stg_zero_in= d1stg_zero_in1 || d1stg_zero_in2;
 
assign d1stg_2zero_in= d1stg_zero_in1 && d1stg_zero_in2;
dff_s #(1) i_d2stg_zero_in1 (
	.din	(d1stg_zero_in1),
	.clk	(rclk),
	.q	(d2stg_zero_in1),
	.se	(se),
	.si	(),
	.so	()
);
dff_s #(1) i_d2stg_zero_in2 (
	.din	(d1stg_zero_in2),
	.clk	(rclk),
	.q	(d2stg_zero_in2),
	.se	(se),
	.si	(),
	.so	()
);
dff_s #(1) i_d2stg_zero_in (
	.din	(d1stg_zero_in),
	.clk	(rclk),
	.q	(d2stg_zero_in),
	.se	(se),
	.si	(),
	.so	()
);
dff_s #(1) i_d2stg_2zero_in (
	.din	(d1stg_2zero_in),
	.clk	(rclk),
	.q	(d2stg_2zero_in),
	.se	(se),
	.si	(),
	.so	()
);
assign d1stg_hold= d1stg_div 
		|| d234stg_fdiv
		|| divs_cnt_lt_23
		|| divd_cnt_lt_52;
assign d1stg_holda= d1stg_div
        	|| d234stg_fdiv
        	|| divs_cnt_lt_23a
		|| divd_cnt_lt_52a;
assign d1stg_step= (!d1stg_hold);
assign d1stg_stepa= (!d1stg_holda);
assign d1stg_op_in[7:0]= ({8{d1stg_stepa}}
			    & (inq_op[7:0] & {8{inq_div}}));
dffr_s #(8) i_d1stg_op (
	.din	(d1stg_op_in[7:0]),
	.rst	(reset),
	.clk	(rclk),
	.q	(d1stg_op[7:0]),
	.se	(se),
	.si	(),
	.so	()
);
assign d1stg_div_in= inq_div && d1stg_stepa;
dffr_s #(1) i_d1stg_div (
	.din	(d1stg_div_in),
	.rst	(reset),
        .clk	(rclk),
 
        .q	(d1stg_div),
 
        .se	(se),
        .si	(),
        .so	()
);
dffe_s #(5) i_d1stg_sngopa (
        .din	({5{inq_op[0]}}),
        .en	(d1stg_stepa),
        .clk	(rclk),
 
        .q	(d1stg_sngopa[4:0]),
 
        .se	(se),
        .si	(),
        .so	()
);
dffe_s #(1) i_d1stg_dblop (
        .din    (inq_op[1]),
        .en     (d1stg_stepa),
        .clk    (rclk),
 
        .q      (d1stg_dblop),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(5) i_d1stg_dblopa (
        .din	({5{inq_op[1]}}),
        .en	(d1stg_stepa),
        .clk	(rclk),
 
        .q	(d1stg_dblopa[4:0]),
 
        .se	(se),
        .si	(),
        .so	()
);
assign d1stg_fdiv= (d1stg_op[7:0]==FDIVS) || (d1stg_op[7:0]==FDIVD);
assign d1stg_fdivs= (d1stg_op[7:0]==FDIVS);
assign d1stg_fdivd= (d1stg_op[7:0]==FDIVD);
assign d1stg_opdec[2:0]= {d1stg_fdiv,
			d1stg_fdivs,
			d1stg_fdivd};
assign d234stg_fdiv_in= d1stg_fdiv || d2stg_fdiv || d3stg_fdiv;
dffr_s #(3) i_d2stg_opdec (
	.din	(d1stg_opdec[2:0]),
	.rst	(reset),
	.clk	(rclk),
	.q	(d2stg_opdec[2:0]),
	.se     (se),
        .si     (),
        .so     ()
);
dffr_s #(1) i_d234stg_fdiv (
	.din	(d234stg_fdiv_in),
	.rst    (reset),
        .clk    (rclk),
	.q	(d234stg_fdiv),
	.se     (se),
        .si     (),
        .so     ()
);
assign d2stg_fdiv= d2stg_opdec[2];
assign d2stg_fdivs= d2stg_opdec[1];
assign d2stg_fdivd= d2stg_opdec[0];
dffr_s #(3) i_d3stg_opdec (
        .din    (d2stg_opdec[2:0]),
        .rst    (reset),
        .clk    (rclk),
        .q      (d3stg_opdec[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign d3stg_fdiv= d3stg_opdec[2];
dffr_s #(3) i_d4stg_opdec (
        .din    (d3stg_opdec[2:0]),
        .rst    (reset),
        .clk    (rclk),
 
        .q      (d4stg_opdec[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
 
assign d4stg_fdiv= d4stg_opdec[2];
assign d4stg_fdivs= d4stg_opdec[1];
assign d4stg_fdivd= d4stg_opdec[0];
 
assign d5stg_step= (!d5stg_fdiv) || d6stg_step;
dffre_s #(3) i_d5stg_opdec (
	.din	(d4stg_opdec[2:0]),
	.en	(d5stg_step),
	.rst    (reset),
        .clk    (rclk),
        .q	(d5stg_opdec[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(1) i_d5stg_fdiva (
	.din	(d4stg_fdiv),
	.en	(d5stg_step),
	.rst	(reset),
	.clk	(rclk),
	.q	(d5stg_fdiva),
	.se	(se),
	.si	(),
	.so	()
);
assign d5stg_fdivb_in= ((d5stg_step && d4stg_fdiv)
			|| ((!d5stg_step) && d5stg_fdiv))
		&& (!reset);
dff_s #(1) i_d5stg_fdivb (
	.din	(d5stg_fdivb_in),
	.clk	(rclk),
	.q	(d5stg_fdivb),
	.se	(se),
	.si	(),
	.so	()
);
assign d5stg_fdiv= d5stg_opdec[2];
assign d5stg_fdivs= d5stg_opdec[1];
assign d5stg_fdivd= d5stg_opdec[0];
assign d6stg_step= (d5stg_fdivd && (div_cnt[5:0]==6'h36))
		|| (d5stg_fdivs && (div_cnt[5:0]==6'h19))
		|| (d5stg_fdiv && ((({7'b0, div_cnt[5:0]}==div_exp1[12:0])
					&& (div_exp1[12:0]!=13'b0))
				|| (({7'b0, div_cnt[5:0]}==div_exp1[12:0])
					&& (div_exp1[12:0]==13'b0)
					&& d8stg_step)
				|| (div_exp1[12] && d8stg_step)));
assign d6stg_opdec_in[2:0]= ({3{d6stg_step}}
			    & d5stg_opdec[2:0]);
dffr_s #(3) i_d6stg_opdec (
	.din	(d6stg_opdec_in[2:0]),
	.rst    (reset),
        .clk    (rclk),
        .q      (d6stg_opdec[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign d6stg_fdiv= d6stg_opdec[2];
assign d6stg_fdivs= d6stg_opdec[1];
assign d6stg_fdivd= d6stg_opdec[0];
dffr_s #(3) i_d7stg_opdec (
        .din    (d6stg_opdec[2:0]),
	.rst    (reset),
        .clk    (rclk),
        .q      (d7stg_opdec[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign d7stg_fdiv= d7stg_opdec[2];
assign d7stg_fdivs= d7stg_opdec[1];
assign d7stg_fdivd= d7stg_opdec[0];
assign d8stg_fdiv_in= (d8stg_step && (!reset) && d7stg_fdiv)
                || ((!d8stg_step) && (!reset) && d8stg_fdiv);
dffre_s #(3) i_d8stg_opdec (
        .din    (d7stg_opdec[2:0]),
	.en	(d8stg_step),
	.rst    (reset),
        .clk    (rclk),
        .q      (d8stg_opdec[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign d8stg_fdiv= d8stg_opdec[2];
assign d8stg_fdivs= d8stg_opdec[1];
assign d8stg_fdivd= d8stg_opdec[0];
assign d8stg_hold= d8stg_fdiv && (!div_dest_rdy);
assign d8stg_step= (!d8stg_hold);
assign div_pipe_active_in =  
   d1stg_fdiv || d2stg_fdiv || d3stg_fdiv || d4stg_fdiv |
   d5stg_fdiv || d6stg_fdiv || d7stg_fdiv || d8stg_fdiv ;
dffre_s #(1) i_div_pipe_active (
	.din	(div_pipe_active_in),
	.en     (1'b1),
        .rst    (reset),
        .clk    (rclk),
        .q      (div_pipe_active),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(2) i_d1stg_rnd_mode (
	.din	(inq_rnd_mode[1:0]),
	.en	(d1stg_stepa),
	.clk	(rclk),
	.q	(d1stg_rnd_mode[1:0]),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(5) i_d1stg_id (
        .din    (inq_id[4:0]),
        .en     (d1stg_stepa),
        .clk    (rclk),
        .q      (d1stg_id[4:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_d1stg_sign1 (
	.din	(inq_in1_63),
	.en	(d1stg_stepa),
        .clk    (rclk),
        .q      (d1stg_sign1),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_d1stg_sign2 (
        .din    (inq_in2_63),
        .en     (d1stg_stepa),
        .clk    (rclk),
        .q      (d1stg_sign2),
        .se     (se),
        .si     (),
        .so     ()
);
assign d1stg_sign= ((d1stg_sign1
				&& (!d2stg_snan_in2)
				&& (!(d2stg_qnan_in2 && (!d2stg_snan_in1))))
			^ (d1stg_sign2
				&& (!(d2stg_snan_in1 && (!d2stg_snan_in2)))
				&& (!(d2stg_qnan_in1 && (!d2stg_nan_in2)))))
		&& (!(d2stg_2inf_in || d2stg_2zero_in));
 
assign div_bkend_step= (d5stg_fdiv && (div_cnt[5:0]==6'b0) && d8stg_step);
dffe_s #(2) i_div_rnd_mode (
	.din	(d1stg_rnd_mode[1:0]),
	.en	(div_bkend_step),
	.clk    (rclk),
        .q      (div_rnd_mode[1:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign div_id_out_in[9:0]= ({10{div_bkend_step}}
			    & {(d1stg_id[4:2]==3'o7),
				(d1stg_id[4:2]==3'o6),
				(d1stg_id[4:2]==3'o5),
				(d1stg_id[4:2]==3'o4),
				(d1stg_id[4:2]==3'o3),
				(d1stg_id[4:2]==3'o2),
				(d1stg_id[4:2]==3'o1),
				(d1stg_id[4:2]==3'o0),
				d1stg_id[1:0]})
		| ({10{(!div_bkend_step)}}
			    & div_id_out[9:0]);
dff_s #(10) i_div_id_out (
	.din	(div_id_out_in[9:0]),
	.clk    (rclk),
 
        .q      (div_id_out[9:0]),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_div_sign_out (
	.din	(d1stg_sign),
	.en	(div_bkend_step),
	.clk    (rclk),
 
        .q      (div_sign_out),
	.se     (se),
        .si     (),
        .so     ()
);
assign div_cnt_plus1[5:0]= (div_cnt[5:0] + 6'h01);
assign div_cnt_in[5:0]= ({6{(d5stg_fdiv && d8stg_step)}}
			    & div_cnt_plus1[5:0])
		| ({6{d4stg_fdiv}}
			    & 6'b0);
assign div_cnt_step= (d5stg_fdiv && d8stg_step)
		|| d4stg_fdiv;
dffre_s #(6) i_div_cnt (
	.din	(div_cnt_in[5:0]),
	.en	(div_cnt_step),
	.rst	(reset),
	.clk    (rclk),
 
        .q      (div_cnt[5:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign div_cnt_lt_step= (!d5stg_fdiv) || d6stg_step || d8stg_step;
assign divs_cnt_lt_23_in= d4stg_fdivs
		|| (d5stg_fdivs && (!d6stg_step) && (div_cnt_plus1[5:0]<6'h17));
dffre_s #(1) i_divs_cnt_lt_23 (
	.din	(divs_cnt_lt_23_in),
	.en	(div_cnt_lt_step),
	.rst	(reset),
	.clk	(rclk),
	.q	(divs_cnt_lt_23),
 
        .se	(se),
        .si	(),
        .so	()
);
dffre_s #(1) i_divs_cnt_lt_23a (
        .din	(divs_cnt_lt_23_in),
        .en	(div_cnt_lt_step),
        .rst	(reset),
        .clk	(rclk),
 
        .q	(divs_cnt_lt_23a),
 
        .se	(se),
        .si	(),
        .so	()
);
assign divd_cnt_lt_52_in= d4stg_fdivd
		|| (d5stg_fdivd && (!d6stg_step) && (div_cnt_plus1[5:0]<6'h34));
dffre_s #(1) i_divd_cnt_lt_52 (
	.din	(divd_cnt_lt_52_in),
	.en	(div_cnt_lt_step),
	.rst	(reset),
	.clk	(rclk),
	.q	(divd_cnt_lt_52),
 
        .se	(se),
        .si	(),
        .so	()
);
dffre_s #(1) i_divd_cnt_lt_52a (
        .din	(divd_cnt_lt_52_in),
        .en	(div_cnt_lt_step),
        .rst	(reset),
        .clk	(rclk),
 
        .q	(divd_cnt_lt_52a),
 
        .se	(se),
        .si	(),
        .so	()
);
assign div_exc_step= d5stg_fdiv && (div_cnt[5:0]==6'b0) && d8stg_step;
assign div_of_mask_in= (!(d1stg_infnan_in || d1stg_zero_in));
dffe_s #(1) i_div_of_mask (
	.din	(div_of_mask_in),
	.en	(div_exc_step),
	.clk    (rclk),
        .q      (div_of_mask),
	.se     (se),
        .si     (),
        .so     ()
);
assign div_nv_out_in= d1stg_snan_in1 || d1stg_snan_in2 || d1stg_2inf_in
		|| d1stg_2zero_in;
dffe_s #(1) i_div_nv_out (
	.din	(div_nv_out_in),
	.en	(div_exc_step),
	.clk    (rclk),
        .q      (div_nv_out),
	.se     (se),
        .si     (),
        .so     ()
);
assign div_dz_out_in= d1stg_zero_in2 && (!d1stg_zero_in1)
		&& (!d1stg_infnan_in1);
dffe_s #(1) i_div_dz_out (
        .din    (div_dz_out_in),
        .en     (div_exc_step),
        .clk    (rclk),
 
        .q      (div_dz_out),
	.se     (se),
        .si     (),
        .so     ()
);
assign d7stg_in_of= ((!div_exp_out[12])
			&& d7stg_fdivd
			&& (div_exp_out[11] || (&div_exp_out[10:0]))
			&& div_of_mask)
		|| ((!div_exp_out[12])
			&& d7stg_fdivs
			&& ((|div_exp_out[11:8]) || (&div_exp_out[7:0]))
			&& div_of_mask);
assign div_of_out_tmp1_in= ((!div_exp_out[12])
			&& d7stg_fdivd
			&& (&div_exp_out[10:1])
			&& d7stg_rndup
			&& div_of_mask)
		|| ((!div_exp_out[12])
	                && d7stg_fdivs
			&& (&div_exp_out[7:1])
	                && d7stg_rndup
	                && div_of_mask);
dffe_s #(1) i_div_of_out_tmp1 (
	.din	(div_of_out_tmp1_in),
	.en	(d7stg_fdiv),
	.clk    (rclk),
        .q      (div_of_out_tmp1),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_div_of_out_tmp2 (
	.din	(d7stg_in_of),
	.en	(d7stg_fdiv),
	.clk	(rclk),
	.q	(div_of_out_tmp2),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_div_out_52_inv (
	.din	(div_frac_add_52_inva),
	.en	(d7stg_fdiv),
        .clk	(rclk),
 
        .q	(div_out_52_inv),
	.se	(se),
	.si	(),
        .so	()
);
assign div_of_out= div_of_out_tmp2
		|| (div_of_out_tmp1 && (!div_out_52_inv));
assign div_uf_out_in= ((!(|div_exp_out[11:0]))
			&& (div_frac_add_in1_neq_0
				|| d7stg_grd
				|| d7stg_stk)
			&& div_of_mask)
		|| (div_exp_out[12]
			&& div_of_mask);
dffe_s #(1) i_div_uf_out (
        .din    (div_uf_out_in),
        .en     (d7stg_fdiv),
        .clk    (rclk),
 
        .q      (div_uf_out),
        .se     (se),
        .si     (),
        .so     ()
);
assign div_nx_out_in= d7stg_grd || d7stg_stk;
dffe_s #(1) i_div_nx_out (
        .din    (div_nx_out_in),
        .en     (d7stg_fdiv),
        .clk    (rclk),
        .q      (div_nx_out),
        .se     (se),
        .si     (),
        .so     ()
);
assign div_exc_out[4:0] =
  {div_nv_out,
   div_of_out,
   div_uf_out,
   div_dz_out,
   (div_nx_out || div_of_out)};  
 
assign d1stg_spc_rslt= (d1stg_inf_in || d1stg_zero_in) && (!d1stg_nan_in);
assign div_norm_frac_in1_dbl_norm= d1stg_fdiv && d1stg_norm_dbl_in1
		&& (!d1stg_snan_dbl_in2)
		&& ((!d1stg_qnan_dbl_in2) || d1stg_snan_dbl_in1)
		&& (!d1stg_spc_rslt);
assign div_norm_frac_in1_dbl_dnrm= d1stg_fdiv && d1stg_denorm_dbl_in1
		&& (!d1stg_snan_dbl_in2)
		&& (!d1stg_qnan_dbl_in2)
		&& (!d1stg_spc_rslt);
assign div_norm_frac_in1_sng_norm= d1stg_fdiv && d1stg_norm_sng_in1
		&& (!d1stg_snan_sng_in2)
		&& ((!d1stg_qnan_sng_in2) || d1stg_snan_sng_in1)
		&& (!d1stg_spc_rslt);
assign div_norm_frac_in1_sng_dnrm= d1stg_fdiv && d1stg_denorm_sng_in1
		&& (!d1stg_snan_sng_in2)
		&& (!d1stg_qnan_sng_in2)
		&& (!d1stg_spc_rslt);
assign div_norm_frac_in2_dbl_norm= (d2stg_fdiv && d2stg_norm_dbl_in2
			&& (!d2stg_infnan_in) && (!d2stg_zero_in))
		|| (d1stg_fdiv && d1stg_snan_dbl_in2)
		|| (d1stg_fdiv && d1stg_qnan_dbl_in2 && (!d1stg_snan_dbl_in1));
assign div_norm_frac_in2_dbl_dnrm= d2stg_fdiv && d2stg_denorm_dbl_in2
			&& (!d2stg_infnan_in) && (!d2stg_zero_in);
assign div_norm_frac_in2_sng_norm= (d2stg_fdiv && d2stg_norm_sng_in2
			&& (!d2stg_infnan_in) && (!d2stg_zero_in))
		|| (d1stg_fdiv && d1stg_snan_sng_in2)
		|| (d1stg_fdiv && d1stg_qnan_sng_in2 && (!d1stg_snan_sng_in1));
assign div_norm_frac_in2_sng_dnrm= d2stg_fdiv && d2stg_denorm_sng_in2
			&& (!d2stg_infnan_in) && (!d2stg_zero_in);
assign div_norm_inf= (d2stg_fdiv && (d2stg_infnan_in || d2stg_zero_in))
		|| (d1stg_fdiv && ((d1stg_inf_in1 && (!d1stg_infnan_in2))
				|| (d1stg_zero_in2 && (!d1stg_infnan_in1)
					&& (!d1stg_zero_in1))));
assign div_norm_qnan= d1stg_fdiv && (d1stg_2inf_in || d1stg_2zero_in);
assign div_norm_zero= d1stg_fdiv
		&& ((d1stg_inf_in2 && (!d1stg_infnan_in1))
			|| (d1stg_zero_in1 && (!d1stg_infnan_in2)
				&& (!d1stg_zero_in2)));
assign div_frac_add_in2_load= d4stg_fdiv || d6stg_fdiv;
assign d6stg_frac_out_shl1= (!div_frac_out_54) && (!div_exp_out[12])
		&& (div_exp_out[11:1]!=11'b0);
assign d6stg_frac_out_nosh= (!d6stg_frac_out_shl1);
assign div_frac_add_in1_add= d5stg_fdiv && (!div_exp1[12]) && d8stg_step;
assign div_frac_add_in1_load= d4stg_fdiv
		|| (d5stg_fdiv && (!div_exp1[12]) && d8stg_step)
		|| d6stg_fdiv;
assign d7stg_lsb_in= (d6stg_fdivd && d6stg_frac_2)
		|| ((!d6stg_fdivd) && d6stg_frac_31);
assign d7stg_grd_in= (d6stg_fdivd && d6stg_frac_1)
		|| ((!d6stg_fdivd) && d6stg_frac_30);
assign d7stg_stk_in= (d6stg_fdivd && d6stg_frac_0)
		|| ((!d6stg_fdivd) && d6stg_frac_29)
		|| div_frac_add_in1_neq_0;
dffe_s #(1) i_d7stg_lsb (
	.din	(d7stg_lsb_in),
	.en	(d6stg_fdiv),
	.clk    (rclk),
        .q      (d7stg_lsb),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_d7stg_grd (
        .din    (d7stg_grd_in),
        .en     (d6stg_fdiv),
        .clk    (rclk),
 
        .q      (d7stg_grd),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_d7stg_stk (
        .din    (d7stg_stk_in),
        .en     (d6stg_fdiv),
        .clk    (rclk),
 
        .q      (d7stg_stk),
        .se     (se),
        .si     (),
        .so     ()
);
assign d7stg_rndup= ((div_rnd_mode[1:0]==2'b10) && (!div_sign_out)
			&& (d7stg_grd || d7stg_stk))
		|| ((div_rnd_mode[1:0]==2'b11) && div_sign_out
			&& (d7stg_grd || d7stg_stk))
		|| ((div_rnd_mode[1:0]==2'b00)
			&& ((d7stg_grd && d7stg_stk)
				|| (d7stg_grd && (!d7stg_stk) && d7stg_lsb)));
assign d7stg_rndup_inv= (!d7stg_rndup);
assign d7stg_to_0= (div_rnd_mode[1:0]==2'b01)
		|| ((div_rnd_mode[1:0]==2'b10) && div_sign_out)
		|| ((div_rnd_mode[1:0]==2'b11) && (!div_sign_out));
assign d7stg_to_0_inv= (!d7stg_to_0);
assign div_frac_out_add_in1= d7stg_fdiv && (!d7stg_rndup) && (!d7stg_in_of);
assign div_frac_out_add= d7stg_fdiv && d7stg_rndup && (!d7stg_in_of);
assign div_frac_out_shl1_dbl= d5stg_fdivd && (!div_exp1[12]) && d8stg_step;
assign div_frac_out_shl1_sng= d5stg_fdivs && (!div_exp1[12]) && d8stg_step;
assign div_frac_out_of= d7stg_fdiv && d7stg_in_of;
assign div_frac_out_load= d4stg_fdiv
		|| d7stg_fdiv
		|| div_frac_out_shl1_dbl
		|| div_frac_out_shl1_sng;
assign div_expadd1_in1_dbl_in= ((d1stg_stepa && inq_op[1])
			|| ((!d1stg_stepa) && d1stg_dblopa[4]))
		&& (!((d1stg_fdiv || d2stg_fdiv || d3stg_fdiv) && (!reset)));
dff_s #(1) i_div_expadd1_in1_dbl (
	.din	(div_expadd1_in1_dbl_in),
        .clk    (rclk),
	.q	(div_expadd1_in1_dbl),
	.se     (se),
        .si     (),
        .so     ()
);
assign div_expadd1_in1_sng_in= ((d1stg_stepa && inq_op[0])
			|| ((!d1stg_stepa) && d1stg_sngopa[4]))
		&& (!((d1stg_fdiv || d2stg_fdiv || d3stg_fdiv) && (!reset)));
dff_s #(1) i_div_expadd1_in1_sng (
	.din	(div_expadd1_in1_sng_in),
	.clk	(rclk),
	.q	(div_expadd1_in1_sng),
	.se	(se),
	.si	(),
	.so	()
);
assign div_expadd1_in2_exp_in2_dbl= d2stg_fdivd;
assign div_expadd1_in2_exp_in2_sng= d2stg_fdivs;
assign div_exp1_expadd1= d1stg_fdiv
		|| (d2stg_fdiv && (!d2stg_infnan_in) && (!d2stg_zero_in))
		|| d3stg_fdiv
		|| d4stg_fdiv;
assign div_exp1_0835= d2stg_fdivd && d2stg_max_exp;
assign div_exp1_0118= d2stg_fdivs && d2stg_max_exp;
assign div_exp1_zero= d2stg_fdiv && d2stg_zero_exp;
assign d2stg_max_exp= d2stg_nan_in || d2stg_inf_in1 || d2stg_zero_in2;
assign d2stg_zero_exp= (d2stg_inf_in2 && (!d2stg_infnan_in1))
		|| (d2stg_zero_in1 && (!d2stg_infnan_in2) && (!d2stg_zero_in2));
assign div_exp1_load= d1stg_fdiv || d2stg_fdiv || d3stg_fdiv || d4stg_fdiv;
assign div_expadd2_in1_exp_out_in= d6stg_opdec_in[2] || d6stg_fdiv;
dffr_s #(1) i_div_expadd2_in1_exp_out (
	.din	(div_expadd2_in1_exp_out_in),
	.rst	(reset),
	.clk	(rclk),
	.q	(div_expadd2_in1_exp_out),
	.se	(se),
	.si	(),
	.so	()
);
assign div_expadd2_no_decr_inv_in= (!(div_frac_out_53
		|| (div_exp1[11:0]==(({12{(!d5stg_fdivs)}} & 12'h035)
					| ({12{d5stg_fdivs}} & 12'h018)))
		|| div_expadd2_12));
assign div_expadd2_no_decr_load= d5stg_fdiv && d8stg_step;
dffe_s #(1) i_div_expadd2_no_decr_inv (
	.din	(div_expadd2_no_decr_inv_in),
	.en	(div_expadd2_no_decr_load),
	.clk	(rclk),
	.q	(div_expadd2_no_decr_inv),
	.se     (se),
        .si     (),
        .so     ()
);
assign div_expadd2_cin= d5stg_fdiv || d7stg_fdiv;
assign div_exp_out_zero= d7stg_fdiv && div_exp_out[12];
assign div_exp_out_expadd22_inv= (!(d6stg_fdiv
			|| (d5stg_fdiv && (div_cnt[5:0]==6'b0) && d8stg_step)));
assign div_exp_out_expadd2= ((d7stg_fdiv && d7stg_rndup && (!d7stg_in_of))
			|| (d5stg_fdiv && (div_cnt[5:0]==6'b0) && d8stg_step)
			|| d6stg_fdiv)
		&& (!div_exp_out_zero);
assign div_exp_out_of= d7stg_fdiv && d7stg_in_of;
assign div_exp_out_exp_out= d7stg_fdiv
		&& (!d7stg_in_of)
		&& (!div_exp_out_zero);
assign div_exp_out_load= (d5stg_fdiv && (div_cnt[5:0]==6'b0) && d8stg_step)
		|| d6stg_fdiv
		|| d7stg_fdiv;
endmodule
module fpu_div_exp_dp (
	inq_in1,
	inq_in2,
	d1stg_step,
	d234stg_fdiv,
	div_expadd1_in1_dbl,
	div_expadd1_in1_sng,
	div_expadd1_in2_exp_in2_dbl,
	div_expadd1_in2_exp_in2_sng,
	d3stg_fdiv,
	d4stg_fdiv,
	div_shl_cnt,
	div_exp1_expadd1,
	div_exp1_0835,
	div_exp1_0118,
	div_exp1_zero,
	div_exp1_load,
	div_expadd2_in1_exp_out,
	d5stg_fdiva,
	d5stg_fdivd,
	d5stg_fdivs,
	d6stg_fdiv,
	d7stg_fdiv,
	div_expadd2_no_decr_inv,
	div_expadd2_cin,
	div_exp_out_expadd2,
	div_exp_out_expadd22_inv,
	div_exp_out_of,
	d7stg_to_0_inv,
	d7stg_fdivd,
	div_exp_out_exp_out,
	d7stg_rndup_inv,
	div_frac_add_52_inv,
	div_exp_out_load,
	fdiv_clken_l,
	rclk,
	
	div_exp1,
	div_expadd2_12,
	div_exp_out,
	div_exp_outa,
	se,
	si,
	so
);
input [62:52]	inq_in1;		
input [62:52]	inq_in2;		
input		d1stg_step;		
input		d234stg_fdiv;		
input		div_expadd1_in1_dbl;	
input		div_expadd1_in1_sng;	
input		div_expadd1_in2_exp_in2_dbl; 
input		div_expadd1_in2_exp_in2_sng; 
input		d3stg_fdiv;		
input		d4stg_fdiv;		
input [5:0]	div_shl_cnt;		
input		div_exp1_expadd1;	
input		div_exp1_0835;		
input		div_exp1_0118;		
input		div_exp1_zero;		
input		div_exp1_load;		
input		div_expadd2_in1_exp_out; 
input		d5stg_fdiva;		
input		d5stg_fdivd;		
input		d5stg_fdivs;		
input		d6stg_fdiv;		
input		d7stg_fdiv;		
input		div_expadd2_no_decr_inv; 
input		div_expadd2_cin;	
input		div_exp_out_expadd2;	
input		div_exp_out_expadd22_inv; 
input		div_exp_out_of;		
input		d7stg_to_0_inv;		
input		d7stg_fdivd;		
input		div_exp_out_exp_out;	
input		d7stg_rndup_inv;	
input		div_frac_add_52_inv;	
input		div_exp_out_load;	
input		fdiv_clken_l;           
input		rclk;		
output [12:0]	div_exp1;		
output        	div_expadd2_12;		
output [12:0]	div_exp_out;		
output [10:0]	div_exp_outa;		
input           se;                     
input           si;                     
output          so;                     
wire [10:0]	div_exp_in1;
wire [10:0]	div_exp_in2;
wire [12:0]	div_expadd1_in1;
wire [12:0]	div_expadd1_in2;
wire [12:0]	div_expadd1;
wire [12:0]	div_exp1_in;
wire [12:0]	div_exp1;
wire [12:0]	div_expadd2_in1;
wire [12:0]	div_expadd2_in2;
wire [12:0]     div_expadd2;
wire         	div_expadd2_12;
wire [12:0]	div_exp_out_in;
wire [12:0]	div_exp_out;
wire [10:0]	div_exp_outa;
wire se_l;
wire        clk;
assign se_l = ~se;
    clken_buf  ckbuf_div_exp_dp (
      .clk(clk),
      .rclk(rclk),
      .enb_l(fdiv_clken_l),
      .tmb_l(se_l)
      );
dffe_s #(11) i_div_exp_in1 (
        .din    (inq_in1[62:52]),
        .en     (d1stg_step),
        .clk    (clk),
 
        .q      (div_exp_in1[10:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(11) i_div_exp_in2 (
        .din    (inq_in2[62:52]),
        .en     (d1stg_step),
        .clk    (clk),
 
        .q      (div_exp_in2[10:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign div_expadd1_in1[12:0]= ({13{d234stg_fdiv}}
			    & div_exp1[12:0])
		| ({13{div_expadd1_in1_dbl}}
			    & {2'b0, div_exp_in1[10:0]})
		| ({13{div_expadd1_in1_sng}}
			    & {5'b0, div_exp_in1[10:3]});
assign div_expadd1_in2[12:0]= ({13{div_expadd1_in1_dbl}}
			    & 13'h0436)
		| ({13{div_expadd1_in1_sng}}
			    & 13'h0099)
		| ({13{div_expadd1_in2_exp_in2_dbl}}
			    & (~{2'b0, div_exp_in2[10:0]}))
		| ({13{div_expadd1_in2_exp_in2_sng}}
			    & (~{5'b0, div_exp_in2[10:3]}))
		| ({13{d3stg_fdiv}}
			    & (~{7'b0, div_shl_cnt[5:0]}))
		| ({13{d4stg_fdiv}}
			    & {7'b0, div_shl_cnt[5:0]});
assign div_expadd1[12:0]= (div_expadd1_in1[12:0]
			+ div_expadd1_in2[12:0]);
assign div_exp1_in[12:0]= ({13{div_exp1_expadd1}}
			    & div_expadd1[12:0])
		| ({13{div_exp1_0835}}
			    & 13'h0835)
		| ({13{div_exp1_0118}}
			    & 13'h0118)
		| ({13{div_exp1_zero}}
			    & 13'h0000);
dffe_s #(13) i_div_exp1 (
	.din	(div_exp1_in[12:0]),
	.en	(div_exp1_load),
	.clk    (clk),
        .q      (div_exp1[12:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign div_expadd2_in1[12:0]= ({13{div_expadd2_in1_exp_out}}
			    & div_exp_out[12:0])
		| ({13{d5stg_fdiva}}
			    & div_exp1[12:0]);
assign div_expadd2_in2[12:0]= ({13{d5stg_fdiva}}
			    & {7'h7f, d5stg_fdivs, 1'b0, d5stg_fdivd,
				d5stg_fdivs, 1'b1, d5stg_fdivs})
		| ({13{d6stg_fdiv}}
			    & {13{div_expadd2_no_decr_inv}})
		| ({13{d7stg_fdiv}}
			    & 13'h0000);
assign div_expadd2[12:0]= (div_expadd2_in1[12:0]
			+ div_expadd2_in2[12:0]
			+ {12'b0, div_expadd2_cin});
assign div_expadd2_12 = div_expadd2[12];
assign div_exp_out_in[12:0]= ({13{(div_exp_out_expadd2
				&& (!(div_frac_add_52_inv
					&& div_exp_out_expadd22_inv)))}}
			    & div_expadd2[12:0])
		| ({13{div_exp_out_of}}
			    & {2'b00, {3{d7stg_fdivd}}, 7'h7f, d7stg_to_0_inv})
		| ({13{(div_exp_out_exp_out
			&& (div_frac_add_52_inv || d7stg_rndup_inv))}}
			    & div_exp_out[12:0]);
dffe_s #(13) i_div_exp_out (
	.din	(div_exp_out_in[12:0]),
	.en	(div_exp_out_load),
	.clk    (clk),
        .q      (div_exp_out[12:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign div_exp_outa[10:0]= div_exp_out[10:0];
endmodule
module fpu_div_frac_dp (
	inq_in1,
	inq_in2,
	d1stg_step,
	div_norm_frac_in1_dbl_norm,
	div_norm_frac_in1_dbl_dnrm,
	div_norm_frac_in1_sng_norm,
	div_norm_frac_in1_sng_dnrm,
	div_norm_frac_in2_dbl_norm,
	div_norm_frac_in2_dbl_dnrm,
	div_norm_frac_in2_sng_norm,
	div_norm_frac_in2_sng_dnrm,
	div_norm_inf,
	div_norm_qnan,
	d1stg_dblop,
	div_norm_zero,
	d1stg_snan_dbl_in1,
	d1stg_snan_sng_in1,
	d1stg_snan_dbl_in2,
	d1stg_snan_sng_in2,
	d3stg_fdiv,
	d6stg_fdiv,
	d6stg_fdivd,
	d6stg_fdivs,
	div_frac_add_in2_load,
	d6stg_frac_out_shl1,
	d6stg_frac_out_nosh,
	d4stg_fdiv,
	div_frac_add_in1_add,
	div_frac_add_in1_load,
	d5stg_fdivb,
	div_frac_out_add_in1,
	div_frac_out_add,
	div_frac_out_shl1_dbl,
	div_frac_out_shl1_sng,
	div_frac_out_of,
	d7stg_to_0,
	div_frac_out_load,
	fdiv_clken_l,
	rclk,
	
	div_shl_cnt,
	d6stg_frac_0,
	d6stg_frac_1,
	d6stg_frac_2,
	d6stg_frac_29,
	d6stg_frac_30,
	d6stg_frac_31,
	div_frac_add_in1_neq_0,
	div_frac_add_52_inv,
	div_frac_add_52_inva,
	div_frac_out_54_53,
	div_frac_outa,
	se,
	si,
	so
);
input [54:0]	inq_in1;		
input [54:0]	inq_in2;		
input		d1stg_step;		
input		div_norm_frac_in1_dbl_norm; 
input		div_norm_frac_in1_dbl_dnrm; 
input		div_norm_frac_in1_sng_norm; 
input		div_norm_frac_in1_sng_dnrm; 
input		div_norm_frac_in2_dbl_norm; 
input		div_norm_frac_in2_dbl_dnrm; 
input		div_norm_frac_in2_sng_norm; 
input		div_norm_frac_in2_sng_dnrm; 
input		div_norm_inf;		
input		div_norm_qnan;		
input		d1stg_dblop;		
input		div_norm_zero;		
input		d1stg_snan_dbl_in1;	
input		d1stg_snan_sng_in1;	
input		d1stg_snan_dbl_in2;	
input		d1stg_snan_sng_in2;	
input		d3stg_fdiv;		
input		d6stg_fdiv;		
input		d6stg_fdivd;		
input		d6stg_fdivs;		
input		div_frac_add_in2_load;	
input		d6stg_frac_out_shl1;	
input		d6stg_frac_out_nosh;	
input		d4stg_fdiv;		
input		div_frac_add_in1_add;	
input		div_frac_add_in1_load;	
input		d5stg_fdivb;		
input		div_frac_out_add_in1;	
input		div_frac_out_add;	
input		div_frac_out_shl1_dbl;	
input		div_frac_out_shl1_sng;	
input		div_frac_out_of;	
input		d7stg_to_0;		
input		div_frac_out_load;	
input		fdiv_clken_l;           
input		rclk;		
output [5:0]	div_shl_cnt;		
output		d6stg_frac_0;		
output		d6stg_frac_1;		
output		d6stg_frac_2;		
output		d6stg_frac_29;		
output		d6stg_frac_30;		
output		d6stg_frac_31;		
output		div_frac_add_in1_neq_0;	
output		div_frac_add_52_inv;	
output		div_frac_add_52_inva;	
output [1:0]  	div_frac_out_54_53;	
output [51:0]	div_frac_outa;		
input           se;                     
input           si;                     
output          so;                     
wire [54:0]	div_frac_in1;
wire [54:0]	div_frac_in2;
wire [52:0]	div_norm_inv_in;
wire [52:0]	div_norm_inv;
wire [52:0]	div_norm;
wire [5:0]	div_lead0;
wire [5:0]	div_shl_cnt;
wire [5:0]	div_shl_cnta;
wire [52:0]	div_shl_data;
wire [105:53]	div_shl_tmp;
wire [52:0]	div_shl;
wire [54:0]	div_shl_save;
wire [54:0]	div_frac_add_in2_in;
wire [54:0]	div_frac_add_in2;
wire [53:0]	d6stg_frac;
wire		d6stg_frac_0;
wire		d6stg_frac_1;
wire		d6stg_frac_2;
wire		d6stg_frac_29;
wire		d6stg_frac_30;
wire		d6stg_frac_31;
wire [54:0]	div_frac_add_in1_in;
wire [54:0]	div_frac_add_in1;
wire [54:0]	div_frac_add_in1a;
wire		div_frac_add_in1_neq_0;
wire [54:0]	div_frac_add;
wire		div_frac_add_52_inv;
wire		div_frac_add_52_inva;
wire [54:0]	div_frac_out_in;
wire  [1:0]     div_frac_out_54_53;
wire [54:0]	div_frac_out;
wire [51:0]	div_frac_outa;
wire se_l;
wire        clk;
assign se_l = ~se;
    clken_buf  ckbuf_div_frac_dp (
      .clk(clk),
      .rclk(rclk),
      .enb_l(fdiv_clken_l),
      .tmb_l(se_l)
      );
dffe_s #(55) i_div_frac_in1 (
	.din	(inq_in1[54:0]),
	.en	(d1stg_step),
	.clk    (clk),
 
        .q      (div_frac_in1[54:0]),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(55) i_div_frac_in2 (
        .din    (inq_in2[54:0]),
        .en     (d1stg_step),
        .clk    (clk),
 
        .q      (div_frac_in2[54:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign div_norm_inv_in[52:0]= (~(({53{div_norm_frac_in1_dbl_norm}}
			    & {1'b1, (div_frac_in1[51] || d1stg_snan_dbl_in1),
				div_frac_in1[50:0]})
		| ({53{div_norm_frac_in1_dbl_dnrm}}
			    & {div_frac_in1[51:0], 1'b0})
		| ({53{div_norm_frac_in1_sng_norm}}
			    & {1'b1, (div_frac_in1[54] || d1stg_snan_sng_in1),
				div_frac_in1[53:32], 29'b0})
		| ({53{div_norm_frac_in1_sng_dnrm}}
			    & {div_frac_in1[54:32], 30'b0})
		| ({53{div_norm_frac_in2_dbl_norm}}
			    & {1'b1, (div_frac_in2[51] || d1stg_snan_dbl_in2),
				div_frac_in2[50:0]})
		| ({53{div_norm_frac_in2_dbl_dnrm}}
			    & {div_frac_in2[51:0], 1'b0})
		| ({53{div_norm_frac_in2_sng_norm}}
			    & {1'b1, (div_frac_in2[54] || d1stg_snan_sng_in2),
				div_frac_in2[53:32], 29'b0})
		| ({53{div_norm_frac_in2_sng_dnrm}}
			    & {div_frac_in2[54:32], 30'b0})
		| ({53{div_norm_inf}}
			    & 53'h10000000000000)
		| ({53{div_norm_qnan}}
			    & {24'hffffff, {29{d1stg_dblop}}})
		| ({53{div_norm_zero}}
			    & 53'h00000000000000)));
dff_s #(53) i_div_norm_inv (
	.din	(div_norm_inv_in[52:0]),
	.clk	(clk),
	.q	(div_norm_inv[52:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign div_norm[52:0]= (~div_norm_inv);
fpu_cnt_lead0_53b i_div_lead0 (
	.din	(div_norm[52:0]),
	.lead0 (div_lead0[5:0])
);
dff_s #(12) i_dstg_xtra_regs (
        .din    ({div_lead0[5:0], div_lead0[5:0]}),
        .clk    (clk),
        .q      ({div_shl_cnta[5:0], div_shl_cnt[5:0]}),
        .se     (se),
        .si     (),
        .so     ()
);
dff_s #(53) i_div_shl_data (
	.din	(div_norm[52:0]),
	.clk    (clk),
        .q      (div_shl_data[52:0]),
	.se     (se),
        .si     (),
        .so     ()
);
  assign div_shl_tmp[105:53]= div_shl_data[52:0]         << div_shl_cnta[5:0];
assign div_shl[52:0]= div_shl_tmp[105:53];
dffe_s #(55) i_div_shl_save (
	.din	({2'b0, div_shl[52:0]}),
	.en	(d3stg_fdiv),
        .clk    (clk),
 
        .q      (div_shl_save[54:0]),
 
        .se     (se),
        .si     (),
        .so     ()
);
assign div_frac_add_in2_in[54:0]= ({55{d4stg_fdiv}}
			    & (~{2'b0, div_shl[52:0]}))
		| ({55{d6stg_fdiv}}
			    & {25'b0, d6stg_fdivs, 28'b0, d6stg_fdivd});
dffe_s #(55) i_div_frac_add_in2 (
	.din	(div_frac_add_in2_in[54:0]),
	.en	(div_frac_add_in2_load),
	.clk    (clk),
        .q      (div_frac_add_in2[54:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign d6stg_frac[53:0]= ({54{d6stg_frac_out_shl1}}
			    & {div_frac_out[52:0], 1'b0})
		| ({54{d6stg_frac_out_nosh}}
			    & div_frac_out[53:0]);
assign d6stg_frac_0= d6stg_frac[0];
assign d6stg_frac_1= d6stg_frac[1];
assign d6stg_frac_2= d6stg_frac[2];
assign d6stg_frac_29= d6stg_frac[29];
assign d6stg_frac_30= d6stg_frac[30];
assign d6stg_frac_31= d6stg_frac[31];
assign div_frac_add_in1_in[54:0]= ({55{d4stg_fdiv}}
			    & div_shl_save[54:0])
		| ({55{(div_frac_add_in1_add && (!div_frac_add[54]))}}
			    & {div_frac_add[53:0], 1'b0})
		| ({55{(div_frac_add_in1_add && div_frac_add[54])}}
			    & {div_frac_add_in1[53:0], 1'b0})
		| ({55{d6stg_fdiv}}
			    & {3'b0, d6stg_frac[53:31],
				(d6stg_frac[30:2] & {29{d6stg_fdivd}})});
dffe_s #(55) i_div_frac_add_in1 (
	.din	(div_frac_add_in1_in[54:0]),
	.en	(div_frac_add_in1_load),
	.clk    (clk),
        .q      (div_frac_add_in1[54:0]),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(55) i_div_frac_add_in1a (
	.din	(div_frac_add_in1_in[54:0]),
	.en	(div_frac_add_in1_load),
	.clk	(clk),
	.q	(div_frac_add_in1a[54:0]),
	.se	(se),
	.si	(),
	.so	()
);
assign div_frac_add_in1_neq_0= (|div_frac_add_in1[54:0]);
assign div_frac_add[54:0]= (div_frac_add_in1a[54:0]
			+ div_frac_add_in2[54:0]
			+ {54'b0, d5stg_fdivb});
assign div_frac_add_52_inv= (!div_frac_add[52]);
assign div_frac_add_52_inva= (!div_frac_add[52]);
assign div_frac_out_in[54:0]= ({55{d4stg_fdiv}}
			    & 55'b0)
		| ({55{div_frac_out_add_in1}}
			    & div_frac_add_in1[54:0])
		| ({55{div_frac_out_add}}
			    & div_frac_add[54:0])
		| ({55{div_frac_out_shl1_dbl}}
			    & {div_frac_out[53:0], (!div_frac_add[54])})
		| ({55{div_frac_out_shl1_sng}}
			    & {div_frac_out[53:29], (!div_frac_add[54]), 29'b0})
		| ({55{div_frac_out_of}}
			    & {55{d7stg_to_0}});
dffe_s #(55) i_div_frac_out (
	.din	(div_frac_out_in[54:0]),
	.en	(div_frac_out_load),
	.clk    (clk),
        .q      (div_frac_out[54:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign div_frac_out_54_53[1:0] = div_frac_out[54:53];
assign div_frac_outa[51:0]= div_frac_out[51:0];
endmodule
module fpu_in (
	pcx_fpio_data_rdy_px2,
	pcx_fpio_data_px2,
	a1stg_step,
	m1stg_step,
	d1stg_step,
	add_pipe_active,
	mul_pipe_active,
	div_pipe_active,
	inq_dout,
	sehold,
	arst_l,
	grst_l,
	rclk,
	fadd_clken_l,
	fmul_clken_l,
	fdiv_clken_l,
	
	inq_add,
	inq_mul,
	inq_div,
	inq_id,
	inq_rnd_mode,
	inq_fcc,
	inq_op,
	inq_in1_exp_neq_ffs,
	inq_in1_exp_eq_0,
	inq_in1_53_0_neq_0,
	inq_in1_50_0_neq_0,
	inq_in1_53_32_neq_0,
	inq_in1,
	inq_in2_exp_neq_ffs,
	inq_in2_exp_eq_0,
	inq_in2_53_0_neq_0,
	inq_in2_50_0_neq_0,
	inq_in2_53_32_neq_0,
	inq_in2,
	fp_id_in,
	fp_rnd_mode_in,
	fp_fcc_in,
	fp_op_in,
	fp_src1_in,
	fp_src2_in,
	inq_rdaddr,
	inq_wraddr,
	inq_read_en,
	inq_we,
	se,
	si,
	so
);
input		pcx_fpio_data_rdy_px2;	
input [123:0]	pcx_fpio_data_px2;	
input		a1stg_step;		
input		m1stg_step;		
input		d1stg_step;		
input 		add_pipe_active;        
input 		mul_pipe_active;        
input 		div_pipe_active;        
input [154:0] inq_dout; 
input sehold; 
input		arst_l;			
input		grst_l;			
input		rclk;			
output		fadd_clken_l;		
output		fmul_clken_l;		
output		fdiv_clken_l;		
output		inq_add;		
output		inq_mul;		
output		inq_div;		
output [4:0]	inq_id;			
output [1:0]	inq_rnd_mode;		
output [1:0]	inq_fcc;		
output [7:0]	inq_op;			
output		inq_in1_exp_neq_ffs;	
output		inq_in1_exp_eq_0;	
output		inq_in1_53_0_neq_0;	
output		inq_in1_50_0_neq_0;	
output		inq_in1_53_32_neq_0;	
output [63:0]	inq_in1;		
output		inq_in2_exp_neq_ffs;	
output		inq_in2_exp_eq_0;	
output		inq_in2_53_0_neq_0;	
output		inq_in2_50_0_neq_0;	
output		inq_in2_53_32_neq_0;	
output [63:0]	inq_in2;		
output [4:0] fp_id_in; 
output [1:0] fp_rnd_mode_in; 
output [1:0] fp_fcc_in; 
output [7:0] fp_op_in; 
output [68:0] fp_src1_in; 
output [68:0] fp_src2_in; 
output [3:0] inq_rdaddr; 
output [3:0] inq_wraddr; 
output inq_read_en; 
output inq_we; 
input           se;                     
input           si;                     
output          so;                     
wire		inq_we;			
wire [3:0]	inq_wraddr;		
wire            inq_read_en;            
wire [3:0]	inq_rdaddr;		
wire		inq_bp;			
wire		inq_bp_inv;		
wire		inq_fwrd;		
wire		inq_fwrd_inv;		
wire		inq_add;		
wire		inq_mul;		
wire		inq_div;		
wire  		fadd_clken_l;		
wire 		fmul_clken_l;		
wire 		fdiv_clken_l;		
wire [7:0]	fp_op_in;		
wire            fp_op_in_7in;           
wire [4:0]	inq_id;			
wire [1:0]	inq_rnd_mode;		
wire [1:0]	inq_fcc;		
wire [7:0]	inq_op;			
wire		inq_in1_exp_neq_ffs;	
wire		inq_in1_exp_eq_0;	
wire		inq_in1_53_0_neq_0;	
wire		inq_in1_50_0_neq_0;	
wire		inq_in1_53_32_neq_0;	
wire [63:0]	inq_in1;		
wire		inq_in2_exp_neq_ffs;	
wire		inq_in2_exp_eq_0;	
wire		inq_in2_53_0_neq_0;	
wire		inq_in2_50_0_neq_0;	
wire		inq_in2_53_32_neq_0;	
wire [63:0]	inq_in2;		
wire [4:0] fp_id_in; 
wire [1:0] fp_rnd_mode_in; 
wire [1:0] fp_fcc_in; 
wire [68:0] fp_src1_in; 
wire [68:0] fp_src2_in; 
wire fp_data_rdy;
wire        scan_out_fpu_in_ctl;
fpu_in_ctl fpu_in_ctl (
	.pcx_fpio_data_rdy_px2		(pcx_fpio_data_rdy_px2),
	.pcx_fpio_data_px2		(pcx_fpio_data_px2[123:118]),
	.fp_op_in    			(fp_op_in[3:2]),
        .fp_op_in_7in                   (fp_op_in_7in),
	.a1stg_step			(a1stg_step),
	.m1stg_step			(m1stg_step),
	.d1stg_step			(d1stg_step),
	.add_pipe_active		(add_pipe_active),
	.mul_pipe_active		(mul_pipe_active),
	.div_pipe_active		(div_pipe_active),
	.sehold (sehold),
	.arst_l				(arst_l),
	.grst_l				(grst_l),
	.rclk			(rclk),
        .fp_data_rdy			(fp_data_rdy),
	.fadd_clken_l			(fadd_clken_l),
	.fmul_clken_l			(fmul_clken_l),
	.fdiv_clken_l			(fdiv_clken_l),
	.inq_we				(inq_we),
	.inq_wraddr			(inq_wraddr[3:0]),
	.inq_read_en			(inq_read_en),
	.inq_rdaddr			(inq_rdaddr[3:0]),
	.inq_bp				(inq_bp),
	.inq_bp_inv			(inq_bp_inv),
	.inq_fwrd			(inq_fwrd),
	.inq_fwrd_inv			(inq_fwrd_inv),
	.inq_add			(inq_add),
	.inq_mul			(inq_mul),
	.inq_div			(inq_div),
	.se           (se),
  .si           (si),
  .so           (scan_out_fpu_in_ctl)
);
fpu_in_dp fpu_in_dp (
        .fp_data_rdy			(fp_data_rdy),
        .fpio_data_px2_116_112          (pcx_fpio_data_px2[116:112]),
        .fpio_data_px2_79_72            (pcx_fpio_data_px2[79:72]),
        .fpio_data_px2_67_0             (pcx_fpio_data_px2[67:0]),
	.inq_fwrd			(inq_fwrd),
	.inq_fwrd_inv			(inq_fwrd_inv),
	.inq_bp				(inq_bp),
	.inq_bp_inv			(inq_bp_inv),
	.inq_dout    (inq_dout[154:0]),
	.rclk			(rclk),
        .fp_op_in_7in                   (fp_op_in_7in),
	.inq_id				(inq_id[4:0]),
	.inq_rnd_mode			(inq_rnd_mode[1:0]),
	.inq_fcc			(inq_fcc[1:0]),
	.inq_op				(inq_op[7:0]),
	.inq_in1_exp_neq_ffs		(inq_in1_exp_neq_ffs),
	.inq_in1_exp_eq_0		(inq_in1_exp_eq_0),
	.inq_in1_53_0_neq_0		(inq_in1_53_0_neq_0),
	.inq_in1_50_0_neq_0		(inq_in1_50_0_neq_0),
	.inq_in1_53_32_neq_0		(inq_in1_53_32_neq_0),
	.inq_in1			(inq_in1[63:0]),
	.inq_in2_exp_neq_ffs		(inq_in2_exp_neq_ffs),
	.inq_in2_exp_eq_0		(inq_in2_exp_eq_0),
	.inq_in2_53_0_neq_0		(inq_in2_53_0_neq_0),
	.inq_in2_50_0_neq_0		(inq_in2_50_0_neq_0),
	.inq_in2_53_32_neq_0		(inq_in2_53_32_neq_0),
	.inq_in2			(inq_in2[63:0]),
	.fp_id_in (fp_id_in[4:0]),
	.fp_rnd_mode_in (fp_rnd_mode_in[1:0]),
	.fp_fcc_in (fp_fcc_in[1:0]),
	.fp_op_in (fp_op_in[7:0]),
	.fp_src1_in (fp_src1_in[68:0]),
	.fp_src2_in (fp_src2_in[68:0]),
	.se                             (se),
        .si                             (scan_out_fpu_in_ctl),
        .so                             (so)
);
endmodule
 
module fpu_in_ctl (
	pcx_fpio_data_rdy_px2,
	pcx_fpio_data_px2,
	fp_op_in,
        fp_op_in_7in,
	a1stg_step,
	m1stg_step,
	d1stg_step,
	add_pipe_active,
	mul_pipe_active,
	div_pipe_active,
	sehold,
	arst_l,
	grst_l,
	rclk,
        fp_data_rdy,
	fadd_clken_l,
	fmul_clken_l,
	fdiv_clken_l,
	
	inq_we,
	inq_wraddr,
	inq_read_en,
	inq_rdaddr,
	inq_bp,
	inq_bp_inv,
	inq_fwrd,
	inq_fwrd_inv,
	inq_add,
	inq_mul,
	inq_div,
	se,
	si,
	so
);
input		pcx_fpio_data_rdy_px2;	
input [123:118]	pcx_fpio_data_px2;	
input [3:2]	fp_op_in;		
input         	fp_op_in_7in;		
input		a1stg_step;		
input		m1stg_step;		
input		d1stg_step;		
input 		add_pipe_active;        
input 		mul_pipe_active;        
input 		div_pipe_active;        
input sehold; 
input		arst_l;			
input		grst_l;			
input		rclk;		
output          fp_data_rdy;
output		fadd_clken_l;		
output		fmul_clken_l;		
output		fdiv_clken_l;		
output		inq_we;			
output [3:0]	inq_wraddr;		
output          inq_read_en;            
output [3:0]	inq_rdaddr;		
output		inq_bp;			
output		inq_bp_inv;		
output		inq_fwrd;		
output		inq_fwrd_inv;		
output		inq_add;		
output		inq_mul;		
output		inq_div;		
input           se;                     
input           si;                     
output          so;                     
wire		reset;
wire		fp_data_rdy;
wire		fp_vld_in;
wire [4:0]	fp_type_in;
wire  		fadd_clken_l;
wire 		fmul_clken_l;
wire 		fdiv_clken_l;
wire		fp_op_in_7;
wire		fp_op_in_7_inv;
wire		inq_we;
wire            inq_read_en;
wire [3:0]	inq_wrptr_plus1;
wire		inq_wrptr_step;
wire [3:0]	inq_wrptr;
wire [3:0]	inq_div_wrptr_plus1;
wire		inq_div_wrptr_step;
wire [3:0]	inq_div_wrptr;
wire [3:0]	inq_wraddr;
wire [3:0]	inq_wraddr_del;
wire		inq_re;
wire [3:0]	inq_rdptr_plus1;
wire [3:0]	inq_rdptr_in;
wire [3:0]	inq_rdptr;
wire		inq_div_re;
wire [3:0]	inq_div_rdptr_plus1;
wire [3:0]	inq_div_rdptr_in;
wire [3:0]	inq_div_rdptr;
wire		inq_div_rd_in;
wire		inq_div_rd;
wire [3:0]	inq_rdaddr;
wire [3:0]	inq_rdaddr_del;
wire		inq_bp;
wire		inq_bp_inv;
wire		inq_empty;
wire		inq_div_empty;
wire		inq_fwrd;
wire		inq_fwrd_inv;
wire		fp_add_in;
wire		fp_mul_in;
wire		fp_div_in;
wire [7:0]	inq_rdptr_dec_in;
wire [7:0]	inq_rdptr_dec;
wire [7:0]	inq_div_rdptr_dec_in;
wire [7:0]	inq_div_rdptr_dec;
wire [15:0]	inq_rdaddr_del_dec_in;
wire [15:0]	inq_rdaddr_del_dec;
wire		inq_pipe0_we;
wire		inq_pipe1_we;
wire		inq_pipe2_we;
wire		inq_pipe3_we;
wire		inq_pipe4_we;
wire		inq_pipe5_we;
wire		inq_pipe6_we;
wire		inq_pipe7_we;
wire		inq_pipe8_we;
wire		inq_pipe9_we;
wire		inq_pipe10_we;
wire		inq_pipe11_we;
wire		inq_pipe12_we;
wire		inq_pipe13_we;
wire		inq_pipe14_we;
wire		inq_pipe15_we;
wire [2:0]	inq_pipe0;
wire [2:0]	inq_pipe1;
wire [2:0]	inq_pipe2;
wire [2:0]	inq_pipe3;
wire [2:0]	inq_pipe4;
wire [2:0]	inq_pipe5;
wire [2:0]	inq_pipe6;
wire [2:0]	inq_pipe7;
wire [2:0]	inq_pipe8;
wire [2:0]	inq_pipe9;
wire [2:0]	inq_pipe10;
wire [2:0]	inq_pipe11;
wire [2:0]	inq_pipe12;
wire [2:0]	inq_pipe13;
wire [2:0]	inq_pipe14;
wire [2:0]	inq_pipe15;
wire [2:0]	inq_pipe;
wire		inq_div;
wire		inq_diva;
wire		inq_diva_dly;
wire		d1stg_step_dly;
wire		inq_mul;
wire		inq_mula;
wire		inq_add;
wire		inq_adda;
wire		valid_packet;
wire            valid_packet_dly;
wire		tag_sel;
wire sehold_inv;
wire        in_ctl_rst_l;
wire        inq_adda_dly;
wire        inq_mula_dly;
dffrl_async #(1)  dffrl_in_ctl (
  .din  (grst_l),
  .clk  (rclk),
  .rst_l(arst_l),
  .q    (in_ctl_rst_l),
	.se (se),
	.si (),
	.so ()
  );
assign reset= (!in_ctl_rst_l);
dffr_s #(1) i_fp_data_rdy (
	.din	(pcx_fpio_data_rdy_px2),
	.rst    (reset),
        .clk    (rclk),
        .q      (fp_data_rdy),
	.se     (se),
        .si     (),
        .so     ()
);
dff_s #(1) i_fp_vld_in (
	.din	(pcx_fpio_data_px2[123]),
	.clk    (rclk),
        .q      (fp_vld_in),
	.se     (se),
        .si     (),
        .so     ()
);
dff_s #(5) i_fp_type_in (
	.din	(pcx_fpio_data_px2[122:118]),
        .clk    (rclk),
 
        .q      (fp_type_in[4:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign fp_op_in_7= fp_op_in_7in;
assign fp_op_in_7_inv= (!fp_op_in_7);
assign inq_we= fp_data_rdy && fp_vld_in
		&& (((fp_type_in[4:0]==5'h0a) && fp_op_in_7)
			|| ((fp_type_in[4:0]==5'h0b) && fp_op_in_7_inv));
assign inq_wrptr_plus1[3:0]= inq_wrptr[3:0] + 4'h1;
assign inq_wrptr_step= inq_we && (!fp_div_in);
dffre_s #(4) i_inq_wrptr (
	.din	(inq_wrptr_plus1[3:0]),
	.en	(inq_wrptr_step),
	.rst	(reset),
	.clk    (rclk),
        .q      (inq_wrptr[3:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign inq_div_wrptr_plus1[3:0]= inq_div_wrptr[3:0] + 4'h1;
assign inq_div_wrptr_step= inq_we && fp_div_in;
dffre_s #(4) i_inq_div_wrptr (
        .din    (inq_div_wrptr_plus1[3:0]),
        .en     (inq_div_wrptr_step),
        .rst    (reset),
        .clk    (rclk),
 
        .q      (inq_div_wrptr[3:0]),
 
        .se     (se),
        .si     (),
        .so     ()
);
assign inq_wraddr[3:0]= {fp_div_in,
		(({3{fp_div_in}}
			    & inq_div_wrptr[2:0])
		    | ({3{(!fp_div_in)}}
			    & inq_wrptr[2:0]))};
dff_s #(4) i_inq_wraddr_del (
	.din	(inq_wraddr[3:0]),
	.clk	(rclk),
	.q	(inq_wraddr_del[3:0]),
	.se	(se),
	.si	(),
	.so	()
);
assign inq_read_en = ~inq_empty | ~inq_div_empty;
assign inq_re= (inq_adda && a1stg_step)
		|| (inq_mula && m1stg_step);
assign inq_rdptr_plus1[3:0]= inq_rdptr[3:0] + 4'h1;
assign inq_rdptr_in[3:0]= ({4{(inq_re && (!reset))}}
			    & inq_rdptr_plus1[3:0])
		| ({4{((!inq_re) && (!reset))}}
			    & inq_rdptr[3:0]);
dff_s #(4) i_inq_rdptr (
	.din	(inq_rdptr_in[3:0]),
	.clk    (rclk),
 
        .q      (inq_rdptr[3:0]),
 
        .se     (se),
        .si     (),
        .so     ()
);
assign inq_div_re= (inq_diva && d1stg_step);
assign inq_div_rdptr_plus1[3:0]= inq_div_rdptr[3:0] + 4'h1;
assign inq_div_rdptr_in[3:0]= ({4{(inq_div_re && (!reset))}}
                            & inq_div_rdptr_plus1[3:0])
                | ({4{((!inq_div_re) && (!reset))}}
                            & inq_div_rdptr[3:0]);
 
dff_s #(4) i_inq_div_rdptr (
        .din    (inq_div_rdptr_in[3:0]),
        .clk    (rclk),
        .q      (inq_div_rdptr[3:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign inq_div_rd_in= (!inq_div_empty) && d1stg_step && (!inq_diva);
dff_s #(1) i_inq_div_rd (
	.din	(inq_div_rd_in),
	.clk    (rclk),
        .q      (inq_div_rd),
        .se     (se),
        .si     (),
        .so     ()
);
assign inq_rdaddr[3:0]= {inq_div_rd_in,
		(({3{inq_div_rd_in}}
			    & (inq_div_rdptr[2:0] & {3{(!reset)}}))
		    | ({3{(!inq_div_rd_in)}}
			    & inq_rdptr_in[2:0]))};
dff_s #(4) i_inq_rdaddr_del (
	.din	(inq_rdaddr[3:0]),
        .clk	(rclk),
 
        .q	(inq_rdaddr_del[3:0]),
 
        .se	(se),
        .si	(),
        .so	()
);
assign valid_packet = fp_data_rdy && fp_vld_in &&
                      ((fp_type_in[4:0]==5'h0a) || (fp_type_in[4:0]==5'h0b));
dffre_s #(1) i_valid_packet_dly (
	.din	(valid_packet),
	.en     (1'b1),
        .rst    (reset),
        .clk    (rclk),
        .q      (valid_packet_dly),
        .se     (se),
        .si     (),
        .so     ()
);
assign sehold_inv = ~sehold;
assign inq_bp= (inq_wraddr_del[3:0]==inq_rdaddr_del[3:0]) && valid_packet_dly && sehold_inv;
assign inq_bp_inv= (!inq_bp);
assign inq_empty= (inq_wrptr[3:0]==inq_rdptr[3:0]);
assign inq_div_empty= (inq_div_wrptr[3:0]==inq_div_rdptr[3:0]);
assign inq_fwrd= ((inq_empty && (!inq_div_rd))
  		|| (inq_div_empty && fp_div_in
  			&& d1stg_step)) && valid_packet && sehold_inv;
assign inq_fwrd_inv= (!inq_fwrd);
assign fp_add_in= fp_data_rdy && fp_vld_in && (fp_type_in[4:1]==4'h5)
		&& ((fp_op_in_7 && (!fp_type_in[0]))
			|| (fp_op_in_7_inv && (!fp_op_in[3]) && fp_type_in[0]));
assign fp_mul_in= fp_data_rdy && fp_vld_in && (fp_type_in[4:0]==5'h0b)
		&& fp_op_in_7_inv && (fp_op_in[3:2]==2'b10);
assign fp_div_in= fp_data_rdy && fp_vld_in && (fp_type_in[4:0]==5'h0b)
                && fp_op_in_7_inv && (fp_op_in[3:2]==2'b11);
assign inq_rdptr_dec_in[7:0]= ({8{reset}}
			    & 8'h01)
		| ({8{(inq_re && (!reset))}}
			    & {inq_rdptr_dec[6:0], inq_rdptr_dec[7]})
		| ({8{((!inq_re) && (!reset))}}
			    & inq_rdptr_dec[7:0]);
dff_s #(8) i_inq_rdptr_dec (
	.din	(inq_rdptr_dec_in[7:0]),
	.clk	(rclk),
	.q	(inq_rdptr_dec[7:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign inq_div_rdptr_dec_in[7:0]= ({8{reset}}
                            & 8'h01)
                | ({8{(inq_div_re && (!reset))}}
                            & {inq_div_rdptr_dec[6:0], inq_div_rdptr_dec[7]})
                | ({8{((!inq_div_re) && (!reset))}}
                            & inq_div_rdptr_dec[7:0]);
 
dff_s #(8) i_inq_div_rdptr_dec (
        .din    (inq_div_rdptr_dec_in[7:0]),
        .clk    (rclk),
        .q      (inq_div_rdptr_dec[7:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign inq_rdaddr_del_dec_in[15:0]= ({16{((!inq_div_empty) && d1stg_step
					&& (!inq_diva))}}
			    & {(inq_div_rdptr_dec[7:1] & {7{(!reset)}}),
				(inq_div_rdptr_dec[0] || reset), 8'b0})
		| ({16{(!((!inq_div_empty) && d1stg_step && (!inq_diva)))}}
			    & {8'b0, inq_rdptr_dec_in[7:0]});
dff_s #(16) i_inq_rdaddr_del_dec (
	.din	(inq_rdaddr_del_dec_in[15:0]),
	.clk	(rclk),
	.q	(inq_rdaddr_del_dec[15:0]),
 
        .se     (se),
        .si     (),
        .so     ()
);
assign inq_pipe0_we= inq_we && (!fp_div_in) && (inq_wrptr[2:0]==3'h0);
assign inq_pipe1_we= inq_we && (!fp_div_in) && (inq_wrptr[2:0]==3'h1);
assign inq_pipe2_we= inq_we && (!fp_div_in) && (inq_wrptr[2:0]==3'h2);
assign inq_pipe3_we= inq_we && (!fp_div_in) && (inq_wrptr[2:0]==3'h3);
assign inq_pipe4_we= inq_we && (!fp_div_in) && (inq_wrptr[2:0]==3'h4);
assign inq_pipe5_we= inq_we && (!fp_div_in) && (inq_wrptr[2:0]==3'h5);
assign inq_pipe6_we= inq_we && (!fp_div_in) && (inq_wrptr[2:0]==3'h6);
assign inq_pipe7_we= inq_we && (!fp_div_in) && (inq_wrptr[2:0]==3'h7);
assign inq_pipe8_we= inq_we && fp_div_in && (inq_div_wrptr[2:0]==3'h0);
assign inq_pipe9_we= inq_we && fp_div_in && (inq_div_wrptr[2:0]==3'h1);
assign inq_pipe10_we= inq_we && fp_div_in && (inq_div_wrptr[2:0]==3'h2);
assign inq_pipe11_we= inq_we && fp_div_in && (inq_div_wrptr[2:0]==3'h3);
assign inq_pipe12_we= inq_we && fp_div_in && (inq_div_wrptr[2:0]==3'h4);
assign inq_pipe13_we= inq_we && fp_div_in && (inq_div_wrptr[2:0]==3'h5);
assign inq_pipe14_we= inq_we && fp_div_in && (inq_div_wrptr[2:0]==3'h6);
assign inq_pipe15_we= inq_we && fp_div_in && (inq_div_wrptr[2:0]==3'h7);
dffre_s #(3) i_inq_pipe0 (
	.din	({fp_div_in, fp_mul_in, fp_add_in}),
	.en	(inq_pipe0_we),
        .rst    (reset),
	.clk    (rclk),
        .q      (inq_pipe0[2:0]),
 
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(3) i_inq_pipe1 (
        .din    ({fp_div_in, fp_mul_in, fp_add_in}),
        .en     (inq_pipe1_we),
        .rst    (reset),
        .clk    (rclk),
        .q      (inq_pipe1[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(3) i_inq_pipe2 (
        .din    ({fp_div_in, fp_mul_in, fp_add_in}),
        .en     (inq_pipe2_we),
        .rst    (reset),
        .clk    (rclk),
        .q      (inq_pipe2[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(3) i_inq_pipe3 (
        .din    ({fp_div_in, fp_mul_in, fp_add_in}),
        .en     (inq_pipe3_we),
        .rst    (reset),
        .clk    (rclk),
        .q      (inq_pipe3[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(3) i_inq_pipe4 (
        .din    ({fp_div_in, fp_mul_in, fp_add_in}),
        .en     (inq_pipe4_we),
        .rst    (reset),
        .clk    (rclk),
        .q      (inq_pipe4[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(3) i_inq_pipe5 (
        .din    ({fp_div_in, fp_mul_in, fp_add_in}),
        .en     (inq_pipe5_we),
        .rst    (reset),
        .clk    (rclk),
        .q      (inq_pipe5[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(3) i_inq_pipe6 (
        .din    ({fp_div_in, fp_mul_in, fp_add_in}),
        .en     (inq_pipe6_we),
        .rst    (reset),
        .clk    (rclk),
        .q      (inq_pipe6[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(3) i_inq_pipe7 (
        .din    ({fp_div_in, fp_mul_in, fp_add_in}),
        .en     (inq_pipe7_we),
        .rst    (reset),
        .clk    (rclk),
        .q      (inq_pipe7[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(3) i_inq_pipe8 (
        .din    ({fp_div_in, fp_mul_in, fp_add_in}),
        .en     (inq_pipe8_we),
        .rst    (reset),
        .clk    (rclk),
        .q      (inq_pipe8[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(3) i_inq_pipe9 (
        .din    ({fp_div_in, fp_mul_in, fp_add_in}),
        .en     (inq_pipe9_we),
        .rst    (reset),
        .clk    (rclk),
        .q      (inq_pipe9[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(3) i_inq_pipe10 (
        .din    ({fp_div_in, fp_mul_in, fp_add_in}),
        .en     (inq_pipe10_we),
        .rst    (reset),
        .clk    (rclk),
        .q      (inq_pipe10[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(3) i_inq_pipe11 (
        .din    ({fp_div_in, fp_mul_in, fp_add_in}),
        .en     (inq_pipe11_we),
        .rst    (reset),
        .clk    (rclk),
        .q      (inq_pipe11[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(3) i_inq_pipe12 (
        .din    ({fp_div_in, fp_mul_in, fp_add_in}),
        .en     (inq_pipe12_we),
        .rst    (reset),
        .clk    (rclk),
        .q      (inq_pipe12[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(3) i_inq_pipe13 (
        .din    ({fp_div_in, fp_mul_in, fp_add_in}),
        .en     (inq_pipe13_we),
        .rst    (reset),
        .clk    (rclk),
        .q      (inq_pipe13[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(3) i_inq_pipe14 (
        .din    ({fp_div_in, fp_mul_in, fp_add_in}),
        .en     (inq_pipe14_we),
        .rst    (reset),
        .clk    (rclk),
        .q      (inq_pipe14[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(3) i_inq_pipe15 (
        .din    ({fp_div_in, fp_mul_in, fp_add_in}),
        .en     (inq_pipe15_we),
        .rst    (reset),
        .clk    (rclk),
        .q      (inq_pipe15[2:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign tag_sel = (inq_empty && (!inq_div_rd))
  		|| (inq_div_empty && fp_div_in && fp_data_rdy && fp_vld_in
  			&& d1stg_step);
assign inq_pipe[2:0]= ({3{tag_sel}}
                                
                                
			    & {(inq_div_empty && fp_div_in && fp_data_rdy && fp_vld_in
				&& d1stg_step
				&& d1stg_step_dly && (!inq_diva_dly)),
                                fp_mul_in,
				fp_add_in})
		| ({3{(!tag_sel)}}
			    & (({3{inq_rdaddr_del_dec[0]}}
					& inq_pipe0[2:0])
				| ({3{inq_rdaddr_del_dec[1]}}
                                        & inq_pipe1[2:0])
                                | ({3{inq_rdaddr_del_dec[2]}}
                                        & inq_pipe2[2:0])
                                | ({3{inq_rdaddr_del_dec[3]}}
                                        & inq_pipe3[2:0])
                                | ({3{inq_rdaddr_del_dec[4]}}
                                        & inq_pipe4[2:0])
                                | ({3{inq_rdaddr_del_dec[5]}}
                                        & inq_pipe5[2:0])
                                | ({3{inq_rdaddr_del_dec[6]}}
                                        & inq_pipe6[2:0])
                                | ({3{inq_rdaddr_del_dec[7]}}
                                        & inq_pipe7[2:0])
                                | ({3{inq_rdaddr_del_dec[8]}}
                                        & inq_pipe8[2:0])
                                | ({3{inq_rdaddr_del_dec[9]}}
                                        & inq_pipe9[2:0])
                                | ({3{inq_rdaddr_del_dec[10]}}
                                        & inq_pipe10[2:0])
                                | ({3{inq_rdaddr_del_dec[11]}}
                                        & inq_pipe11[2:0])
                                | ({3{inq_rdaddr_del_dec[12]}}
                                        & inq_pipe12[2:0])
                                | ({3{inq_rdaddr_del_dec[13]}}
                                        & inq_pipe13[2:0])
                                | ({3{inq_rdaddr_del_dec[14]}}
                                        & inq_pipe14[2:0])
                                | ({3{inq_rdaddr_del_dec[15]}}
                                        & inq_pipe15[2:0])));
assign inq_div= inq_pipe[2];
assign inq_diva= inq_pipe[2];
assign inq_mul= inq_pipe[1];
assign inq_mula= inq_pipe[1];
assign inq_add= inq_pipe[0];
assign inq_adda= inq_pipe[0];
dffre_s #(1) i_inq_adda_dly (
	.din	(inq_adda),
	.en     (1'b1),
        .rst    (reset),
        .clk    (rclk),
        .q      (inq_adda_dly),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(1) i_inq_mula_dly (
	.din	(inq_mula),
	.en     (1'b1),
        .rst    (reset),
        .clk    (rclk),
        .q      (inq_mula_dly),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(1) i_inq_diva_dly (
	.din	(inq_diva),
	.en     (1'b1),
        .rst    (reset),
        .clk    (rclk),
        .q      (inq_diva_dly),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(1) i_d1stg_step_dly (
	.din	(d1stg_step),
	.en     (1'b1),
        .rst    (reset),
        .clk    (rclk),
        .q      (d1stg_step_dly),
        .se     (se),
        .si     (),
        .so     ()
);
assign fadd_clken_l = !(add_pipe_active || inq_adda || inq_adda_dly || reset);
assign fmul_clken_l = !(mul_pipe_active || inq_mula || inq_mula_dly || reset);
assign fdiv_clken_l = !(div_pipe_active || inq_diva || inq_diva_dly || reset);
endmodule
module fpu_in_dp (
	fp_data_rdy,
        fpio_data_px2_116_112,
        fpio_data_px2_79_72,
        fpio_data_px2_67_0,
	inq_fwrd,
	inq_fwrd_inv,
	inq_bp,
	inq_bp_inv,
	inq_dout,
	rclk,
	
        fp_op_in_7in,
	inq_id,
	inq_rnd_mode,
	inq_fcc,
	inq_op,
	inq_in1_exp_neq_ffs,
	inq_in1_exp_eq_0,
	inq_in1_53_0_neq_0,
	inq_in1_50_0_neq_0,
	inq_in1_53_32_neq_0,
	inq_in1,
	inq_in2_exp_neq_ffs,
	inq_in2_exp_eq_0,
	inq_in2_53_0_neq_0,
	inq_in2_50_0_neq_0,
	inq_in2_53_32_neq_0,
	inq_in2,
	fp_id_in,
	fp_rnd_mode_in,
	fp_fcc_in,
	fp_op_in,
	fp_src1_in,
	fp_src2_in,
	se,
	si,
	so
);
input           fp_data_rdy;
input [116:112] fpio_data_px2_116_112;  
input [79:72]   fpio_data_px2_79_72;    
input [67:0]    fpio_data_px2_67_0;     
input		inq_fwrd;		
input		inq_fwrd_inv;		
input		inq_bp;			
input		inq_bp_inv;		
input [154:0] inq_dout; 
input		rclk;		
output          fp_op_in_7in;           
output [4:0]	inq_id;			
output [1:0]	inq_rnd_mode;		
output [1:0]	inq_fcc;		
output [7:0]	inq_op;			
output		inq_in1_exp_neq_ffs;	
output		inq_in1_exp_eq_0;	
output		inq_in1_53_0_neq_0;	
output		inq_in1_50_0_neq_0;	
output		inq_in1_53_32_neq_0;	
output [63:0]	inq_in1;		
output		inq_in2_exp_neq_ffs;	
output		inq_in2_exp_eq_0;	
output		inq_in2_53_0_neq_0;	
output		inq_in2_50_0_neq_0;	
output		inq_in2_53_32_neq_0;	
output [63:0]	inq_in2;		
output [4:0] fp_id_in; 
output [1:0] fp_rnd_mode_in; 
output [1:0] fp_fcc_in; 
output [7:0] fp_op_in; 
output [68:0] fp_src1_in; 
output [68:0] fp_src2_in; 
input           se;                     
input           si;                     
output          so;                     
wire [154:0]	inq_dout;
wire [4:0]	fp_id_in;
wire [7:0]	fp_op_in;
wire		fp_op_in_7;		
wire		fp_op_in_7_inv;		
wire            fp_op_in_7in;
wire [1:0]	fp_fcc_in;
wire [1:0]	fp_rnd_mode_in;
wire [63:0]	fp_srca_in;
wire		fp_srca_53_0_neq_0;
wire		fp_srca_50_0_neq_0;
wire		fp_srca_53_32_neq_0;
wire		fp_srca_exp_eq_0;
wire		fp_srca_exp_neq_ffs;
wire [68:0]	fp_srcb_in;
wire [68:0]	fp_src1_in;
wire [68:0]	fp_src2_in;
wire [154:0]	inq_din_d1;
wire [154:0]	inq_data;
wire [4:0]	inq_id;
wire [1:0]	inq_rnd_mode;
wire [1:0]	inq_fcc;
wire [7:0]	inq_op;
wire		inq_in1_exp_neq_ffs;
wire		inq_in1_exp_eq_0;
wire		inq_in1_53_0_neq_0;
wire		inq_in1_50_0_neq_0;
wire		inq_in1_53_32_neq_0;
wire [63:0]	inq_in1;
wire		inq_in2_exp_neq_ffs;
wire		inq_in2_exp_eq_0;
wire		inq_in2_53_0_neq_0;
wire		inq_in2_50_0_neq_0;
wire		inq_in2_53_32_neq_0;
wire [63:0]	inq_in2;
wire clk;
wire se_l;
assign se_l = ~se;
clken_buf  ckbuf_in_dp (
  .clk(clk),
  .rclk(rclk),
  .enb_l(1'b0),
  .tmb_l(se_l)
  );
dff_s #(5) i_fp_id_in (
	.din	(fpio_data_px2_116_112[116:112]),
	.clk    (clk),
 
        .q      (fp_id_in[4:0]),
 
        .se     (se),
        .si     (),
        .so     ()
);
dff_s #(8) i_fp_op_in (
        .din    (fpio_data_px2_79_72[79:72]),
        .clk    (clk),
        .q      (fp_op_in[7:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign fp_op_in_7in = fp_op_in[7];
assign fp_op_in_7 = fp_op_in[7];
assign fp_op_in_7_inv = ~fp_op_in[7];
dff_s #(2) i_fp_fcc_in (
        .din    (fpio_data_px2_67_0[67:66]),
        .clk    (clk),
        .q      (fp_fcc_in[1:0]),
 
        .se     (se),
        .si     (),
        .so     ()
);
dff_s #(2) i_fp_rnd_mode_in (
        .din    (fpio_data_px2_67_0[65:64]),
        .clk    (clk),
        .q      (fp_rnd_mode_in[1:0]),
 
        .se     (se),
        .si     (),
        .so     ()
);
dff_s #(64) i_fp_srca_in (
	.din    (fpio_data_px2_67_0[63:0]),
        .clk    (clk),
        .q      (fp_srca_in[63:0]),
 
        .se     (se),
        .si     (),
        .so     ()
);
assign fp_srca_53_0_neq_0= (|fp_srca_in[53:0]);
assign fp_srca_50_0_neq_0= (|fp_srca_in[50:0]);
assign fp_srca_53_32_neq_0= (|fp_srca_in[53:32]);
assign fp_srca_exp_eq_0= (!((|fp_srca_in[62:55])
		|| (fp_op_in[1] && (|fp_srca_in[54:52]))));
assign fp_srca_exp_neq_ffs= (!((&fp_srca_in[62:55])
		&& (fp_op_in[0] || (&fp_srca_in[54:52]))));
dffe_s #(69) i_fp_srcb_in (
	.din	({fp_srca_exp_neq_ffs, fp_srca_exp_eq_0, fp_srca_53_0_neq_0,
			fp_srca_50_0_neq_0, fp_srca_53_32_neq_0,
			fp_srca_in[63:0]}),
        .en     (fp_data_rdy),
	.clk    (clk),
        .q      (fp_srcb_in[68:0]),
 
        .se     (se),
        .si     (),
        .so     ()
);
assign fp_src1_in[68:0]= ({69{fp_op_in_7_inv}}
			    & {fp_srca_exp_neq_ffs, fp_srca_exp_eq_0,
				fp_srca_53_0_neq_0, fp_srca_50_0_neq_0,
				fp_srca_53_32_neq_0, fp_srca_in[63:0]})
		| ({69{fp_op_in_7}}
			    & 69'h180000000000000000);
assign fp_src2_in[68:0]= ({69{fp_op_in_7_inv}}
			    & fp_srcb_in[68:0])
		| ({69{fp_op_in_7}}
			    & {fp_srca_exp_neq_ffs, fp_srca_exp_eq_0,
				fp_srca_53_0_neq_0, fp_srca_50_0_neq_0,
				fp_srca_53_32_neq_0, fp_srca_in[63:0]});
dff_s #(155) i_inq_din_d1 (
	.din	({fp_id_in[4:0], fp_rnd_mode_in[1:0], fp_fcc_in[1:0],
                        fp_op_in[7:0], fp_src1_in[68:0], fp_src2_in[68:0]}),
	.clk    (clk),
        .q      (inq_din_d1[154:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign inq_data[154:0]= ({155{inq_fwrd}}
			    & {fp_id_in[4:0], fp_rnd_mode_in[1:0],
				fp_fcc_in[1:0], fp_op_in[7:0],
				fp_src1_in[68:0], fp_src2_in[68:0]})
		| ({155{inq_fwrd_inv}}
			    & (({155{inq_bp}}
					& inq_din_d1[154:0])
				| ({155{inq_bp_inv}}
					& inq_dout[154:0])));
assign inq_id[4:0]= inq_data[154:150];
assign inq_rnd_mode[1:0]= inq_data[149:148];
assign inq_fcc[1:0]= inq_data[147:146];
assign inq_op[7:0]= inq_data[145:138];
assign inq_in1_exp_neq_ffs= inq_data[137];
assign inq_in1_exp_eq_0= inq_data[136];
assign inq_in1_53_0_neq_0= inq_data[135];
assign inq_in1_50_0_neq_0= inq_data[134];
assign inq_in1_53_32_neq_0= inq_data[133];
assign inq_in1[63:0]= inq_data[132:69];
assign inq_in2_exp_neq_ffs= inq_data[68];
assign inq_in2_exp_eq_0= inq_data[67];
assign inq_in2_53_0_neq_0= inq_data[66];
assign inq_in2_50_0_neq_0= inq_data[65];
assign inq_in2_53_32_neq_0= inq_data[64];
assign inq_in2[63:0]= inq_data[63:0];
endmodule
module fpu_in2_gt_in1_2b (
	din1,
	din2,
	din2_neq_din1,
	din2_gt_din1
);
input [1:0]	din1;			
input [1:0]	din2;			
output		din2_neq_din1;		
output		din2_gt_din1;		
wire [1:0]	din2_eq_din1;
wire		din2_neq_din1;
wire		din2_gt_din1;
assign din2_eq_din1[1:0]= (~(din1 ^ din2));
assign din2_neq_din1= (!(&din2_eq_din1));
assign din2_gt_din1= ((!din1[1]) && din2[1])
		|| (din2_eq_din1[1] && (!din1[0]) && din2[0]);
endmodule
module fpu_in2_gt_in1_3b (
	din1,
	din2,
	din2_neq_din1,
	din2_gt_din1
);
input [2:0]	din1;			
input [2:0]	din2;			
output		din2_neq_din1;		
output		din2_gt_din1;		
wire [2:0]	din2_eq_din1;
wire		din2_neq_din1;
wire		din2_gt_din1;
assign din2_eq_din1[2:0]= (~(din1 ^ din2));
assign din2_neq_din1= (!(&din2_eq_din1));
assign din2_gt_din1= ((!din1[2]) && din2[2])
		|| (din2_eq_din1[2] && (!din1[1]) && din2[1])
		|| ((&din2_eq_din1[2:1]) && (!din1[0]) && din2[0]);
endmodule
module fpu_in2_gt_in1_3to1 (
	din2_neq_din1_hi,
	din2_gt_din1_hi,
	din2_neq_din1_mid,
	din2_gt_din1_mid,
	din2_neq_din1_lo,
	din2_gt_din1_lo,
	din2_neq_din1,
	din2_gt_din1
);
input		din2_neq_din1_hi;	
input		din2_gt_din1_hi;	
input		din2_neq_din1_mid;	
input		din2_gt_din1_mid;	
input		din2_neq_din1_lo;	
input		din2_gt_din1_lo;	
output		din2_neq_din1;		
output		din2_gt_din1;		
wire		din2_neq_din1;
wire		din2_gt_din1;
assign din2_neq_din1= din2_neq_din1_hi || din2_neq_din1_mid || din2_neq_din1_lo;
assign din2_gt_din1= (din2_neq_din1_hi && din2_gt_din1_hi)
		|| ((!din2_neq_din1_hi) && din2_neq_din1_mid
			&& din2_gt_din1_mid)
		|| ((!din2_neq_din1_hi) && (!din2_neq_din1_mid)
			&& din2_gt_din1_lo);
endmodule
module fpu_in2_gt_in1_frac (
	din1,
	din2,
	sngop,
	expadd11,
	expeq,
	din2_neq_din1,
	din2_gt_din1,
	din2_gt1_din1
);
input [54:0]	din1;			
input [54:0]	din2;			
input		sngop;			
input		expadd11;		
input		expeq;			
output		din2_neq_din1;		
output		din2_gt_din1;		
output		din2_gt1_din1;		
wire		din2_neq_din1_54_52;
wire		din2_gt_din1_54_52;
wire		din2_neq_din1_51_50;
wire		din2_gt_din1_51_50;
wire		din2_neq_din1_49_48;
wire		din2_gt_din1_49_48;
wire		din2_neq_din1_47_45;
wire		din2_gt_din1_47_45;
wire		din2_neq_din1_44_42;
wire		din2_gt_din1_44_42;
wire		din2_neq_din1_41_39;
wire		din2_gt_din1_41_39;
wire		din2_neq_din1_38_36;
wire		din2_gt_din1_38_36;
wire		din2_neq_din1_35_33;
wire		din2_gt_din1_35_33;
wire		din2_neq_din1_32_30;
wire		din2_gt_din1_32_30;
wire		din2_neq_din1_29_27;
wire		din2_gt_din1_29_27;
wire		din2_neq_din1_26_24;
wire		din2_gt_din1_26_24;
wire		din2_neq_din1_23_21;
wire		din2_gt_din1_23_21;
wire		din2_neq_din1_20_18;
wire		din2_gt_din1_20_18;
wire		din2_neq_din1_17_15;
wire		din2_gt_din1_17_15;
wire		din2_neq_din1_14_12;
wire		din2_gt_din1_14_12;
wire		din2_neq_din1_11_9;
wire		din2_gt_din1_11_9;
wire		din2_neq_din1_8_6;
wire		din2_gt_din1_8_6;
wire		din2_neq_din1_5_3;
wire		din2_gt_din1_5_3;
wire		din2_neq_din1_2_0;
wire		din2_gt_din1_2_0;
wire		din2_neq_din1_51_45;
wire		din2_gt_din1_51_45;
wire		din2_neq_din1_44_36;
wire		din2_gt_din1_44_36;
wire		din2_neq_din1_35_27;
wire		din2_gt_din1_35_27;
wire		din2_neq_din1_26_18;
wire		din2_gt_din1_26_18;
wire		din2_neq_din1_17_9;
wire		din2_gt_din1_17_9;
wire		din2_neq_din1_8_0;
wire		din2_gt_din1_8_0;
wire		din2_neq_din1_51_27;
wire		din2_gt_din1_51_27;
wire		din2_neq_din1_26_0;
wire		din2_gt_din1_26_0;
wire		din2_neq_din1;
wire		din2_gt_din1;
wire		din2_gt1_din1;
fpu_in2_gt_in1_3b fpu_in2_gt_in1_54_52 (
	.din1			(din1[54:52]),
	.din2			(din2[54:52]),
	.din2_neq_din1		(din2_neq_din1_54_52),
	.din2_gt_din1		(din2_gt_din1_54_52)
);
fpu_in2_gt_in1_2b fpu_in2_gt_in1_51_50 (
	.din1			(din1[51:50]),
	.din2			(din2[51:50]),
	.din2_neq_din1		(din2_neq_din1_51_50),
	.din2_gt_din1		(din2_gt_din1_51_50)
);
fpu_in2_gt_in1_2b fpu_in2_gt_in1_49_48 (
        .din1                   (din1[49:48]),
        .din2                   (din2[49:48]),
        .din2_neq_din1          (din2_neq_din1_49_48),
        .din2_gt_din1           (din2_gt_din1_49_48)
);
fpu_in2_gt_in1_3b fpu_in2_gt_in1_47_45 (
        .din1                   (din1[47:45]),
        .din2                   (din2[47:45]),
        .din2_neq_din1          (din2_neq_din1_47_45),
        .din2_gt_din1           (din2_gt_din1_47_45)
);
fpu_in2_gt_in1_3b fpu_in2_gt_in1_44_42 (
        .din1                   (din1[44:42]),
        .din2                   (din2[44:42]),
        .din2_neq_din1          (din2_neq_din1_44_42),
        .din2_gt_din1           (din2_gt_din1_44_42)
);
fpu_in2_gt_in1_3b fpu_in2_gt_in1_41_39 (
        .din1                   (din1[41:39]),
        .din2                   (din2[41:39]),
        .din2_neq_din1          (din2_neq_din1_41_39),
        .din2_gt_din1           (din2_gt_din1_41_39)
);
fpu_in2_gt_in1_3b fpu_in2_gt_in1_38_36 (
        .din1                   (din1[38:36]),
        .din2                   (din2[38:36]),
        .din2_neq_din1          (din2_neq_din1_38_36),
        .din2_gt_din1           (din2_gt_din1_38_36)
);
fpu_in2_gt_in1_3b fpu_in2_gt_in1_35_33 (
        .din1                   (din1[35:33]),
        .din2                   (din2[35:33]),
        .din2_neq_din1          (din2_neq_din1_35_33),
        .din2_gt_din1           (din2_gt_din1_35_33)
);
fpu_in2_gt_in1_3b fpu_in2_gt_in1_32_30 (
        .din1                   (din1[32:30]),
        .din2                   (din2[32:30]),
        .din2_neq_din1          (din2_neq_din1_32_30),
        .din2_gt_din1           (din2_gt_din1_32_30)
);
fpu_in2_gt_in1_3b fpu_in2_gt_in1_29_27 (
        .din1                   (din1[29:27]),
        .din2                   (din2[29:27]),
        .din2_neq_din1          (din2_neq_din1_29_27),
        .din2_gt_din1           (din2_gt_din1_29_27)
);
fpu_in2_gt_in1_3b fpu_in2_gt_in1_26_24 (
        .din1                   (din1[26:24]),
        .din2                   (din2[26:24]),
        .din2_neq_din1          (din2_neq_din1_26_24),
        .din2_gt_din1           (din2_gt_din1_26_24)
);
fpu_in2_gt_in1_3b fpu_in2_gt_in1_23_21 (
        .din1                   (din1[23:21]),
        .din2                   (din2[23:21]),
        .din2_neq_din1          (din2_neq_din1_23_21),
        .din2_gt_din1           (din2_gt_din1_23_21)
);
fpu_in2_gt_in1_3b fpu_in2_gt_in1_20_18 (
        .din1                   (din1[20:18]),
        .din2                   (din2[20:18]),
        .din2_neq_din1          (din2_neq_din1_20_18),
        .din2_gt_din1           (din2_gt_din1_20_18)
);
fpu_in2_gt_in1_3b fpu_in2_gt_in1_17_15 (
        .din1                   (din1[17:15]),
        .din2                   (din2[17:15]),
        .din2_neq_din1          (din2_neq_din1_17_15),
        .din2_gt_din1           (din2_gt_din1_17_15)
);
fpu_in2_gt_in1_3b fpu_in2_gt_in1_14_12 (
        .din1                   (din1[14:12]),
        .din2                   (din2[14:12]),
        .din2_neq_din1          (din2_neq_din1_14_12),
        .din2_gt_din1           (din2_gt_din1_14_12)
);
fpu_in2_gt_in1_3b fpu_in2_gt_in1_11_9 (
        .din1                   (din1[11:9]),
        .din2                   (din2[11:9]),
        .din2_neq_din1          (din2_neq_din1_11_9),
        .din2_gt_din1           (din2_gt_din1_11_9)
);
fpu_in2_gt_in1_3b fpu_in2_gt_in1_8_6 (
        .din1                   (din1[8:6]),
        .din2                   (din2[8:6]),
        .din2_neq_din1          (din2_neq_din1_8_6),
        .din2_gt_din1           (din2_gt_din1_8_6)
);
fpu_in2_gt_in1_3b fpu_in2_gt_in1_5_3 (
        .din1                   (din1[5:3]),
        .din2                   (din2[5:3]),
        .din2_neq_din1          (din2_neq_din1_5_3),
        .din2_gt_din1           (din2_gt_din1_5_3)
);
fpu_in2_gt_in1_3b fpu_in2_gt_in1_2_0 (
        .din1                   (din1[2:0]),
        .din2                   (din2[2:0]),
        .din2_neq_din1          (din2_neq_din1_2_0),
        .din2_gt_din1           (din2_gt_din1_2_0)
);
fpu_in2_gt_in1_3to1 fpu_in2_gt_in1_51_45 (
	.din2_neq_din1_hi	(din2_neq_din1_51_50),
	.din2_gt_din1_hi	(din2_gt_din1_51_50),
	.din2_neq_din1_mid	(din2_neq_din1_49_48),
	.din2_gt_din1_mid	(din2_gt_din1_49_48),
	.din2_neq_din1_lo	(din2_neq_din1_47_45),
	.din2_gt_din1_lo	(din2_gt_din1_47_45),
	.din2_neq_din1		(din2_neq_din1_51_45),
	.din2_gt_din1		(din2_gt_din1_51_45)
);
fpu_in2_gt_in1_3to1 fpu_in2_gt_in1_44_36 (
        .din2_neq_din1_hi       (din2_neq_din1_44_42),
        .din2_gt_din1_hi        (din2_gt_din1_44_42),
        .din2_neq_din1_mid      (din2_neq_din1_41_39),
        .din2_gt_din1_mid       (din2_gt_din1_41_39),
        .din2_neq_din1_lo       (din2_neq_din1_38_36),
        .din2_gt_din1_lo        (din2_gt_din1_38_36),
        .din2_neq_din1          (din2_neq_din1_44_36),
	.din2_gt_din1           (din2_gt_din1_44_36)
);
fpu_in2_gt_in1_3to1 fpu_in2_gt_in1_35_27 (
        .din2_neq_din1_hi       (din2_neq_din1_35_33),
        .din2_gt_din1_hi        (din2_gt_din1_35_33),
        .din2_neq_din1_mid      (din2_neq_din1_32_30),
        .din2_gt_din1_mid       (din2_gt_din1_32_30),
        .din2_neq_din1_lo       (din2_neq_din1_29_27),
        .din2_gt_din1_lo        (din2_gt_din1_29_27),
        .din2_neq_din1          (din2_neq_din1_35_27),
        .din2_gt_din1           (din2_gt_din1_35_27)
);
fpu_in2_gt_in1_3to1 fpu_in2_gt_in1_26_18 (
        .din2_neq_din1_hi       (din2_neq_din1_26_24),
        .din2_gt_din1_hi        (din2_gt_din1_26_24),
        .din2_neq_din1_mid      (din2_neq_din1_23_21),
        .din2_gt_din1_mid       (din2_gt_din1_23_21),
        .din2_neq_din1_lo       (din2_neq_din1_20_18),
        .din2_gt_din1_lo        (din2_gt_din1_20_18),
        .din2_neq_din1          (din2_neq_din1_26_18),
        .din2_gt_din1           (din2_gt_din1_26_18)
);
fpu_in2_gt_in1_3to1 fpu_in2_gt_in1_17_9 (
        .din2_neq_din1_hi       (din2_neq_din1_17_15),
        .din2_gt_din1_hi        (din2_gt_din1_17_15),
        .din2_neq_din1_mid      (din2_neq_din1_14_12),
        .din2_gt_din1_mid       (din2_gt_din1_14_12),
        .din2_neq_din1_lo       (din2_neq_din1_11_9),
        .din2_gt_din1_lo        (din2_gt_din1_11_9),
        .din2_neq_din1          (din2_neq_din1_17_9),
        .din2_gt_din1           (din2_gt_din1_17_9)
);
fpu_in2_gt_in1_3to1 fpu_in2_gt_in1_8_0 (
        .din2_neq_din1_hi       (din2_neq_din1_8_6),
        .din2_gt_din1_hi        (din2_gt_din1_8_6),
        .din2_neq_din1_mid      (din2_neq_din1_5_3),
        .din2_gt_din1_mid       (din2_gt_din1_5_3),
        .din2_neq_din1_lo       (din2_neq_din1_2_0),
        .din2_gt_din1_lo        (din2_gt_din1_2_0),
        .din2_neq_din1          (din2_neq_din1_8_0),
        .din2_gt_din1           (din2_gt_din1_8_0)
);
fpu_in2_gt_in1_3to1 fpu_in2_gt_in1_51_27 (
	.din2_neq_din1_hi       (din2_neq_din1_51_45),
	.din2_gt_din1_hi	(din2_gt_din1_51_45),
	.din2_neq_din1_mid      (din2_neq_din1_44_36),
	.din2_gt_din1_mid       (din2_gt_din1_44_36),
	.din2_neq_din1_lo       (din2_neq_din1_35_27),
	.din2_gt_din1_lo        (din2_gt_din1_35_27),
	.din2_neq_din1          (din2_neq_din1_51_27),
	.din2_gt_din1           (din2_gt_din1_51_27)
);
fpu_in2_gt_in1_3to1 fpu_in2_gt_in1_26_0 (
	.din2_neq_din1_hi       (din2_neq_din1_26_18),
	.din2_gt_din1_hi        (din2_gt_din1_26_18),
	.din2_neq_din1_mid      (din2_neq_din1_17_9),
	.din2_gt_din1_mid       (din2_gt_din1_17_9),
	.din2_neq_din1_lo       (din2_neq_din1_8_0),
	.din2_gt_din1_lo        (din2_gt_din1_8_0),
	.din2_neq_din1          (din2_neq_din1_26_0),
	.din2_gt_din1           (din2_gt_din1_26_0)
);
assign din2_neq_din1= din2_neq_din1_51_27
		|| din2_neq_din1_26_0
		|| (din2_neq_din1_54_52 && sngop);
assign din2_gt_din1= (din2_neq_din1_54_52 && din2_gt_din1_54_52
			&& sngop)
		|| ((!(din2_neq_din1_54_52 && sngop))
			&& din2_neq_din1_51_27 && din2_gt_din1_51_27)
		|| ((!(din2_neq_din1_54_52 && sngop))
			&& (!din2_neq_din1_51_27)
			&& din2_gt_din1_26_0);
assign din2_gt1_din1= expadd11
		|| (din2_gt_din1 && expeq);
endmodule
module fpu_mul (
	inq_op,
	inq_rnd_mode,
	inq_id,
	inq_in1,
	inq_in1_53_0_neq_0,
	inq_in1_50_0_neq_0,
	inq_in1_53_32_neq_0,
	inq_in1_exp_eq_0,
	inq_in1_exp_neq_ffs,
	inq_in2,
	inq_in2_53_0_neq_0,
	inq_in2_50_0_neq_0,
	inq_in2_53_32_neq_0,
	inq_in2_exp_eq_0,
	inq_in2_exp_neq_ffs,
	inq_mul,
	mul_dest_rdy,
	mul_dest_rdya,
	fmul_clken_l,
	fmul_clken_l_buf1,
	arst_l,
	grst_l,
	rclk,
	
	mul_pipe_active,
	m1stg_step,
	m6stg_fmul_in,
	m6stg_id_in,
	mul_exc_out,
	m6stg_fmul_dbl_dst,
	m6stg_fmuls,
	mul_sign_out,
	mul_exp_out,
	mul_frac_out,
	se_mul,
	se_mul64,
	si,
	so
);
input [7:0]	inq_op;			
input [1:0]	inq_rnd_mode;		
input [4:0]	inq_id;			
input [63:0]	inq_in1;		
input		inq_in1_53_0_neq_0;	
input		inq_in1_50_0_neq_0;	
input		inq_in1_53_32_neq_0;	
input		inq_in1_exp_eq_0;	
input		inq_in1_exp_neq_ffs;	
input [63:0]	inq_in2;		
input		inq_in2_53_0_neq_0;	
input		inq_in2_50_0_neq_0;	
input		inq_in2_53_32_neq_0;	
input		inq_in2_exp_eq_0;	
input		inq_in2_exp_neq_ffs;	
input		inq_mul;		
input		mul_dest_rdy;		
input		mul_dest_rdya;		
input		fmul_clken_l;           
input		fmul_clken_l_buf1;           
input		arst_l;			
input		grst_l;			
input		rclk;			
output		mul_pipe_active;        
output		m1stg_step;		
output		m6stg_fmul_in;		
output [9:0]	m6stg_id_in;		
output [4:0]	mul_exc_out;		
output		m6stg_fmul_dbl_dst;	
output		m6stg_fmuls;		
output		mul_sign_out;		
output [10:0]	mul_exp_out;		
output [51:0]	mul_frac_out;		
input           se_mul;     
input           se_mul64;       
input           si;                     
output          so;                     
wire		m1stg_snan_sng_in1;	
wire		m1stg_snan_dbl_in1;	
wire		m1stg_snan_sng_in2;	
wire		m1stg_snan_dbl_in2;	
wire		m1stg_step;		
wire		m1stg_sngop;		
wire		m1stg_dblop;		
wire		m1stg_dblop_inv;	
wire		m1stg_fmul;		
wire		m1stg_fsmuld;		
wire		m2stg_fmuls;		
wire		m2stg_fmuld;		
wire		m2stg_fsmuld;		
wire		m5stg_fmuls;		
wire		m5stg_fmuld;		
wire		m5stg_fmulda;		
wire		m6stg_fmul_in;		
wire [9:0]	m6stg_id_in;		
wire		m6stg_fmul_dbl_dst;	
wire		m6stg_fmuls;		
wire		m6stg_step;		
wire		mul_sign_out;		
wire		m5stg_in_of;		
wire [4:0]	mul_exc_out;		
wire		m2stg_frac1_dbl_norm;	
wire		m2stg_frac1_dbl_dnrm;	
wire		m2stg_frac1_sng_norm;	
wire		m2stg_frac1_sng_dnrm;	
wire		m2stg_frac1_inf;	
wire		m2stg_frac2_dbl_norm;	
wire		m2stg_frac2_dbl_dnrm;	
wire		m2stg_frac2_sng_norm;	
wire		m2stg_frac2_sng_dnrm;	
wire		m2stg_frac2_inf;	
wire		m1stg_inf_zero_in;	
wire		m1stg_inf_zero_in_dbl;	
wire		m2stg_exp_expadd;	
wire		m2stg_exp_0bff;		
wire		m2stg_exp_017f;		
wire		m2stg_exp_04ff;		
wire		m2stg_exp_zero;		
wire [6:0]	m3bstg_ld0_inv;		
wire [5:0]	m4stg_sh_cnt_in;	
wire            m4stg_inc_exp_54;       
wire            m4stg_inc_exp_55;       
wire            m4stg_inc_exp_105;      
wire		m4stg_left_shift_step;	
wire		m4stg_right_shift_step;	
wire		m5stg_to_0;		
wire		m5stg_to_0_inv;		
wire		mul_frac_out_fracadd;	
wire		mul_frac_out_frac;	
wire		mul_exp_out_exp_plus1;	
wire		mul_exp_out_exp;	
wire		mul_pipe_active;        
wire mul_rst_l; 
wire [12:0]	m3stg_exp;		
wire		m3stg_expadd_eq_0;	
wire		m3stg_expadd_lte_0_inv;	
wire [12:0]	m4stg_exp;		
wire [12:0]	m5stg_exp;		
wire [10:0]	mul_exp_out;		
wire [52:0]	m2stg_frac1_array_in;	
wire [52:0]	m2stg_frac2_array_in;	
wire [5:0]	m1stg_ld0_1;		
wire [5:0]	m1stg_ld0_2;		
wire		m4stg_frac_105;		
wire [6:0]	m3stg_ld0_inv;		
wire		m4stg_shl_54;		
wire		m4stg_shl_55;		
wire [32:0]	m5stg_frac_32_0;	
wire		m5stg_frac_dbl_nx;	
wire		m5stg_frac_sng_nx;	
wire		m5stg_frac_neq_0;	
wire		m5stg_fracadd_cout;	
wire [51:0]	mul_frac_out;		
wire [105:0]	m4stg_frac;		
wire [29:0] m4stg_frac_unused; 
wire        scan_out_fpu_mul_ctl;
wire        scan_out_fpu_mul_exp_dp;
wire        scan_out_fpu_mul_frac_dp;
fpu_mul_ctl fpu_mul_ctl (
	.inq_in1_51			(inq_in1[51]),
	.inq_in1_54			(inq_in1[54]),
	.inq_in1_53_0_neq_0		(inq_in1_53_0_neq_0),
	.inq_in1_50_0_neq_0		(inq_in1_50_0_neq_0),
	.inq_in1_53_32_neq_0		(inq_in1_53_32_neq_0),
	.inq_in1_exp_eq_0		(inq_in1_exp_eq_0),
	.inq_in1_exp_neq_ffs		(inq_in1_exp_neq_ffs),
	.inq_in2_51			(inq_in2[51]),
	.inq_in2_54			(inq_in2[54]),
	.inq_in2_53_0_neq_0		(inq_in2_53_0_neq_0),
	.inq_in2_50_0_neq_0		(inq_in2_50_0_neq_0),
	.inq_in2_53_32_neq_0		(inq_in2_53_32_neq_0),
	.inq_in2_exp_eq_0		(inq_in2_exp_eq_0),
	.inq_in2_exp_neq_ffs		(inq_in2_exp_neq_ffs),
	.inq_op				(inq_op[7:0]),
	.inq_mul			(inq_mul),
	.inq_rnd_mode			(inq_rnd_mode[1:0]),
	.inq_id				(inq_id[4:0]),
	.inq_in1_63			(inq_in1[63]),
	.inq_in2_63			(inq_in2[63]),
	.mul_dest_rdy			(mul_dest_rdy),
	.mul_dest_rdya			(mul_dest_rdya),
	.m5stg_exp			(m5stg_exp[12:0]),
	.m5stg_fracadd_cout		(m5stg_fracadd_cout),
	.m5stg_frac_neq_0		(m5stg_frac_neq_0),
	.m5stg_frac_dbl_nx		(m5stg_frac_dbl_nx),
	.m5stg_frac_sng_nx		(m5stg_frac_sng_nx),
	.m1stg_ld0_1			(m1stg_ld0_1[5:0]),
	.m1stg_ld0_2			(m1stg_ld0_2[5:0]),
	.m3stg_exp			(m3stg_exp[12:0]),
	.m3stg_expadd_eq_0		(m3stg_expadd_eq_0),
	.m3stg_expadd_lte_0_inv		(m3stg_expadd_lte_0_inv),
	.m3stg_ld0_inv			(m3stg_ld0_inv[5:0]),
	.m4stg_exp			(m4stg_exp[12:0]),
	.m4stg_frac_105			(m4stg_frac_105),
	.m5stg_frac			(m5stg_frac_32_0[32:0]),
	.arst_l				(arst_l),
	.grst_l				(grst_l),
	.mula_rst_l    (mul_rst_l),
	.rclk			(rclk),
	.mul_pipe_active                (mul_pipe_active),
	.m1stg_snan_sng_in1		(m1stg_snan_sng_in1),
	.m1stg_snan_dbl_in1		(m1stg_snan_dbl_in1),
	.m1stg_snan_sng_in2		(m1stg_snan_sng_in2),
	.m1stg_snan_dbl_in2		(m1stg_snan_dbl_in2),
	.m1stg_step			(m1stg_step),
	.m1stg_sngop			(m1stg_sngop),
	.m1stg_dblop			(m1stg_dblop),
	.m1stg_dblop_inv		(m1stg_dblop_inv),
	.m1stg_fmul			(m1stg_fmul),
	.m1stg_fsmuld			(m1stg_fsmuld),
	.m2stg_fmuls			(m2stg_fmuls),
	.m2stg_fmuld			(m2stg_fmuld),
	.m2stg_fsmuld			(m2stg_fsmuld),
	.m5stg_fmuls			(m5stg_fmuls),
	.m5stg_fmuld			(m5stg_fmuld),
	.m5stg_fmulda			(m5stg_fmulda),
	.m6stg_fmul_in			(m6stg_fmul_in),
	.m6stg_id_in			(m6stg_id_in[9:0]),
	.m6stg_fmul_dbl_dst		(m6stg_fmul_dbl_dst),
	.m6stg_fmuls			(m6stg_fmuls),
	.m6stg_step			(m6stg_step),
	.mul_sign_out			(mul_sign_out),
	.m5stg_in_of			(m5stg_in_of),
	.mul_exc_out			(mul_exc_out[4:0]),
	.m2stg_frac1_dbl_norm		(m2stg_frac1_dbl_norm),
	.m2stg_frac1_dbl_dnrm		(m2stg_frac1_dbl_dnrm),
	.m2stg_frac1_sng_norm		(m2stg_frac1_sng_norm),
	.m2stg_frac1_sng_dnrm		(m2stg_frac1_sng_dnrm),
	.m2stg_frac1_inf		(m2stg_frac1_inf),
	.m2stg_frac2_dbl_norm		(m2stg_frac2_dbl_norm),
	.m2stg_frac2_dbl_dnrm		(m2stg_frac2_dbl_dnrm),
	.m2stg_frac2_sng_norm		(m2stg_frac2_sng_norm),
	.m2stg_frac2_sng_dnrm		(m2stg_frac2_sng_dnrm),
	.m2stg_frac2_inf		(m2stg_frac2_inf),
	.m1stg_inf_zero_in		(m1stg_inf_zero_in),
	.m1stg_inf_zero_in_dbl		(m1stg_inf_zero_in_dbl),
	.m2stg_exp_expadd		(m2stg_exp_expadd),
	.m2stg_exp_0bff			(m2stg_exp_0bff),
	.m2stg_exp_017f			(m2stg_exp_017f),
	.m2stg_exp_04ff			(m2stg_exp_04ff),
	.m2stg_exp_zero			(m2stg_exp_zero),
	.m3bstg_ld0_inv			(m3bstg_ld0_inv[6:0]),
	.m4stg_sh_cnt_in		(m4stg_sh_cnt_in[5:0]),
	.m4stg_inc_exp_54		(m4stg_inc_exp_54),
	.m4stg_inc_exp_55		(m4stg_inc_exp_55),
	.m4stg_inc_exp_105		(m4stg_inc_exp_105),
	.m4stg_left_shift_step		(m4stg_left_shift_step),
	.m4stg_right_shift_step		(m4stg_right_shift_step),
	.m5stg_to_0			(m5stg_to_0),
	.m5stg_to_0_inv			(m5stg_to_0_inv),
	.mul_frac_out_fracadd		(mul_frac_out_fracadd),
	.mul_frac_out_frac		(mul_frac_out_frac),
	.mul_exp_out_exp_plus1		(mul_exp_out_exp_plus1),
	.mul_exp_out_exp		(mul_exp_out_exp),
	.se                             (se_mul),
        .si                             (si),
        .so                             (scan_out_fpu_mul_ctl)
);
fpu_mul_exp_dp fpu_mul_exp_dp (
	.inq_in1			(inq_in1[62:52]),
	.inq_in2			(inq_in2[62:52]),
	.m6stg_step			(m6stg_step),
	.m1stg_dblop			(m1stg_dblop),
	.m1stg_sngop			(m1stg_sngop),
	.m2stg_exp_expadd		(m2stg_exp_expadd),
	.m2stg_exp_0bff			(m2stg_exp_0bff),
	.m2stg_exp_017f			(m2stg_exp_017f),
	.m2stg_exp_04ff			(m2stg_exp_04ff),
	.m2stg_exp_zero			(m2stg_exp_zero),
	.m1stg_fsmuld			(m1stg_fsmuld),
	.m2stg_fmuld			(m2stg_fmuld),
	.m2stg_fmuls			(m2stg_fmuls),
	.m2stg_fsmuld			(m2stg_fsmuld),
	.m3stg_ld0_inv			(m3stg_ld0_inv[6:0]),
	.m4stg_inc_exp_54		(m4stg_inc_exp_54),
	.m4stg_inc_exp_55		(m4stg_inc_exp_55),
	.m4stg_inc_exp_105		(m4stg_inc_exp_105),
	.m5stg_fracadd_cout		(m5stg_fracadd_cout),
	.mul_exp_out_exp_plus1		(mul_exp_out_exp_plus1),
	.mul_exp_out_exp		(mul_exp_out_exp),
	.m5stg_in_of			(m5stg_in_of),
	.m5stg_fmuld			(m5stg_fmuld),
	.m5stg_to_0_inv			(m5stg_to_0_inv),
	.m4stg_shl_54			(m4stg_shl_54),
	.m4stg_shl_55			(m4stg_shl_55),
	.fmul_clken_l			(fmul_clken_l_buf1),
	.rclk			(rclk),
	.m3stg_exp			(m3stg_exp[12:0]),
	.m3stg_expadd_eq_0		(m3stg_expadd_eq_0),
	.m3stg_expadd_lte_0_inv		(m3stg_expadd_lte_0_inv),
	.m4stg_exp			(m4stg_exp[12:0]),
	.m5stg_exp			(m5stg_exp[12:0]),
	.mul_exp_out			(mul_exp_out[10:0]),
	.se                             (se_mul),
        .si                             (scan_out_fpu_mul_ctl),
        .so                             (scan_out_fpu_mul_exp_dp)
);
fpu_mul_frac_dp fpu_mul_frac_dp (
	.inq_in1			(inq_in1[54:0]),
	.inq_in2			(inq_in2[54:0]),
	.m6stg_step			(m6stg_step),
	.m2stg_frac1_dbl_norm		(m2stg_frac1_dbl_norm),
	.m2stg_frac1_dbl_dnrm		(m2stg_frac1_dbl_dnrm),
	.m2stg_frac1_sng_norm		(m2stg_frac1_sng_norm),
	.m2stg_frac1_sng_dnrm		(m2stg_frac1_sng_dnrm),
	.m2stg_frac1_inf		(m2stg_frac1_inf),
	.m1stg_snan_dbl_in1		(m1stg_snan_dbl_in1),
	.m1stg_snan_sng_in1		(m1stg_snan_sng_in1),
	.m2stg_frac2_dbl_norm		(m2stg_frac2_dbl_norm),
	.m2stg_frac2_dbl_dnrm		(m2stg_frac2_dbl_dnrm),
	.m2stg_frac2_sng_norm		(m2stg_frac2_sng_norm),
	.m2stg_frac2_sng_dnrm		(m2stg_frac2_sng_dnrm),
	.m2stg_frac2_inf		(m2stg_frac2_inf),
	.m1stg_snan_dbl_in2		(m1stg_snan_dbl_in2),
	.m1stg_snan_sng_in2		(m1stg_snan_sng_in2),
	.m1stg_inf_zero_in		(m1stg_inf_zero_in),
	.m1stg_inf_zero_in_dbl		(m1stg_inf_zero_in_dbl),
	.m1stg_dblop			(m1stg_dblop),
	.m1stg_dblop_inv		(m1stg_dblop_inv),
	.m4stg_frac			(m4stg_frac),
	.m4stg_sh_cnt_in		(m4stg_sh_cnt_in[5:0]),
	.m3bstg_ld0_inv			(m3bstg_ld0_inv[6:0]),
	.m4stg_left_shift_step		(m4stg_left_shift_step),
	.m4stg_right_shift_step		(m4stg_right_shift_step),
	.m5stg_fmuls			(m5stg_fmuls),
	.m5stg_fmulda			(m5stg_fmulda),
	.mul_frac_out_fracadd		(mul_frac_out_fracadd),
	.mul_frac_out_frac		(mul_frac_out_frac),
	.m5stg_in_of			(m5stg_in_of),
	.m5stg_to_0			(m5stg_to_0),
	.fmul_clken_l			(fmul_clken_l),
	.rclk			(rclk),
	.m2stg_frac1_array_in		(m2stg_frac1_array_in),
	.m2stg_frac2_array_in		(m2stg_frac2_array_in),
	.m1stg_ld0_1			(m1stg_ld0_1),
	.m1stg_ld0_2			(m1stg_ld0_2),
	.m4stg_frac_105			(m4stg_frac_105),
	.m3stg_ld0_inv			(m3stg_ld0_inv[6:0]),
	.m4stg_shl_54			(m4stg_shl_54),
	.m4stg_shl_55			(m4stg_shl_55),
	.m5stg_frac_32_0		(m5stg_frac_32_0[32:0]),
	.m5stg_frac_dbl_nx		(m5stg_frac_dbl_nx),
	.m5stg_frac_sng_nx		(m5stg_frac_sng_nx),
	.m5stg_frac_neq_0		(m5stg_frac_neq_0),
	.m5stg_fracadd_cout		(m5stg_fracadd_cout),
	.mul_frac_out			(mul_frac_out[51:0]),
	.se                             (se_mul),
        .si                             (scan_out_fpu_mul_exp_dp),
        .so                             (scan_out_fpu_mul_frac_dp)
);
mul64 i_m4stg_frac (
	.rs1_l ({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
		1'b1, 1'b1, 1'b1, m2stg_frac1_array_in[52:0]}),
	.rs2 ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, m2stg_frac2_array_in[52:0]}),
	.valid(m1stg_fmul),
	.areg ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0}),
	.accreg ({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
	.x2 (1'b0),
	.rclk (rclk),
	.si (scan_out_fpu_mul_frac_dp),
	.se (se_mul64),
	.mul_rst_l (mul_rst_l),
	.mul_step (m6stg_step),
	.so (so),
	.out ({m4stg_frac_unused[29:0], m4stg_frac[105:0]})
);
endmodule
module fpu_mul_ctl (
	inq_in1_51,
	inq_in1_54,
	inq_in1_53_0_neq_0,
	inq_in1_50_0_neq_0,
	inq_in1_53_32_neq_0,
	inq_in1_exp_eq_0,
	inq_in1_exp_neq_ffs,
	inq_in2_51,
	inq_in2_54,
	inq_in2_53_0_neq_0,
	inq_in2_50_0_neq_0,
	inq_in2_53_32_neq_0,
	inq_in2_exp_eq_0,
	inq_in2_exp_neq_ffs,
	inq_op,
	inq_mul,
	inq_rnd_mode,
	inq_id,
	inq_in1_63,
	inq_in2_63,
	mul_dest_rdy,
	mul_dest_rdya,
	m5stg_exp,
	m5stg_fracadd_cout,
	m5stg_frac_neq_0,
	m5stg_frac_dbl_nx,
	m5stg_frac_sng_nx,
	m1stg_ld0_1,
	m1stg_ld0_2,
	m3stg_exp,
	m3stg_expadd_eq_0,
	m3stg_expadd_lte_0_inv,
	m3stg_ld0_inv,
	m4stg_exp,
	m4stg_frac_105,
	m5stg_frac,
	arst_l,
	grst_l,
	rclk,
	mul_pipe_active,
	m1stg_snan_sng_in1,
	m1stg_snan_dbl_in1,
	m1stg_snan_sng_in2,
	m1stg_snan_dbl_in2,
	m1stg_step,
	m1stg_sngop,
	m1stg_dblop,
	m1stg_dblop_inv,
	m1stg_fmul,
	m1stg_fsmuld,
	m2stg_fmuls,
	m2stg_fmuld,
	m2stg_fsmuld,
	m5stg_fmuls,
	m5stg_fmuld,
	m5stg_fmulda,
	m6stg_fmul_in,
	m6stg_id_in,
	m6stg_fmul_dbl_dst,
	m6stg_fmuls,
	m6stg_step,
	mul_sign_out,
	m5stg_in_of,
	mul_exc_out,
	m2stg_frac1_dbl_norm,
	m2stg_frac1_dbl_dnrm,
	m2stg_frac1_sng_norm,
	m2stg_frac1_sng_dnrm,
	m2stg_frac1_inf,
	m2stg_frac2_dbl_norm,
	m2stg_frac2_dbl_dnrm,
	m2stg_frac2_sng_norm,
	m2stg_frac2_sng_dnrm,
	m2stg_frac2_inf,
	m1stg_inf_zero_in,
	m1stg_inf_zero_in_dbl,
	m2stg_exp_expadd,
	m2stg_exp_0bff,
	m2stg_exp_017f,
	m2stg_exp_04ff,
	m2stg_exp_zero,
	m3bstg_ld0_inv,
	m4stg_sh_cnt_in,
	m4stg_inc_exp_54,
	m4stg_inc_exp_55,
	m4stg_inc_exp_105,
	m4stg_left_shift_step,
	m4stg_right_shift_step,
	m5stg_to_0,
	m5stg_to_0_inv,
	mul_frac_out_fracadd,
	mul_frac_out_frac,
	mul_exp_out_exp_plus1,
	mul_exp_out_exp,
	mula_rst_l,
	se,
	si,
	so
);
parameter
		FMULS=  8'h49,
		FMULD=	8'h4a,
		FSMULD=	8'h69;
input		inq_in1_51;		
input		inq_in1_54;		
input		inq_in1_53_0_neq_0;	
input		inq_in1_50_0_neq_0;	
input		inq_in1_53_32_neq_0;	
input		inq_in1_exp_eq_0;	
input		inq_in1_exp_neq_ffs;	
input		inq_in2_51;		
input		inq_in2_54;		
input		inq_in2_53_0_neq_0;	
input		inq_in2_50_0_neq_0;	
input		inq_in2_53_32_neq_0;	
input		inq_in2_exp_eq_0;	
input		inq_in2_exp_neq_ffs;	
input [7:0]	inq_op;			
input		inq_mul;		
input [1:0]	inq_rnd_mode;		
input [4:0]	inq_id;			
input		inq_in1_63;		
input		inq_in2_63;		
input		mul_dest_rdy;		
input		mul_dest_rdya;		
input [12:0]	m5stg_exp;		
input		m5stg_fracadd_cout;	
input		m5stg_frac_neq_0;	
input		m5stg_frac_dbl_nx;	
input		m5stg_frac_sng_nx;	
input [5:0]	m1stg_ld0_1;		
input [5:0]	m1stg_ld0_2;		
input [12:0]	m3stg_exp;		
input		m3stg_expadd_eq_0;	
input		m3stg_expadd_lte_0_inv;	
input [5:0]	m3stg_ld0_inv;		
input [12:0]	m4stg_exp;		
input		m4stg_frac_105;	
input [32:0]	m5stg_frac;		
input		arst_l;			
input		grst_l;			
input		rclk;		
output		mul_pipe_active;        
output		m1stg_snan_sng_in1;	
output		m1stg_snan_dbl_in1;	
output		m1stg_snan_sng_in2;	
output		m1stg_snan_dbl_in2;	
output		m1stg_step;		
output		m1stg_sngop;		
output		m1stg_dblop;		
output		m1stg_dblop_inv;	
output		m1stg_fmul;		
output		m1stg_fsmuld;		
output		m2stg_fmuls;		
output		m2stg_fmuld;		
output		m2stg_fsmuld;		
output		m5stg_fmuls;		
output		m5stg_fmuld;		
output		m5stg_fmulda;		
output		m6stg_fmul_in;		
output [9:0]	m6stg_id_in;		
output		m6stg_fmul_dbl_dst;	
output		m6stg_fmuls;		
output		m6stg_step;		
output		mul_sign_out;		
output		m5stg_in_of;		
output [4:0]	mul_exc_out;		
output		m2stg_frac1_dbl_norm;	
output		m2stg_frac1_dbl_dnrm;	
output		m2stg_frac1_sng_norm;	
output		m2stg_frac1_sng_dnrm;	
output		m2stg_frac1_inf;	
output		m2stg_frac2_dbl_norm;	
output		m2stg_frac2_dbl_dnrm;	
output		m2stg_frac2_sng_norm;	
output		m2stg_frac2_sng_dnrm;	
output		m2stg_frac2_inf;	
output		m1stg_inf_zero_in;	
output		m1stg_inf_zero_in_dbl;	
output		m2stg_exp_expadd;	
output		m2stg_exp_0bff;		
output		m2stg_exp_017f;		
output		m2stg_exp_04ff;		
output		m2stg_exp_zero;		
output [6:0]	m3bstg_ld0_inv;		
output [5:0]	m4stg_sh_cnt_in;	
output          m4stg_inc_exp_54;       
output          m4stg_inc_exp_55;       
output          m4stg_inc_exp_105;      
output		m4stg_left_shift_step;	
output		m4stg_right_shift_step;	
output		m5stg_to_0;		
output		m5stg_to_0_inv;		
output		mul_frac_out_fracadd;	
output		mul_frac_out_frac;	
output		mul_exp_out_exp_plus1;	
output		mul_exp_out_exp;	
output    mula_rst_l; 
input           se;                     
input           si;                     
output          so;                     
wire		reset;
wire		mul_frac_in1_51;
wire		mul_frac_in1_54;
wire		mul_frac_in1_53_0_neq_0;
wire		mul_frac_in1_50_0_neq_0;
wire		mul_frac_in1_53_32_neq_0;
wire		mul_exp_in1_exp_eq_0;
wire		mul_exp_in1_exp_neq_ffs;
wire		mul_frac_in2_51;
wire		mul_frac_in2_54;
wire		mul_frac_in2_53_0_neq_0;
wire		mul_frac_in2_50_0_neq_0;
wire		mul_frac_in2_53_32_neq_0;
wire		mul_exp_in2_exp_eq_0;
wire		mul_exp_in2_exp_neq_ffs;
wire		m1stg_denorm_sng_in1;
wire		m1stg_denorm_dbl_in1;
wire		m1stg_denorm_sng_in2;
wire		m1stg_denorm_dbl_in2;
wire		m1stg_denorm_in1;
wire		m1stg_denorm_in2;
wire		m1stg_norm_sng_in1;
wire		m1stg_norm_dbl_in1;
wire		m1stg_norm_sng_in2;
wire		m1stg_norm_dbl_in2;
wire		m1stg_snan_sng_in1;
wire		m1stg_snan_dbl_in1;
wire		m1stg_snan_sng_in2;
wire		m1stg_snan_dbl_in2;
wire		m1stg_qnan_sng_in1;
wire		m1stg_qnan_dbl_in1;
wire		m1stg_qnan_sng_in2;
wire		m1stg_qnan_dbl_in2;
wire		m1stg_snan_in1;
wire		m1stg_snan_in2;
wire		m1stg_qnan_in1;
wire		m1stg_qnan_in2;
wire		m2stg_snan_in1;
wire		m2stg_snan_in2;
wire		m2stg_qnan_in1;
wire		m2stg_qnan_in2;
wire		m1stg_nan_sng_in1;
wire		m1stg_nan_dbl_in1;
wire		m1stg_nan_sng_in2;
wire		m1stg_nan_dbl_in2;
wire		m1stg_nan_in1;
wire		m1stg_nan_in2;
wire		m2stg_nan_in2;
wire		m1stg_inf_sng_in1;
wire		m1stg_inf_dbl_in1;
wire		m1stg_inf_sng_in2;
wire		m1stg_inf_dbl_in2;
wire		m1stg_inf_in1;
wire		m1stg_inf_in2;
wire		m1stg_inf_in;
wire		m2stg_inf_in1;
wire		m2stg_inf_in2;
wire		m2stg_inf_in;
wire		m1stg_infnan_sng_in1;
wire		m1stg_infnan_dbl_in1;
wire		m1stg_infnan_sng_in2;
wire		m1stg_infnan_dbl_in2;
wire		m1stg_infnan_in1;
wire		m1stg_infnan_in2;
wire		m1stg_infnan_in;
wire		m1stg_zero_in1;
wire		m1stg_zero_in2;
wire		m1stg_zero_in;
wire		m2stg_zero_in1;
wire		m2stg_zero_in2;
wire		m2stg_zero_in;
wire		m1stg_step;
wire [7:0]	m1stg_op_in;
wire [7:0]	m1stg_op;
wire		m1stg_mul_in;
wire		m1stg_mul;
wire		m1stg_sngop;
wire [3:0]	m1stg_sngopa;
wire		m1stg_dblop;
wire [3:0]	m1stg_dblopa;
wire		m1stg_dblop_inv_in;
wire		m1stg_dblop_inv;
wire [1:0]	m1stg_rnd_mode;
wire [4:0]	m1stg_id;
wire		m1stg_fmul;
wire		m1stg_fmul_dbl_dst;
wire		m1stg_fmuls;
wire		m1stg_fmuld;
wire		m1stg_fsmuld;
wire [4:0]	m1stg_opdec;
wire [4:0]	m2stg_opdec;
wire [1:0]	m2stg_rnd_mode;
wire [4:0]	m2stg_id;
wire		m2stg_fmul;
wire		m2stg_fmuls;
wire		m2stg_fmuld;
wire		m2stg_fsmuld;
wire [4:1]	m3astg_opdec;
wire [1:0]	m3astg_rnd_mode;
wire [4:0]	m3astg_id;
wire [4:1]	m3bstg_opdec;
wire [1:0]	m3bstg_rnd_mode;
wire [4:0]	m3bstg_id;
wire [4:1]	m3stg_opdec;
wire [1:0]	m3stg_rnd_mode;
wire [4:0]	m3stg_id;
wire		m3stg_fmul;
wire [4:1]	m4stg_opdec;
wire [1:0]	m4stg_rnd_mode;
wire [4:0]	m4stg_id;
wire		m4stg_fmul;
wire		m4stg_fmuld;
wire [4:1]	m5stg_opdec;
wire [1:0]	m5stg_rnd_mode;
wire [4:0]	m5stg_id;
wire		m5stg_fmul;
wire		m5stg_fmuls;
wire		m5stg_fmuld;
wire		m5stg_fmulda;
wire		m6stg_fmul_in;
wire [4:2]	m6stg_opdec;
wire [9:0]	m6stg_id_in;
wire [9:0]	m6stg_id;
wire		m6stg_fmul;
wire		m6stg_fmul_dbl_dst;
wire		m6stg_fmuls;
wire		m6stg_hold;
wire		m6stg_holda;
wire		m6stg_step;
wire		m6stg_stepa;
wire		m1stg_sign1;
wire		m1stg_sign2;
wire		m2stg_sign1;
wire		m2stg_sign2;
wire		m1stg_of_mask;
wire		m2stg_of_mask;
wire		m2stg_sign;
wire		m3astg_sign;
wire		m2stg_nv;
wire		m3astg_nv;
wire		m3astg_of_mask;
wire		m3bstg_sign;
wire		m3bstg_nv;
wire		m3stg_sign;
wire		m3stg_nv;
wire		m3stg_of_mask;
wire		m4stg_sign;
wire		m4stg_nv;
wire		m4stg_of_mask;
wire		m5stg_sign;
wire		m5stg_nv;
wire		m5stg_of_mask;
wire		mul_sign_out;
wire		mul_nv_out;
wire		m5stg_in_of;
wire		mul_of_out_tmp1_in;
wire		mul_of_out_tmp1;
wire		mul_of_out_tmp2;
wire		mul_of_out_cout;
wire		mul_of_out;
wire		mul_uf_out_in;
wire		mul_uf_out;
wire		mul_nx_out_in;
wire		mul_nx_out;
wire [4:0]	mul_exc_out;
wire		m2stg_frac1_dbl_norm;
wire		m2stg_frac1_dbl_dnrm;
wire		m2stg_frac1_sng_norm;
wire		m2stg_frac1_sng_dnrm;
wire		m2stg_frac1_inf;
wire		m2stg_frac2_dbl_norm;
wire		m2stg_frac2_dbl_dnrm;
wire		m2stg_frac2_sng_norm;
wire		m2stg_frac2_sng_dnrm;
wire		m2stg_frac2_inf;
wire		m1stg_inf_zero_in;
wire		m1stg_inf_zero_in_dbl;
wire [5:0]	m2stg_ld0_1_in;
wire [5:0]	m2stg_ld0_1;
wire [5:0]	m2stg_ld0_2_in;
wire [5:0]	m2stg_ld0_2;
wire		m2stg_exp_expadd;
wire		m2stg_exp_0bff;
wire		m2stg_exp_017f;
wire		m2stg_exp_04ff;
wire		m2stg_exp_zero;
wire [6:0]	m2stg_ld0;
wire [6:0]	m2stg_ld0_inv;
wire [6:0]	m3astg_ld0_inv;
wire [6:0]	m3bstg_ld0_inv;
wire		m4stg_expadd_eq_0;
wire		m3stg_exp_lte_0;
wire		m4stg_right_shift_in;
wire		m4stg_right_shift;
wire [5:0]	m3stg_exp_minus1;
wire [5:0]	m3stg_exp_inv_plus2;
wire		m3stg_exp_lt_neg57;
wire [5:0]	m4stg_sh_cnt_in;
wire		m4stg_left_shift_step;
wire		m4stg_right_shift_step;
wire		m4stg_inc_exp_54;
wire		m4stg_inc_exp_55;
wire		m4stg_inc_exp_105;
wire		m5stg_rndup;
wire		m5stg_to_0;
wire		m5stg_to_0_inv;
wire		mul_frac_out_fracadd;
wire		mul_frac_out_frac;
wire		mul_exp_out_exp_plus1;
wire		mul_exp_out_exp;
wire		mul_pipe_active_in;
wire		mul_pipe_active;
wire    mula_rst_l;
wire        mul_ctl_rst_l;
wire        m3bstf_of_mask;
dffrl_async #(1)  dffrl_mul_ctl (
  .din  (grst_l),
  .clk  (rclk),
  .rst_l(arst_l),
  .q    (mul_ctl_rst_l),
	.se (se),
	.si (),
	.so ()
  );
assign reset= (!mul_ctl_rst_l);
assign mula_rst_l = mul_ctl_rst_l;
dffe_s #(1) i_mul_frac_in1_51 (
	.din	(inq_in1_51),
	.en     (m6stg_step),
        .clk    (rclk),
 
        .q      (mul_frac_in1_51),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_mul_frac_in1_54 (
	.din	(inq_in1_54),
	.en     (m6stg_step),
        .clk    (rclk),
 
        .q      (mul_frac_in1_54),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_mul_frac_in1_53_0_neq_0 (
	.din	(inq_in1_53_0_neq_0),
	.en     (m6stg_step),
        .clk    (rclk),
 
        .q      (mul_frac_in1_53_0_neq_0),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_mul_frac_in1_50_0_neq_0 (
	.din	(inq_in1_50_0_neq_0),
	.en	(m6stg_step),
	.clk	(rclk),
	.q	(mul_frac_in1_50_0_neq_0),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_mul_frac_in1_53_32_neq_0 (
	.din	(inq_in1_53_32_neq_0),
	.en	(m6stg_step),
	.clk	(rclk),
	.q	(mul_frac_in1_53_32_neq_0),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_mul_exp_in1_exp_eq_0 (
        .din	(inq_in1_exp_eq_0),
        .en	(m6stg_step),
        .clk	(rclk),
 
        .q	(mul_exp_in1_exp_eq_0),
 
        .se	(se),
        .si	(),
        .so	()
);
dffe_s #(1) i_mul_exp_in1_exp_neq_ffs (
	.din	(inq_in1_exp_neq_ffs),
	.en	(m6stg_step),
	.clk	(rclk),
	.q	(mul_exp_in1_exp_neq_ffs),
   	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_mul_frac_in2_51 (
	.din	(inq_in2_51),
	.en	(m6stg_step),
	.clk	(rclk),
	.q	(mul_frac_in2_51),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_mul_frac_in2_54 (
	.din	(inq_in2_54),
	.en	(m6stg_step),
	.clk	(rclk),
	.q	(mul_frac_in2_54),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_mul_frac_in2_53_0_neq_0 (
	.din	(inq_in2_53_0_neq_0),
	.en  	(m6stg_step),
	.clk	(rclk),
	.q	(mul_frac_in2_53_0_neq_0),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_mul_frac_in2_50_0_neq_0 (
	.din	(inq_in2_50_0_neq_0),
	.en	(m6stg_step),
	.clk	(rclk),
	.q	(mul_frac_in2_50_0_neq_0),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_mul_frac_in2_53_32_neq_0 (
	.din	(inq_in2_53_32_neq_0),
	.en	(m6stg_step),
	.clk	(rclk),
	.q	(mul_frac_in2_53_32_neq_0),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_mul_exp_in2_exp_eq_0 (
	.din	(inq_in2_exp_eq_0),
	 .en	(m6stg_step),
	.clk	(rclk),
	.q	(mul_exp_in2_exp_eq_0),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_mul_exp_in2_exp_neq_ffs (
        .din	(inq_in2_exp_neq_ffs),
        .en	(m6stg_step),
        .clk	(rclk),
 
        .q	(mul_exp_in2_exp_neq_ffs),
 
        .se	(se),
        .si	(),
        .so	()
);
assign m1stg_denorm_sng_in1= mul_exp_in1_exp_eq_0 && m1stg_sngopa[0];
assign m1stg_denorm_dbl_in1= mul_exp_in1_exp_eq_0 && m1stg_dblopa[0];
assign m1stg_denorm_sng_in2= mul_exp_in2_exp_eq_0 && m1stg_sngopa[0];
assign m1stg_denorm_dbl_in2= mul_exp_in2_exp_eq_0 && m1stg_dblopa[0];
assign m1stg_denorm_in1= m1stg_denorm_sng_in1 || m1stg_denorm_dbl_in1;
assign m1stg_denorm_in2= m1stg_denorm_sng_in2 || m1stg_denorm_dbl_in2;
assign m1stg_norm_sng_in1= (!mul_exp_in1_exp_eq_0) && m1stg_sngopa[0];
assign m1stg_norm_dbl_in1= (!mul_exp_in1_exp_eq_0) && m1stg_dblopa[0];
assign m1stg_norm_sng_in2= (!mul_exp_in2_exp_eq_0) && m1stg_sngopa[0];
assign m1stg_norm_dbl_in2= (!mul_exp_in2_exp_eq_0) && m1stg_dblopa[0];
assign m1stg_snan_sng_in1= (!mul_exp_in1_exp_neq_ffs) && (!mul_frac_in1_54)
		&& (mul_frac_in1_53_32_neq_0) && m1stg_sngopa[1];
assign m1stg_snan_dbl_in1= (!mul_exp_in1_exp_neq_ffs)
		&& (!mul_frac_in1_51) && mul_frac_in1_50_0_neq_0
		&& m1stg_dblopa[1];
assign m1stg_snan_sng_in2= (!mul_exp_in2_exp_neq_ffs) && (!mul_frac_in2_54)
                && (mul_frac_in2_53_32_neq_0) && m1stg_sngopa[1];
assign m1stg_snan_dbl_in2= (!mul_exp_in2_exp_neq_ffs)
                && (!mul_frac_in2_51) && mul_frac_in2_50_0_neq_0
                && m1stg_dblopa[1];
assign m1stg_qnan_sng_in1= (!mul_exp_in1_exp_neq_ffs) && mul_frac_in1_54
		&& m1stg_sngopa[1];
assign m1stg_qnan_dbl_in1= (!mul_exp_in1_exp_neq_ffs) && mul_frac_in1_51
		&& m1stg_dblopa[1];
assign m1stg_qnan_sng_in2= (!mul_exp_in2_exp_neq_ffs) && mul_frac_in2_54
                && m1stg_sngopa[1];
assign m1stg_qnan_dbl_in2= (!mul_exp_in2_exp_neq_ffs) && mul_frac_in2_51
                && m1stg_dblopa[1];
assign m1stg_snan_in1= m1stg_snan_sng_in1 || m1stg_snan_dbl_in1;
assign m1stg_snan_in2= m1stg_snan_sng_in2 || m1stg_snan_dbl_in2;
assign m1stg_qnan_in1= m1stg_qnan_sng_in1 || m1stg_qnan_dbl_in1;
 
assign m1stg_qnan_in2= m1stg_qnan_sng_in2 || m1stg_qnan_dbl_in2;
dffe_s #(1) i_m2stg_snan_in1 (
	.din	(m1stg_snan_in1),
	.en	(m6stg_step),
	.clk	(rclk),
	.q	(m2stg_snan_in1),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_m2stg_snan_in2 (
	.din	(m1stg_snan_in2),
	.en	(m6stg_step),
	.clk	(rclk),
	.q	(m2stg_snan_in2),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_m2stg_qnan_in1 (
	.din	(m1stg_qnan_in1),
	.en	(m6stg_step),
	.clk	(rclk),
	.q	(m2stg_qnan_in1),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_m2stg_qnan_in2 (
	.din	(m1stg_qnan_in2),
	.en	(m6stg_step),
	.clk	(rclk),
	.q	(m2stg_qnan_in2),
	.se	(se),
	.si	(),
	.so	()
);
assign m1stg_nan_sng_in1= (!mul_exp_in1_exp_neq_ffs)
		&& (mul_frac_in1_54 || mul_frac_in1_53_32_neq_0)
		&& m1stg_sngopa[2];
assign m1stg_nan_dbl_in1= (!mul_exp_in1_exp_neq_ffs)
		&& (mul_frac_in1_51 || mul_frac_in1_50_0_neq_0)
		&& m1stg_dblopa[2];
assign m1stg_nan_sng_in2= (!mul_exp_in2_exp_neq_ffs)
		&& (mul_frac_in2_54 || mul_frac_in2_53_32_neq_0)
		&& m1stg_sngopa[2];
assign m1stg_nan_dbl_in2= (!mul_exp_in2_exp_neq_ffs)
		&& (mul_frac_in2_51 || mul_frac_in2_50_0_neq_0)
		&& m1stg_dblopa[2];
assign m1stg_nan_in1= m1stg_nan_sng_in1 || m1stg_nan_dbl_in1;
assign m1stg_nan_in2= m1stg_nan_sng_in2 || m1stg_nan_dbl_in2;
dffe_s #(1) i_m2stg_nan_in2 (
	.din	(m1stg_nan_in2),
	.en	(m6stg_step),
	.clk	(rclk),
	.q	(m2stg_nan_in2),
	.se	(se),
	.si	(),
	.so	()
);
assign m1stg_inf_sng_in1= (!mul_exp_in1_exp_neq_ffs)
		&& (!mul_frac_in1_54) && (!mul_frac_in1_53_32_neq_0)
		&& m1stg_sngopa[2];
assign m1stg_inf_dbl_in1= (!mul_exp_in1_exp_neq_ffs)
		&& (!mul_frac_in1_51) && (!mul_frac_in1_50_0_neq_0)
		&& m1stg_dblopa[2];
assign m1stg_inf_sng_in2= (!mul_exp_in2_exp_neq_ffs)
		&& (!mul_frac_in2_54) && (!mul_frac_in2_53_32_neq_0)
		&& m1stg_sngopa[2];
assign m1stg_inf_dbl_in2= (!mul_exp_in2_exp_neq_ffs)
		&& (!mul_frac_in2_51) && (!mul_frac_in2_50_0_neq_0)
		&& m1stg_dblopa[2];
assign m1stg_inf_in1= m1stg_inf_sng_in1 || m1stg_inf_dbl_in1;
assign m1stg_inf_in2= m1stg_inf_sng_in2 || m1stg_inf_dbl_in2;
assign m1stg_inf_in= m1stg_inf_in1 || m1stg_inf_in2;
dffe_s #(1) i_m2stg_inf_in1 (
	.din	(m1stg_inf_in1),
	.en	(m6stg_step),
	.clk	(rclk),
	.q	(m2stg_inf_in1),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_m2stg_inf_in2 (
	.din	(m1stg_inf_in2),
	.en	(m6stg_step),
	.clk	(rclk),
	.q	(m2stg_inf_in2),
 
        .se	(se),
        .si	(),
        .so	()
);
dffe_s #(1) i_m2stg_inf_in (
	.din	(m1stg_inf_in),
	.en	(m6stg_step),
	.clk	(rclk),
	.q	(m2stg_inf_in),
 
        .se	(se),
        .si	(),
        .so	()
);
assign m1stg_infnan_sng_in1= (!mul_exp_in1_exp_neq_ffs) && m1stg_sngopa[3];
assign m1stg_infnan_dbl_in1= (!mul_exp_in1_exp_neq_ffs) && m1stg_dblopa[3];
assign m1stg_infnan_sng_in2= (!mul_exp_in2_exp_neq_ffs) && m1stg_sngopa[3];
assign m1stg_infnan_dbl_in2= (!mul_exp_in2_exp_neq_ffs) && m1stg_dblopa[3];
assign m1stg_infnan_in1= m1stg_infnan_sng_in1 || m1stg_infnan_dbl_in1;
assign m1stg_infnan_in2= m1stg_infnan_sng_in2 || m1stg_infnan_dbl_in2;
assign m1stg_infnan_in= m1stg_infnan_in1 || m1stg_infnan_in2;
assign m1stg_zero_in1= mul_exp_in1_exp_eq_0
		&& (!mul_frac_in1_53_0_neq_0) && (!mul_frac_in1_54);
assign m1stg_zero_in2= mul_exp_in2_exp_eq_0
                && (!mul_frac_in2_53_0_neq_0) && (!mul_frac_in2_54);
assign m1stg_zero_in= m1stg_zero_in1 || m1stg_zero_in2;
dffe_s #(1) i_m2stg_zero_in1 (
	.din	(m1stg_zero_in1),
	.en	(m6stg_step),
	.clk	(rclk),
	.q	(m2stg_zero_in1),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_m2stg_zero_in2 (
	.din	(m1stg_zero_in2),
	.en	(m6stg_step),
	.clk	(rclk),
	.q	(m2stg_zero_in2),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_m2stg_zero_in (
	.din	(m1stg_zero_in),
	.en	(m6stg_step),
	.clk	(rclk),
	.q	(m2stg_zero_in),
 
        .se	(se),
        .si	(),
        .so	()
);
 
assign m1stg_step= m6stg_stepa && (!m1stg_mul);
assign m1stg_op_in[7:0]= ({8{(m1stg_step && (!reset))}}
			    & (inq_op[7:0] & {8{inq_mul}}))
		| ({8{((!m6stg_step) && (!reset))}}
			    & m1stg_op[7:0]);
dff_s #(8) i_m1stg_op (
	.din	(m1stg_op_in[7:0]),
	.clk	(rclk),
	.q	(m1stg_op[7:0]),
	.se	(se),
	.si	(),
	.so	()
);
assign m1stg_mul_in= (m1stg_step && (!reset) && inq_mul)
		|| ((!m6stg_step) && (!reset) && m1stg_mul);
dff_s #(1) i_m1stg_mul (
        .din    (m1stg_mul_in),
	.clk    (rclk),
 
        .q      (m1stg_mul),
 
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_m1stg_sngop (
	.din	(inq_op[0]),
	.en	(m6stg_step),
	.clk	(rclk),
	.q	(m1stg_sngop),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(4) i_m1stg_sngopa (
	.din	({4{inq_op[0]}}),
	.en	(m6stg_step),
        .clk	(rclk),
 
        .q	(m1stg_sngopa[3:0]),
 
        .se	(se),
        .si	(),
        .so	()
);
dffe_s #(1) i_m1stg_dblop (
        .din    (inq_op[1]),
        .en     (m6stg_step),
        .clk    (rclk),
 
        .q      (m1stg_dblop),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(4) i_m1stg_dblopa (
	.din	({4{inq_op[1]}}),
	.en	(m6stg_step),
	.clk	(rclk),
	 .q	(m1stg_dblopa[3:0]),
	.se	(se),
	.si	(),
	.so	()
);
assign m1stg_dblop_inv_in= (!inq_op[1]);
dffe_s #(1) i_m1stg_dblop_inv (
        .din	(m1stg_dblop_inv_in),
        .en	(m6stg_step),
        .clk	(rclk),
 
        .q	(m1stg_dblop_inv),
 
        .se	(se),
        .si	(),
        .so	()
);
dffe_s #(2) i_m1stg_rnd_mode (
	.din	(inq_rnd_mode[1:0]),
	.en	(m6stg_step),
	.clk    (rclk),
        .q      (m1stg_rnd_mode[1:0]),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(5) i_m1stg_id (
	.din	(inq_id[4:0]),
	.en     (m6stg_step),
        .clk    (rclk),
 
        .q      (m1stg_id[4:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign m1stg_fmul= (m1stg_op[7:0]==FMULS) || (m1stg_op[7:0]==FMULD)
		|| (m1stg_op[7:0]==FSMULD);
assign m1stg_fmul_dbl_dst= (m1stg_op[7:0]==FMULD) || (m1stg_op[7:0]==FSMULD);
assign m1stg_fmuls= (m1stg_op[7:0]==FMULS);
assign m1stg_fmuld= (m1stg_op[7:0]==FMULD);
assign m1stg_fsmuld= (m1stg_op[7:0]==FSMULD);
assign m1stg_opdec[4:0]= {m1stg_fmul,
			m1stg_fmul_dbl_dst,
			m1stg_fmuls,
			m1stg_fmuld,
			m1stg_fsmuld};
dffre_s #(5) i_m2stg_opdec (
	.din	(m1stg_opdec[4:0]),
	.en	(m6stg_step),
	.rst	(reset),
	.clk	(rclk),
	.q	(m2stg_opdec[4:0]),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(2) i_m2stg_rnd_mode (
        .din    (m1stg_rnd_mode[1:0]),
        .en     (m6stg_step),
        .clk    (rclk),
 
        .q      (m2stg_rnd_mode[1:0]),
        .se     (se),
        .si     (),
        .so     ()
);
 
dffe_s #(5) i_m2stg_id (
        .din    (m1stg_id[4:0]),
        .en     (m6stg_step),
        .clk    (rclk),
 
        .q      (m2stg_id[4:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign m2stg_fmul= m2stg_opdec[4];
assign m2stg_fmuls= m2stg_opdec[2];
assign m2stg_fmuld= m2stg_opdec[1];
assign m2stg_fsmuld= m2stg_opdec[0];
dffre_s #(4) i_m3astg_opdec (
        .din    (m2stg_opdec[4:1]),
        .en     (m6stg_step),
        .rst    (reset),
        .clk    (rclk),
        .q      (m3astg_opdec[4:1]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(2) i_m3astg_rnd_mode (
        .din    (m2stg_rnd_mode[1:0]),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m3astg_rnd_mode[1:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(5) i_m3astg_id (
        .din    (m2stg_id[4:0]),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m3astg_id[4:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(4) i_m3bstg_opdec (
        .din    (m3astg_opdec[4:1]),
        .en     (m6stg_step),
        .rst    (reset),
        .clk    (rclk),
        .q      (m3bstg_opdec[4:1]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(2) i_m3bstg_rnd_mode (
        .din    (m3astg_rnd_mode[1:0]),
        .en     (m6stg_step),
        .clk    (rclk),
 
        .q      (m3bstg_rnd_mode[1:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(5) i_m3bstg_id (
        .din    (m3astg_id[4:0]),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m3bstg_id[4:0]),
 
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(4) i_m3stg_opdec (
        .din    (m3bstg_opdec[4:1]),
        .en     (m6stg_step),
        .rst    (reset),
        .clk    (rclk),
        .q      (m3stg_opdec[4:1]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(2) i_m3stg_rnd_mode (
        .din    (m3bstg_rnd_mode[1:0]),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m3stg_rnd_mode[1:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(5) i_m3stg_id (
        .din    (m3bstg_id[4:0]),
        .en     (m6stg_step),
        .clk    (rclk),
 
        .q      (m3stg_id[4:0]),
 
        .se     (se),
        .si     (),
        .so     ()
);
assign m3stg_fmul= m3stg_opdec[4];
dffre_s #(4) i_m4stg_opdec (
        .din    (m3stg_opdec[4:1]),
        .en     (m6stg_step),
        .rst    (reset),
        .clk    (rclk),
        .q      (m4stg_opdec[4:1]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(2) i_m4stg_rnd_mode (
        .din    (m3stg_rnd_mode[1:0]),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m4stg_rnd_mode[1:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(5) i_m4stg_id (
        .din    (m3stg_id[4:0]),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m4stg_id[4:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign m4stg_fmul= m4stg_opdec[4];
assign m4stg_fmuld= m4stg_opdec[1];
dffre_s #(4) i_m5stg_opdec (
        .din    (m4stg_opdec[4:1]),
        .en     (m6stg_step),
        .rst    (reset),
        .clk    (rclk),
        .q      (m5stg_opdec[4:1]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(2) i_m5stg_rnd_mode (
        .din    (m4stg_rnd_mode[1:0]),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m5stg_rnd_mode[1:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(5) i_m5stg_id (
        .din    (m4stg_id[4:0]),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m5stg_id[4:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffre_s #(1) i_m5stg_fmulda (
	.din	(m4stg_fmuld),
	.en	(m6stg_step),
	.rst	(reset),
	.clk	(rclk),
  	.q	(m5stg_fmulda),
	.se	(se),
	.si	(),
	.so	()
);
assign m5stg_fmul= m5stg_opdec[4];
assign m5stg_fmuls= m5stg_opdec[2];
assign m5stg_fmuld= m5stg_opdec[1];
assign m6stg_fmul_in= (m6stg_stepa && (!reset)
			&& m5stg_fmul)
		|| ((!m6stg_stepa) && (!reset)
			&& m6stg_fmul);
dffre_s #(3) i_m6stg_opdec (
        .din    (m5stg_opdec[4:2]),
        .en     (m6stg_step),
        .rst    (reset),
        .clk    (rclk),
        .q      (m6stg_opdec[4:2]),
        .se     (se),
        .si     (),
        .so     ()
);
assign m6stg_id_in[9:0]= ({10{m6stg_stepa}}
			    & {(m5stg_id[4:2]==3'o7),
				(m5stg_id[4:2]==3'o6),
				(m5stg_id[4:2]==3'o5),
				(m5stg_id[4:2]==3'o4),
				(m5stg_id[4:2]==3'o3),
				(m5stg_id[4:2]==3'o2),
				(m5stg_id[4:2]==3'o1),
				(m5stg_id[4:2]==3'o0),
				m5stg_id[1:0]})
		| ({10{(!m6stg_stepa)}}
			    & m6stg_id[9:0]);
dffe_s #(10) i_m6stg_id (
        .din    (m6stg_id_in[9:0]),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m6stg_id[9:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign m6stg_fmul= m6stg_opdec[4];
assign m6stg_fmul_dbl_dst= m6stg_opdec[3];
assign m6stg_fmuls= m6stg_opdec[2];
assign m6stg_hold= m6stg_fmul && (!mul_dest_rdy);
assign m6stg_holda= m6stg_fmul && (!mul_dest_rdya);
assign m6stg_step= (!m6stg_hold);
assign m6stg_stepa= (!m6stg_holda);
assign mul_pipe_active_in =  
   m1stg_fmul || m2stg_fmul || m3astg_opdec[4] || m3bstg_opdec[4] ||
   m3stg_fmul || m4stg_fmul || m5stg_fmul      || m6stg_fmul;
dffre_s #(1) i_mul_pipe_active (
	.din	(mul_pipe_active_in),
	.en     (1'b1),
        .rst    (reset),
        .clk    (rclk),
        .q      (mul_pipe_active),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_m1stg_sign1 (
        .din    (inq_in1_63),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m1stg_sign1),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_m1stg_sign2 (
        .din    (inq_in2_63),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m1stg_sign2),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_m2stg_sign1 (
        .din	(m1stg_sign1),
        .en	(m6stg_step),
        .clk	(rclk),
 
        .q	(m2stg_sign1),
 
        .se	(se),
        .si	(),
        .so	()
);
 
dffe_s #(1) i_m2stg_sign2 (
        .din	(m1stg_sign2),
        .en	(m6stg_step),
        .clk	(rclk),
 
        .q	(m2stg_sign2),
 
        .se	(se),
        .si	(),
        .so	()
);
assign m1stg_of_mask= (!m1stg_infnan_in);
dffe_s #(1) i_m2stg_of_mask (
        .din    (m1stg_of_mask),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m2stg_of_mask),
 
        .se     (se),
        .si     (),
        .so     ()
);
assign m2stg_sign= ((m2stg_sign1
				&& (!m2stg_snan_in2)
				&& (!(m2stg_qnan_in2 && (!m2stg_snan_in1))))
			^ (m2stg_sign2
				&& (!(m2stg_snan_in1 && (!m2stg_snan_in2)))
				&& (!(m2stg_qnan_in1 && (!m2stg_nan_in2)))))
		&& (!(m2stg_inf_in && m2stg_zero_in));
dffe_s #(1) i_m3astg_sign (
        .din    (m2stg_sign),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m3astg_sign),
        .se     (se),
        .si     (),
        .so     ()
);
assign m2stg_nv= m2stg_snan_in1
		|| m2stg_snan_in2
		|| (m2stg_zero_in1 && m2stg_inf_in2)
		|| (m2stg_inf_in1 && m2stg_zero_in2);
dffe_s #(1) i_m3astg_nv (
        .din    (m2stg_nv),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m3astg_nv),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_m3astg_of_mask (
        .din    (m2stg_of_mask),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m3astg_of_mask),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_m3bstg_sign (
        .din    (m3astg_sign),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m3bstg_sign),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_m3bstg_nv (
        .din    (m3astg_nv),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m3bstg_nv),
        .se     (se),
        .si     (),
        .so     ()
);
wire m3bstg_of_mask;
dffe_s #(1) i_m3bstg_of_mask (
        .din    (m3astg_of_mask),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m3bstg_of_mask),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_m3stg_sign (
        .din    (m3bstg_sign),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m3stg_sign),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_m3stg_nv (
        .din    (m3bstg_nv),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m3stg_nv),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_m3stg_of_mask (
        .din    (m3bstg_of_mask),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m3stg_of_mask),
        .se     (se),
        .si     (),
        .so     ()
);
 
dffe_s #(1) i_m4stg_sign (
        .din    (m3stg_sign),
        .en     (m6stg_step),
        .clk    (rclk),
 
        .q      (m4stg_sign),
 
        .se     (se),
        .si     (),
        .so     ()
);
 
dffe_s #(1) i_m4stg_nv (
        .din    (m3stg_nv),
        .en     (m6stg_step),
        .clk    (rclk),
 
        .q      (m4stg_nv),
 
        .se     (se),
        .si     (),
        .so     ()
);
 
dffe_s #(1) i_m4stg_of_mask (
        .din    (m3stg_of_mask),
        .en     (m6stg_step),
        .clk    (rclk),
 
        .q      (m4stg_of_mask),
 
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_m5stg_sign (
        .din    (m4stg_sign),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m5stg_sign),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_m5stg_nv (
        .din    (m4stg_nv),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m5stg_nv),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_m5stg_of_mask (
        .din    (m4stg_of_mask),
        .en     (m6stg_step),
        .clk    (rclk),
 
        .q      (m5stg_of_mask),
 
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_mul_sign_out (
	.din	(m5stg_sign),
	.en     (m6stg_step),
        .clk    (rclk),
        .q      (mul_sign_out),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_mul_nv_out (
	.din	(m5stg_nv),
	.en     (m6stg_step),
        .clk    (rclk),
        .q      (mul_nv_out),
	.se     (se),
        .si     (),
        .so     ()
);
assign m5stg_in_of= ((!m5stg_exp[12])
                        && m5stg_fmuld
                        && (m5stg_exp[11] || (&m5stg_exp[10:0]))
                        && m5stg_of_mask)
                || ((!m5stg_exp[12])
                        && m5stg_fmuls
                        && ((|m5stg_exp[11:8]) || (&m5stg_exp[7:0]))
                        && m5stg_of_mask);
assign mul_of_out_tmp1_in= ((!m5stg_exp[12])
                        && m5stg_fmuld
                        && (&m5stg_exp[10:1])
                        && m5stg_rndup
                        && m5stg_of_mask)
                || ((!m5stg_exp[12])
                        && m5stg_fmuls
                        && (&m5stg_exp[7:1])
                        && m5stg_rndup
                        && m5stg_of_mask);
dffe_s #(1) i_mul_of_out_tmp1 (
        .din    (mul_of_out_tmp1_in),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (mul_of_out_tmp1),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_mul_of_out_tmp2 (
	.din	(m5stg_in_of),
	.en	(m6stg_step),
    	.clk	(rclk),
	.q	(mul_of_out_tmp2),
	.se	(se),
	.si	(),
	.so	()
);
dffe_s #(1) i_mul_of_out_cout (
	.din	(m5stg_fracadd_cout),
	.en	(m6stg_step),
    	.clk	(rclk),
	.q	(mul_of_out_cout),
	.se	(se),
	.si	(),
	.so	()
);
assign mul_of_out= mul_of_out_tmp2
		|| (mul_of_out_tmp1 && mul_of_out_cout);
assign mul_uf_out_in= (m5stg_exp[12] || (!(|m5stg_exp[11:0])))
		&& m5stg_frac_neq_0;
dffe_s #(1) i_mul_uf_out (
        .din    (mul_uf_out_in),
        .en     (m6stg_step),
        .clk    (rclk),
 
        .q      (mul_uf_out),
 
        .se     (se),
        .si     (),
        .so     ()
);
assign mul_nx_out_in= (m5stg_fmuld && m5stg_frac_dbl_nx)
		|| (m5stg_fmuls && m5stg_frac_sng_nx);
dffe_s #(1) i_mul_nx_out (
        .din    (mul_nx_out_in),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (mul_nx_out),
        .se     (se),
        .si     (),
        .so     ()
);
assign mul_exc_out[4:0] =
  {mul_nv_out,
   mul_of_out,
   mul_uf_out,
   1'b0,
   (mul_nx_out || mul_of_out)};  
 
assign m2stg_frac1_dbl_norm= m1stg_norm_dbl_in1
		&& ((!(m1stg_infnan_dbl_in1 || m1stg_infnan_dbl_in2))
			|| (m1stg_snan_dbl_in1 && (!m1stg_snan_dbl_in2))
			|| (m1stg_qnan_dbl_in1 && (!m1stg_nan_dbl_in2)));
assign m2stg_frac1_dbl_dnrm= m1stg_denorm_dbl_in1
		&& (!(m1stg_infnan_dbl_in1 || m1stg_infnan_dbl_in2));
assign m2stg_frac1_sng_norm= m1stg_norm_sng_in1
		&& ((!(m1stg_infnan_sng_in1 || m1stg_infnan_sng_in2))
                        || (m1stg_snan_sng_in1 && (!m1stg_snan_sng_in2))
                        || (m1stg_qnan_sng_in1 && (!m1stg_nan_sng_in2)));
assign m2stg_frac1_sng_dnrm= m1stg_denorm_sng_in1
		&& (!(m1stg_infnan_sng_in1 || m1stg_infnan_sng_in2));
assign m2stg_frac1_inf= (m1stg_inf_in && (!m1stg_nan_in1) && (!m1stg_nan_in2))
		|| m1stg_snan_in2
		|| (m1stg_qnan_in2 && (!m1stg_snan_in1));
assign m2stg_frac2_dbl_norm= m1stg_norm_dbl_in2
		&& ((!(m1stg_infnan_dbl_in1 || m1stg_infnan_dbl_in2))
			|| m1stg_snan_dbl_in2
			|| (m1stg_qnan_dbl_in2 && (!m1stg_snan_dbl_in1)));
assign m2stg_frac2_dbl_dnrm= m1stg_denorm_dbl_in2
		&& (!(m1stg_infnan_dbl_in1 || m1stg_infnan_dbl_in2));
assign m2stg_frac2_sng_norm= m1stg_norm_sng_in2
		&& ((!(m1stg_infnan_sng_in1 || m1stg_infnan_sng_in2))
                        || m1stg_snan_sng_in2
                        || (m1stg_qnan_sng_in2 && (!m1stg_snan_sng_in1)));
assign m2stg_frac2_sng_dnrm= m1stg_denorm_sng_in2
		&& (!(m1stg_infnan_sng_in1 || m1stg_infnan_sng_in2));
assign m2stg_frac2_inf= (m1stg_inf_in && (!m1stg_nan_in1) && (!m1stg_nan_in2))
		|| (m1stg_snan_in1 && (!m1stg_snan_in2))
		|| (m1stg_qnan_in1 && (!m1stg_nan_in2));
assign m1stg_inf_zero_in= (m1stg_inf_in1 && m1stg_zero_in2)
		|| (m1stg_zero_in1 && m1stg_inf_in2);
assign m1stg_inf_zero_in_dbl= ((m1stg_inf_in1 && m1stg_zero_in2)
			|| (m1stg_zero_in1 && m1stg_inf_in2))
		&& m1stg_fmul_dbl_dst;
assign m2stg_ld0_1_in[5:0]= ({6{(m1stg_denorm_in1 && (!m1stg_infnan_in))}}
		& m1stg_ld0_1[5:0]);
dffe_s #(6) i_m2stg_ld0_1 (
	.din	(m2stg_ld0_1_in[5:0]),
	.en	(m6stg_step),
	.clk    (rclk),
        .q      (m2stg_ld0_1[5:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign m2stg_ld0_2_in[5:0]= ({6{(m1stg_denorm_in2 && (!m1stg_infnan_in))}}
		& m1stg_ld0_2[5:0]);
dffe_s #(6) i_m2stg_ld0_2 (
        .din    (m2stg_ld0_2_in[5:0]),
        .en     (m6stg_step),
        .clk    (rclk),
 
        .q      (m2stg_ld0_2[5:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign m2stg_exp_expadd= (!m1stg_infnan_in) && (!m1stg_zero_in);
assign m2stg_exp_0bff= m1stg_fmuld && m1stg_infnan_in;
assign m2stg_exp_017f= m1stg_fmuls && m1stg_infnan_in;
assign m2stg_exp_04ff= m1stg_fsmuld && m1stg_infnan_in;
 
assign m2stg_exp_zero= m1stg_zero_in && (!m1stg_infnan_in);
assign m2stg_ld0[6:0]= {1'b0, m2stg_ld0_1[5:0]}
			+ {1'b0, m2stg_ld0_2[5:0]};
assign m2stg_ld0_inv[6:0]= (~m2stg_ld0[6:0]);
dffe_s #(7) i_m3astg_ld0_inv (
	.din	(m2stg_ld0_inv[6:0]),
	.en     (m6stg_step),
        .clk    (rclk),
        .q      (m3astg_ld0_inv[6:0]),
	.se     (se),
        .si     (),
        .so     ()
);
dffe_s #(7) i_m3bstg_ld0_inv (
        .din    (m3astg_ld0_inv[6:0]),
        .en     (m6stg_step),
        .clk    (rclk),
        .q      (m3bstg_ld0_inv[6:0]),
 
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(1) i_m4stg_expadd_eq_0 (
        .din    (m3stg_expadd_eq_0),
        .en     (m6stg_step),
        .clk    (rclk),
 
        .q      (m4stg_expadd_eq_0),
 
        .se     (se),
        .si     (),
        .so     ()
);
assign m3stg_exp_lte_0= (!(|m3stg_exp[11:0])) || m3stg_exp[12];
assign m4stg_right_shift_in= (!m3stg_expadd_lte_0_inv) && m3stg_exp_lte_0;
dffe_s #(1) i_m4stg_right_shift (
	.din	(m4stg_right_shift_in),
	.en     (m6stg_step),
        .clk    (rclk),
        .q      (m4stg_right_shift),
	.se     (se),
        .si     (),
        .so     ()
);
assign m3stg_exp_minus1[5:0]= m3stg_exp[5:0]
			+ 6'h3f;
assign m3stg_exp_inv_plus2[5:0]= (~m3stg_exp[5:0])
			+ 6'h02;
assign m3stg_exp_lt_neg57= ((!(&m3stg_exp[11:6]))
			|| (!(|m3stg_exp[5:3])))
		&& m3stg_exp[12];
assign m4stg_sh_cnt_in[5:0]= ({6{((!m3stg_expadd_lte_0_inv)
				&& (!m3stg_exp_lte_0))}}
			    & m3stg_exp_minus1[5:0])
		| ({6{((!m3stg_expadd_lte_0_inv) && m3stg_exp_lte_0
				&& m3stg_exp_lt_neg57)}}
			    & 6'h39)
		| ({6{((!m3stg_expadd_lte_0_inv) && m3stg_exp_lte_0
				&& (!m3stg_exp_lt_neg57))}}
			    & m3stg_exp_inv_plus2[5:0])
		| ({6{m3stg_expadd_lte_0_inv}}
			    & (~m3stg_ld0_inv[5:0]));
assign m4stg_left_shift_step= (!m4stg_right_shift) && m6stg_step;
assign m4stg_right_shift_step= m4stg_right_shift && m6stg_step;
assign m4stg_inc_exp_54  = (!(|m4stg_exp[12:0])) && (!m4stg_right_shift);
assign m4stg_inc_exp_55  = !m4stg_right_shift;
assign m4stg_inc_exp_105 = m4stg_expadd_eq_0 && m4stg_right_shift && m4stg_frac_105;
assign m5stg_rndup= ((((m5stg_rnd_mode[1:0]==2'b10) && (!m5stg_sign)
					&& (m5stg_frac[2:0]!=3'b0))
				|| ((m5stg_rnd_mode[1:0]==2'b11) && m5stg_sign
					&& (m5stg_frac[2:0]!=3'b0))
				|| ((m5stg_rnd_mode[1:0]==2'b00)
					&& m5stg_frac[2]
					&& ((m5stg_frac[1:0]!=2'b0)
						|| m5stg_frac[3])))
			&& m5stg_fmuld)
		|| ((((m5stg_rnd_mode[1:0]==2'b10) && (!m5stg_sign)
					&& (m5stg_frac[31:0]!=32'b0))
				|| ((m5stg_rnd_mode[1:0]==2'b11) && m5stg_sign
                                        && (m5stg_frac[31:0]!=32'b0))
				|| ((m5stg_rnd_mode[1:0]==2'b00)
                                        && m5stg_frac[31]
					&& ((m5stg_frac[30:0]!=31'b0)
						|| m5stg_frac[32])))
			&& m5stg_fmuls);
assign m5stg_to_0= (m5stg_rnd_mode[1:0]==2'b01)
                || ((m5stg_rnd_mode[1:0]==2'b10) && m5stg_sign)
                || ((m5stg_rnd_mode[1:0]==2'b11) && (!m5stg_sign));
assign m5stg_to_0_inv= (!m5stg_to_0);
assign mul_frac_out_fracadd= m5stg_rndup && (!m5stg_in_of);
assign mul_frac_out_frac= (!m5stg_rndup) && (!m5stg_in_of);
assign mul_exp_out_exp_plus1= m5stg_rndup && (!m5stg_in_of);
assign mul_exp_out_exp= (!m5stg_rndup) && (!m5stg_in_of);
endmodule
module fpu_mul_exp_dp (
	inq_in1,
	inq_in2,
	m6stg_step,
	m1stg_dblop,
	m1stg_sngop,
	m2stg_exp_expadd,
	m2stg_exp_0bff,
	m2stg_exp_017f,
	m2stg_exp_04ff,
	m2stg_exp_zero,
	m1stg_fsmuld,
	m2stg_fmuld,
	m2stg_fmuls,
	m2stg_fsmuld,
	m3stg_ld0_inv,
	m5stg_fracadd_cout,
	mul_exp_out_exp_plus1,
	mul_exp_out_exp,
	m5stg_in_of,
	m5stg_fmuld,
	m5stg_to_0_inv,
	m4stg_shl_54,
	m4stg_shl_55,
	m4stg_inc_exp_54,
	m4stg_inc_exp_55,
	m4stg_inc_exp_105,
	fmul_clken_l,
	rclk,
	
	m3stg_exp,
	m3stg_expadd_eq_0,
	m3stg_expadd_lte_0_inv,
	m4stg_exp,
	m5stg_exp,
	mul_exp_out,
	se,
	si,
	so
);
input [62:52]	inq_in1;		
input [62:52]	inq_in2;		
input		m6stg_step;		
input		m1stg_dblop;		
input		m1stg_sngop;		
input		m2stg_exp_expadd;	
input		m2stg_exp_0bff;		
input		m2stg_exp_017f;		
input		m2stg_exp_04ff;		
input		m2stg_exp_zero;		
input		m1stg_fsmuld;		
input		m2stg_fmuld;		
input		m2stg_fmuls;		
input		m2stg_fsmuld;		
input [6:0]	m3stg_ld0_inv;		
input           m4stg_inc_exp_54;       
input           m4stg_inc_exp_55;       
input           m4stg_inc_exp_105;      
input		m5stg_fracadd_cout;	
input		mul_exp_out_exp_plus1;	
input		mul_exp_out_exp;	
input		m5stg_in_of;		
input		m5stg_fmuld;		
input		m5stg_to_0_inv;		
input		m4stg_shl_54;		
input		m4stg_shl_55;		
input		fmul_clken_l;           
input		rclk; 		
output [12:0]	m3stg_exp;		
output		m3stg_expadd_eq_0;	
output		m3stg_expadd_lte_0_inv;	
output [12:0]	m4stg_exp;		
output [12:0]	m5stg_exp;		
output [10:0]	mul_exp_out;		
input           se;                     
input           si;                     
output          so;                     
wire [10:0]	m1stg_exp_in1;
wire [10:0]	m1stg_exp_in2;
wire [12:0]	m1stg_expadd_in1;
wire [12:0]	m1stg_expadd_in2;
wire [12:0]	m1stg_expadd;
wire [12:0]	m2stg_exp_in;
wire [12:0]	m2stg_exp;
wire [12:0]	m2stg_expadd_in2;
wire [12:0]	m2stg_expadd;
wire [12:0]	m3astg_exp;
wire [12:0]	m3bstg_exp;
wire [12:0]	m3stg_exp;
wire [12:0]	m3stg_expa;
wire [12:0]	m3stg_expadd;
wire		m3stg_expadd_eq_0;
wire		m3stg_expadd_lte_0_inv;
wire [12:0]	m4stg_exp_in;
wire [12:0]	m4stg_exp;
wire [12:0]	m4stg_exp_plus1;
wire [12:0]	m5stg_exp_pre1_in;
wire [12:0]	m5stg_exp_pre1;
wire [12:0]	m5stg_exp_pre2_in;
wire [12:0]	m5stg_exp_pre2;
wire [12:0]	m5stg_exp_pre3_in;
wire [12:0]	m5stg_exp_pre3;
wire [12:0]	m5stg_exp;
wire [12:0]	m5stg_expa;
wire [12:0]	m5stg_exp_plus1;
wire [10:0]	mul_exp_out_in;
wire [10:0]	mul_exp_out;
wire se_l;
wire        clk;
wire        m5stg_shl_55;
wire        m5stg_shl_54;
wire        m5stg_inc_exp_54;
wire        m5stg_inc_exp_55;
wire        m5stg_inc_exp_105;
assign se_l = ~se;
    clken_buf  ckbuf_mul_exp_dp (
      .clk(clk),
      .rclk(rclk),
      .enb_l(fmul_clken_l),
      .tmb_l(se_l)
      );
dffe_s #(11) i_m1stg_exp_in1 (
        .din    (inq_in1[62:52]),
        .en     (m6stg_step),
        .clk    (clk),
 
        .q      (m1stg_exp_in1[10:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(11) i_m1stg_exp_in2 (
        .din    (inq_in2[62:52]),
        .en     (m6stg_step),
        .clk    (clk),
 
        .q      (m1stg_exp_in2[10:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign m1stg_expadd_in1[12:0]= ({13{m1stg_dblop}}
			    & {2'b0, m1stg_exp_in1[10:0]})
		| ({13{m1stg_sngop}}
			    & {5'b0, m1stg_exp_in1[10:3]});
assign m1stg_expadd_in2[12:0]= ({13{m1stg_dblop}}
                            & {2'b0, m1stg_exp_in2[10:0]})
                | ({13{m1stg_sngop}}
                            & {5'b0, m1stg_exp_in2[10:3]});
assign m1stg_expadd[12:0]= (m1stg_expadd_in1[12:0]
			+ m1stg_expadd_in2[12:0]
			+ 13'h0001);
assign m2stg_exp_in[12:0]= ({13{m2stg_exp_expadd}}
			    & m1stg_expadd[12:0])
		| ({13{m2stg_exp_0bff}}
			    & 13'h0bff)
		| ({13{m2stg_exp_017f}}
			    & 13'h017f)
		| ({13{m2stg_exp_04ff}}
			    & 13'h04ff)
		| ({13{m2stg_exp_zero}}
			    & {{3{m1stg_fsmuld}}, 10'b0});
dffe_s #(13) i_m2stg_exp (
	.din	(m2stg_exp_in[12:0]),
	.en     (m6stg_step),
        .clk    (clk),
        .q      (m2stg_exp[12:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign m2stg_expadd_in2[12:0]= ({13{m2stg_fmuld}}
			    & 13'h1c00)
		| ({13{m2stg_fmuls}}
			    & 13'h1f80)
		| ({13{m2stg_fsmuld}}
			    & 13'h0300);
assign m2stg_expadd[12:0]= m2stg_exp[12:0]
			+ m2stg_expadd_in2[12:0];
dffe_s #(13) i_m3astg_exp (
	.din	(m2stg_expadd[12:0]),
	.en     (m6stg_step),
        .clk    (clk),
        .q      (m3astg_exp[12:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(13) i_m3bstg_exp (
        .din    (m3astg_exp[12:0]),
	.en     (m6stg_step),
        .clk    (clk),
        .q      (m3bstg_exp[12:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(13) i_m3stg_exp (
        .din    (m3bstg_exp[12:0]),
        .en     (m6stg_step),
        .clk    (clk),
        .q      (m3stg_exp[12:0]),
 
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(13) i_m3stg_expa (
	.din	(m3bstg_exp[12:0]),
	.en	(m6stg_step),
	.clk	(clk),
	.q	(m3stg_expa[12:0]),
	.se	(se),
	.si	(),
  	.so	()
);
assign m3stg_expadd[12:0]= (m3stg_expa[12:0]
			+ {6'h3f, m3stg_ld0_inv[6:0]}
			+ 13'h0001);
assign m3stg_expadd_eq_0= (&(m3stg_exp[12:0] ^ {6'h3f, m3stg_ld0_inv[6:0]}));
assign m3stg_expadd_lte_0_inv= (!(m3stg_expadd[12] || m3stg_expadd_eq_0));
assign m4stg_exp_in[12:0]= (m3stg_expadd[12:0] & {13{(!m3stg_expadd[12])}});
dffe_s #(13) i_m4stg_exp (
        .din    (m4stg_exp_in[12:0]),
	.en     (m6stg_step),
        .clk    (clk),
        .q      (m4stg_exp[12:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign m4stg_exp_plus1[12:0]= m4stg_exp[12:0]
			+ 13'h0001;
assign m5stg_exp_pre1_in[12:0]= ( ({13{m6stg_step}}
			    & m4stg_exp_plus1[12:0]));
dff_s #(13) i_m5stg_exp_pre1 (
	.din	(m5stg_exp_pre1_in[12:0]),
	.clk    (clk),
 
        .q      (m5stg_exp_pre1[12:0]),
 
        .se     (se),
        .si     (),
        .so     ()
);
assign m5stg_exp_pre2_in[12:0]= ( ({13{m6stg_step}}
			    & m4stg_exp[12:0]));
dff_s #(13) i_m5stg_exp_pre2 (
	.din	(m5stg_exp_pre2_in[12:0]),
	.clk	(clk),
	.q	(m5stg_exp_pre2[12:0]),
	.se	(se),
	 .si	(),
	.so	()
);
assign m5stg_exp_pre3_in[12:0]= (~({13{(!m6stg_step)}}
			    & m5stg_expa[12:0]));
dff_s #(13) i_m5stg_exp_pre3 (
	.din	(m5stg_exp_pre3_in[12:0]),
	.clk	(clk),
	.q	(m5stg_exp_pre3[12:0]),
	.se	(se),
	 .si	(),
	.so	()
);
dff_s #(5) i_m5stg_inc_exp (
	.din	({m4stg_shl_55,m4stg_shl_54,
                  m4stg_inc_exp_54,m4stg_inc_exp_55,m4stg_inc_exp_105}),
	.clk	(clk),
	.q	({m5stg_shl_55,m5stg_shl_54,
                  m5stg_inc_exp_54,m5stg_inc_exp_55,m5stg_inc_exp_105}),
	.se	(se),
	.si	(),
	.so	()
);
assign m5stg_exp[12:0] =
          ( {13{((m5stg_shl_54 & m5stg_inc_exp_54) |
                 (m5stg_shl_55 & m5stg_inc_exp_55) |
                 (m5stg_inc_exp_105)                )}} & m5stg_exp_pre1[12:0]) |
          (~{13{((m5stg_shl_54 & m5stg_inc_exp_54) |
                 (m5stg_shl_55 & m5stg_inc_exp_55) |
                 (m5stg_inc_exp_105)                )}} & m5stg_exp_pre2[12:0]) |
         ~(m5stg_exp_pre3[12:0]);
assign m5stg_expa[12:0]= m5stg_exp[12:0];
 
assign m5stg_exp_plus1[12:0]= m5stg_expa[12:0]
                        + 13'h0001;
assign mul_exp_out_in[10:0]= ({11{(mul_exp_out_exp_plus1
					&& m5stg_fracadd_cout)}}
			    & m5stg_exp_plus1[10:0])
		| ({11{mul_exp_out_exp}}
			    & m5stg_expa[10:0])
		| ({11{((!m5stg_fracadd_cout) && (!m5stg_in_of))}}
			    & m5stg_expa[10:0])
		| ({11{m5stg_in_of}}
			    & {{3{m5stg_fmuld}}, 7'h7f, m5stg_to_0_inv});
dffe_s #(11) i_mul_exp_out (
	.din	(mul_exp_out_in[10:0]),
	.en     (m6stg_step),
        .clk    (clk),
        .q      (mul_exp_out[10:0]),
	.se     (se),
        .si     (),
        .so     ()
);
endmodule
module fpu_mul_frac_dp (
	inq_in1,
	inq_in2,
	m6stg_step,
	m2stg_frac1_dbl_norm,
	m2stg_frac1_dbl_dnrm,
	m2stg_frac1_sng_norm,
	m2stg_frac1_sng_dnrm,
	m2stg_frac1_inf,
	m1stg_snan_dbl_in1,
	m1stg_snan_sng_in1,
	m2stg_frac2_dbl_norm,
	m2stg_frac2_dbl_dnrm,
	m2stg_frac2_sng_norm,
	m2stg_frac2_sng_dnrm,
	m2stg_frac2_inf,
	m1stg_snan_dbl_in2,
	m1stg_snan_sng_in2,
	m1stg_inf_zero_in,
	m1stg_inf_zero_in_dbl,
	m1stg_dblop,
	m1stg_dblop_inv,
	m4stg_frac,
	m4stg_sh_cnt_in,
	m3bstg_ld0_inv,
	m4stg_left_shift_step,
	m4stg_right_shift_step,
	m5stg_fmuls,
	m5stg_fmulda,
	mul_frac_out_fracadd,
	mul_frac_out_frac,
	m5stg_in_of,
	m5stg_to_0,
	fmul_clken_l,
	rclk,
	
	m2stg_frac1_array_in,
	m2stg_frac2_array_in,
	m1stg_ld0_1,
	m1stg_ld0_2,
	m4stg_frac_105,
	m3stg_ld0_inv,
	m4stg_shl_54,
	m4stg_shl_55,
	m5stg_frac_32_0,
	m5stg_frac_dbl_nx,
	m5stg_frac_sng_nx,
	m5stg_frac_neq_0,
	m5stg_fracadd_cout,
	mul_frac_out,
	se,
	si,
	so
);
input [54:0]	inq_in1;		
input [54:0]	inq_in2;		
input		m6stg_step;		
input		m2stg_frac1_dbl_norm;	
input		m2stg_frac1_dbl_dnrm;	
input		m2stg_frac1_sng_norm;	
input		m2stg_frac1_sng_dnrm;	
input		m2stg_frac1_inf;	
input		m1stg_snan_dbl_in1;	
input		m1stg_snan_sng_in1;	
input		m2stg_frac2_dbl_norm;	
input		m2stg_frac2_dbl_dnrm;	
input		m2stg_frac2_sng_norm;	
input		m2stg_frac2_sng_dnrm;	
input		m2stg_frac2_inf;	
input		m1stg_snan_dbl_in2;	
input		m1stg_snan_sng_in2;	
input		m1stg_inf_zero_in;	
input		m1stg_inf_zero_in_dbl;	
input		m1stg_dblop;		
input		m1stg_dblop_inv;	
input [105:0]	m4stg_frac;		
input [5:0]	m4stg_sh_cnt_in;	
input [6:0]	m3bstg_ld0_inv;		
input		m4stg_left_shift_step;	
input		m4stg_right_shift_step;	
input		m5stg_fmuls;		
input		m5stg_fmulda;		
input		mul_frac_out_fracadd;	
input		mul_frac_out_frac;	
input		m5stg_in_of;		
input		m5stg_to_0;		
input		fmul_clken_l;           
input		rclk;		
output [52:0]	m2stg_frac1_array_in;	
output [52:0]	m2stg_frac2_array_in;	
output [5:0]	m1stg_ld0_1;		
output [5:0]	m1stg_ld0_2;		
output		m4stg_frac_105;		
output [6:0]	m3stg_ld0_inv;		
output		m4stg_shl_54;		
output		m4stg_shl_55;		
output [32:0]	m5stg_frac_32_0;	
output		m5stg_frac_dbl_nx;	
output		m5stg_frac_sng_nx;	
output		m5stg_frac_neq_0;	
output		m5stg_fracadd_cout;	
output [51:0]	mul_frac_out;		
input           se;                     
input           si;                     
output          so;                     
wire [54:0]	mul_frac_in1;
wire [54:0]	mul_frac_in2;
wire [52:0]	m2stg_frac1_in;
wire [52:0]	m2stg_frac1_array_in;
wire [52:0]	m2stg_frac2_in;
wire [52:0]	m2stg_frac2_array_in;
wire [52:0]	m1stg_ld0_1_din;
wire [5:0]	m1stg_ld0_1;
wire [52:0]	m1stg_ld0_2_din;
wire [5:0]	m1stg_ld0_2;
wire		m4stg_frac_105;
wire [5:0]	m4stg_sh_cnt_5;
wire [5:0]	m4stg_sh_cnt_4;
wire [5:0]	m4stg_sh_cnt;
wire [6:0]	m3stg_ld0_inv;
wire [168:63]	m4stg_shl_tmp;
wire [55:0]	m4stg_shl;
wire		m4stg_shl_54;
wire		m4stg_shl_55;
wire [168:0]	m4stg_shr_tmp;
wire [55:0]	m4stg_shr;
wire [54:0]	m5stg_frac_pre1_in;
wire [54:0]	m5stg_frac_pre1;
wire [54:0]	m5stg_frac_pre2_in;
wire [54:0]	m5stg_frac_pre2;
wire [54:0]	m5stg_frac_pre3_in;
wire [54:0]	m5stg_frac_pre3;
wire [54:0]	m5stg_frac_pre4_in;
wire [54:0]	m5stg_frac_pre4;
wire [54:33]	m5stg_frac_54_33;
wire [32:0]	m5stg_frac_32_0;
wire [54:3]	m5stg_fraca;
wire [54:0]	m5stg_fracb;
wire		m5stg_frac_dbl_nx;
wire		m5stg_frac_sng_nx;
wire		m5stg_frac_neq_0;
wire [52:0]	m5stg_fracadd_tmp;
wire		m5stg_fracadd_cout;
wire [51:0]	m5stg_fracadd;
wire [51:0]	mul_frac_out_in;
wire [51:0]	mul_frac_out;
wire [30:0] mstg_xtra_regs;
wire se_l;
wire        clk;
assign se_l = ~se;
    clken_buf  ckbuf_mul_frac_dp (
      .clk(clk),
      .rclk(rclk),
      .enb_l(fmul_clken_l),
      .tmb_l(se_l)
      );
dffe_s #(55) i_mul_frac_in1 (
        .din    (inq_in1[54:0]),
        .en     (m6stg_step),
        .clk    (clk),
 
        .q      (mul_frac_in1[54:0]),
        .se     (se),
        .si     (),
        .so     ()
);
dffe_s #(55) i_mul_frac_in2 (
        .din    (inq_in2[54:0]),
        .en     (m6stg_step),
        .clk    (clk),
 
        .q      (mul_frac_in2[54:0]),
        .se     (se),
        .si     (),
        .so     ()
);
assign m2stg_frac1_in[52:0]= ({53{m2stg_frac1_dbl_norm}}
			    & {1'b1, (mul_frac_in1[51] || m1stg_snan_dbl_in1),
				mul_frac_in1[50:0]})
		| ({53{m2stg_frac1_dbl_dnrm}}
                            & {mul_frac_in1[51:0], 1'b0})
                | ({53{m2stg_frac1_sng_norm}}
                            & {1'b1, (mul_frac_in1[54] || m1stg_snan_sng_in1),
                                mul_frac_in1[53:32], 29'b0})
                | ({53{m2stg_frac1_sng_dnrm}}
                            & {mul_frac_in1[54:32], 30'b0})
		| ({53{m2stg_frac1_inf}}
			    & 53'h10000000000000);
assign m2stg_frac1_array_in[52:0]= (~m2stg_frac1_in[52:0]);
assign m2stg_frac2_in[52:0]= ({53{m2stg_frac2_dbl_norm}}
                            & {1'b1, (mul_frac_in2[51] || m1stg_snan_dbl_in2),
                                mul_frac_in2[50:0]})
                | ({53{m2stg_frac2_dbl_dnrm}}
                            & {mul_frac_in2[51:0], 1'b0})
                | ({53{m2stg_frac2_sng_norm}}
                            & {1'b1, (mul_frac_in2[54] || m1stg_snan_sng_in2),
                                mul_frac_in2[53:32], 29'b0})
                | ({53{m2stg_frac2_sng_dnrm}}
                            & {mul_frac_in2[54:32], 30'b0})
                | ({53{m2stg_frac2_inf}}
			    & {1'b1, {23{m1stg_inf_zero_in}},
					{29{m1stg_inf_zero_in_dbl}}});
 
assign m2stg_frac2_array_in[52:0]= m2stg_frac2_in[52:0];
assign m1stg_ld0_1_din[52:0]= ({53{m1stg_dblop_inv}}
			    & {mul_frac_in1[54:32], 30'b0})
		| ({53{m1stg_dblop}}
			    & {mul_frac_in1[51:0], 1'b0});
fpu_cnt_lead0_53b i_m1stg_ld0_1 (
	.din	(m1stg_ld0_1_din[52:0]),
	.lead0	(m1stg_ld0_1[5:0])
);
assign m1stg_ld0_2_din[52:0]= ({53{m1stg_dblop_inv}}
			    & {mul_frac_in2[54:32], 30'b0})
		| ({53{m1stg_dblop}}
			    & {mul_frac_in2[51:0], 1'b0});
fpu_cnt_lead0_53b i_m1stg_ld0_2 (
	.din	(m1stg_ld0_2_din[52:0]),
	.lead0	(m1stg_ld0_2[5:0])
);
assign m4stg_frac_105= m4stg_frac[105];
dffe_s #(56) i_mstg_xtra_regs (
	.din	({{6{m4stg_sh_cnt_in[5]}}, 
			{6{m4stg_sh_cnt_in[4]}},
			m4stg_sh_cnt_in[5:0],
			m3bstg_ld0_inv[6:0],
			31'h0000_0000}),
	.en     (m6stg_step),
        .clk    (clk),
	.q	({m4stg_sh_cnt_5[5:0],
			m4stg_sh_cnt_4[5:0],
			m4stg_sh_cnt[5:0],
			m3stg_ld0_inv[6:0],
			mstg_xtra_regs[30:0]}),
	.se     (se),
        .si     (),
        .so     ()
);
  assign m4stg_shl_tmp[168:63]=  m4stg_frac[105:0]
		<< {m4stg_sh_cnt_5[0], m4stg_sh_cnt[4:0]};
assign m4stg_shl[55:0]= {m4stg_shl_tmp[168:114], (|m4stg_shl_tmp[113:63])};
assign m4stg_shl_54= m4stg_shl[54];
assign m4stg_shl_55= m4stg_shl[55];
  assign m4stg_shr_tmp[168:0]= {       m4stg_frac[105:0], 63'b0} >> m4stg_sh_cnt[5:0];
assign m4stg_shr[55:0]= {m4stg_shr_tmp[168:114], (|m4stg_shr_tmp[113:0])};
assign m5stg_frac_pre1_in[54:0]= ~(({55{(m4stg_left_shift_step && m4stg_shl[55])}}
			    & m4stg_shl[54:0])
		| ({55{(!m6stg_step)}}
			    & m5stg_fracb[54:0]));
dff_s #(55) i_m5stg_frac_pre1 (
	.din	(m5stg_frac_pre1_in[54:0]),
	.clk    (clk),
        .q      (m5stg_frac_pre1[54:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign m5stg_frac_pre2_in[54:0]= ~({55{(m4stg_left_shift_step
					&& (!m4stg_shl[55]))}}
			    & {m4stg_shl[53:0], 1'b0});
dff_s #(55) i_m5stg_frac_pre2 (
	.din	(m5stg_frac_pre2_in[54:0]),
	.clk	(clk),
	.q	(m5stg_frac_pre2[54:0]),
	.se	(se),
		.si	(),
	.so	()
);
assign m5stg_frac_pre3_in[54:0]= ~({55{(m4stg_right_shift_step
					&& m4stg_shr[55])}}
			    & m4stg_shr[54:0]);
dff_s #(55) i_m5stg_frac_pre3 (
	.din	(m5stg_frac_pre3_in[54:0]),
	.clk	(clk),
	.q	(m5stg_frac_pre3[54:0]),
	.se	(se),
		.si	(),
	.so	()
);
assign m5stg_frac_pre4_in[54:0]= ~({55{(m4stg_right_shift_step
					&& (!m4stg_shr[55]))}}
			    & {m4stg_shr[53:0], 1'b0});
dff_s #(55) i_m5stg_frac_pre4 (
	.din	(m5stg_frac_pre4_in[54:0]),
	.clk	(clk),
	.q	(m5stg_frac_pre4[54:0]),
	.se	(se),
		.si	(),
	.so	()
);
assign {m5stg_frac_54_33[54:33], m5stg_frac_32_0[32:0]} = ~(m5stg_frac_pre1[54:0]
		& m5stg_frac_pre2[54:0]
		& m5stg_frac_pre3[54:0]
		& m5stg_frac_pre4[54:0]);
assign m5stg_fraca[54:3]= {m5stg_frac_54_33[54:33], m5stg_frac_32_0[32:3]};
assign m5stg_fracb[54:0]= {m5stg_frac_54_33[54:33], m5stg_frac_32_0[32:0]};
assign m5stg_frac_dbl_nx= (|m5stg_fracb[2:0]);
assign m5stg_frac_sng_nx= m5stg_frac_dbl_nx || (|m5stg_fracb[31:3]);
assign m5stg_frac_neq_0= m5stg_frac_sng_nx || (|m5stg_fracb[54:32]);
assign m5stg_fracadd_tmp[52:0]= {1'b0, m5stg_fraca[54:3]}
			+ {23'b0, m5stg_fmuls, 28'b0, m5stg_fmulda};
assign m5stg_fracadd_cout= m5stg_fracadd_tmp[52];
assign m5stg_fracadd[51:0]= m5stg_fracadd_tmp[51:0];
assign mul_frac_out_in[51:0]= ({52{mul_frac_out_fracadd}}
			    & m5stg_fracadd[51:0])
		| ({52{mul_frac_out_frac}}
			    & m5stg_fracb[54:3])
		| ({52{m5stg_in_of}}
			    & {52{m5stg_to_0}});
dffe_s #(52) i_mul_frac_out (
	.din	(mul_frac_out_in[51:0]),
	.en     (m6stg_step),
        .clk    (clk),
        .q      (mul_frac_out[51:0]),
	.se     (se),
        .si     (),
        .so     ()
);
endmodule
module fpu_out (
	d8stg_fdiv_in,
	m6stg_fmul_in,
	a6stg_fadd_in,
	div_id_out_in,
	m6stg_id_in,
	add_id_out_in,
	div_exc_out,
	d8stg_fdivd,
	d8stg_fdivs,
	div_sign_out,
	div_exp_out,
	div_frac_out,
	mul_exc_out,
	m6stg_fmul_dbl_dst,
	m6stg_fmuls,
	mul_sign_out,
	mul_exp_out,
	mul_frac_out,
	add_exc_out,
	a6stg_fcmpop,
	add_cc_out,
	add_fcc_out,
	a6stg_dbl_dst,
	a6stg_sng_dst,
	a6stg_long_dst,
	a6stg_int_dst,
	add_sign_out,
	add_exp_out,
	add_frac_out,
	arst_l,
	grst_l,
	rclk,
	
	fp_cpx_req_cq,
	add_dest_rdy,
	mul_dest_rdy,
	div_dest_rdy,
	fp_cpx_data_ca,
	se,
	si,
	so
);
input		d8stg_fdiv_in;		
input		m6stg_fmul_in;		
input		a6stg_fadd_in;		
input [9:0]	div_id_out_in;		
input [9:0]	m6stg_id_in;		
input [9:0]	add_id_out_in;		
input [4:0]	div_exc_out;		
input		d8stg_fdivd;		
input		d8stg_fdivs;		
input		div_sign_out;		
input [10:0]	div_exp_out;		
input [51:0]	div_frac_out;		
input [4:0]	mul_exc_out;		
input		m6stg_fmul_dbl_dst;	
input		m6stg_fmuls;		
input		mul_sign_out;		
input [10:0]	mul_exp_out;		
input [51:0]	mul_frac_out;		
input [4:0]	add_exc_out;		
input		a6stg_fcmpop;		
input [1:0]	add_cc_out;		
input [1:0]	add_fcc_out;		
input		a6stg_dbl_dst;		
input		a6stg_sng_dst;		
input		a6stg_long_dst;		
input		a6stg_int_dst;		
input		add_sign_out;		
input [10:0]	add_exp_out;		
input [63:0]	add_frac_out;		
input		arst_l;			
input		grst_l;			
input		rclk;			
output [7:0]	fp_cpx_req_cq;		
output		add_dest_rdy;		
output		mul_dest_rdy;		
output		div_dest_rdy;		
output [144:0]	fp_cpx_data_ca;		
input           se;                     
input           si;                     
output          so;                     
wire [7:0]	fp_cpx_req_cq;		
wire [1:0]	req_thread;		
wire [2:0]	dest_rdy;		
wire		add_dest_rdy;		
wire		mul_dest_rdy;		
wire		div_dest_rdy;		
wire [144:0]	fp_cpx_data_ca;		
wire        scan_out_fpu_out_ctl;
fpu_out_ctl fpu_out_ctl (
	.d8stg_fdiv_in			(d8stg_fdiv_in),
	.m6stg_fmul_in			(m6stg_fmul_in),
	.a6stg_fadd_in			(a6stg_fadd_in),
	.div_id_out_in			(div_id_out_in[9:0]),
	.m6stg_id_in			(m6stg_id_in[9:0]),
	.add_id_out_in			(add_id_out_in[9:0]),
	.arst_l				(arst_l),
	.grst_l				(grst_l),
	.rclk			(rclk),
	.fp_cpx_req_cq			(fp_cpx_req_cq[7:0]),
	.req_thread			(req_thread[1:0]),
	.dest_rdy			(dest_rdy[2:0]),
	.add_dest_rdy			(add_dest_rdy),
	.mul_dest_rdy			(mul_dest_rdy),
	.div_dest_rdy			(div_dest_rdy),
	.se                             (se),
        .si                             (si),
        .so                             (scan_out_fpu_out_ctl)
);
fpu_out_dp fpu_out_dp (
	.dest_rdy			(dest_rdy[2:0]),
	.req_thread			(req_thread[1:0]),
	.div_exc_out			(div_exc_out[4:0]),
	.d8stg_fdivd			(d8stg_fdivd),
	.d8stg_fdivs			(d8stg_fdivs),
	.div_sign_out			(div_sign_out),
	.div_exp_out			(div_exp_out[10:0]),
	.div_frac_out			(div_frac_out[51:0]),
	.mul_exc_out			(mul_exc_out[4:0]),
	.m6stg_fmul_dbl_dst		(m6stg_fmul_dbl_dst),
	.m6stg_fmuls			(m6stg_fmuls),
	.mul_sign_out			(mul_sign_out),
	.mul_exp_out			(mul_exp_out[10:0]),
	.mul_frac_out			(mul_frac_out[51:0]),
	.add_exc_out			(add_exc_out[4:0]),
	.a6stg_fcmpop			(a6stg_fcmpop),
	.add_cc_out			(add_cc_out[1:0]),
	.add_fcc_out			(add_fcc_out[1:0]),
	.a6stg_dbl_dst			(a6stg_dbl_dst),
	.a6stg_sng_dst			(a6stg_sng_dst),
	.a6stg_long_dst			(a6stg_long_dst),
	.a6stg_int_dst			(a6stg_int_dst),
	.add_sign_out			(add_sign_out),
	.add_exp_out			(add_exp_out[10:0]),
	.add_frac_out			(add_frac_out[63:0]),
	.rclk			(rclk),
	.fp_cpx_data_ca			(fp_cpx_data_ca[144:0]),
	.se                             (se),
        .si                             (scan_out_fpu_out_ctl),
        .so                             (so)
);
endmodule
 
module fpu_out_ctl (
	d8stg_fdiv_in,
	m6stg_fmul_in,
	a6stg_fadd_in,
	div_id_out_in,
	m6stg_id_in,
	add_id_out_in,
	arst_l,
	grst_l,
	rclk,
	
	fp_cpx_req_cq,
	req_thread,
	dest_rdy,
	add_dest_rdy,
	mul_dest_rdy,
	div_dest_rdy,
	se,
	si,
	so
);
input		d8stg_fdiv_in;		
input		m6stg_fmul_in;		
input		a6stg_fadd_in;		
input [9:0]	div_id_out_in;		
input [9:0]	m6stg_id_in;		
input [9:0]	add_id_out_in;		
input		arst_l;			
input		grst_l;			
input		rclk;		
output [7:0]	fp_cpx_req_cq;		
output [1:0]	req_thread;		
output [2:0]	dest_rdy;		
output		add_dest_rdy;		
output		mul_dest_rdy;		
output		div_dest_rdy;		
input           se;                     
input           si;                     
output          so;                     
wire		reset;
wire		add_req_in;
wire		add_req_step;
wire		add_req;
wire		div_req_sel;
wire		mul_req_sel;
wire		add_req_sel;
wire [9:0]	out_id;
wire [7:0]	fp_cpx_req_cq;
wire [1:0]	req_thread;
wire [2:0]	dest_rdy_in;
wire [2:0]	dest_rdy;
wire		add_dest_rdy;
wire		mul_dest_rdy;
wire		div_dest_rdy;
wire        out_ctl_rst_l;
dffrl_async #(1)  dffrl_out_ctl (
  .din  (grst_l),
  .clk  (rclk),
  .rst_l(arst_l),
  .q    (out_ctl_rst_l),
	.se (se),
	.si (),
	.so ()
  );
assign reset= (!out_ctl_rst_l);
assign add_req_in= (!add_req);
assign add_req_step= add_req_sel || mul_req_sel;
dffre_s #(1) i_add_req (
	.din	(add_req_in),
	.en	(add_req_step),
	.rst    (reset),
        .clk    (rclk),
        .q      (add_req),
	.se     (se),
        .si     (),
        .so     ()
);
assign div_req_sel= d8stg_fdiv_in;
assign mul_req_sel= m6stg_fmul_in
		&& ((!add_req) || (!a6stg_fadd_in))
		&& (!div_req_sel);
assign add_req_sel= a6stg_fadd_in
		&& (add_req || (!m6stg_fmul_in))
		&& (!div_req_sel);
assign out_id[9:0]= ({10{div_req_sel}}
			    & div_id_out_in[9:0])
		| ({10{mul_req_sel}}
			    & m6stg_id_in[9:0])
		| ({10{add_req_sel}}
			    & add_id_out_in[9:0]);
dff_s #(8) i_fp_cpx_req_cq (
	.din	(out_id[9:2]),
	.clk    (rclk),
        .q      (fp_cpx_req_cq[7:0]),
	.se     (se),
        .si     (),
        .so     ()
);
dff_s #(2) i_req_thread (
	.din	(out_id[1:0]),
	.clk    (rclk),
 
        .q      (req_thread[1:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign dest_rdy_in[2:0]= {div_req_sel, mul_req_sel, add_req_sel};
dff_s #(3) i_dest_rdy (
	.din	(dest_rdy_in[2:0]),
	.clk    (rclk),
        .q      (dest_rdy[2:0]),
	.se     (se),
        .si     (),
        .so     ()
);
dff_s i_add_dest_rdy (
	.din	(add_req_sel),
	.clk	(rclk),
	.q	(add_dest_rdy),
	.se	(se),
        .si	(),
        .so	()
);
dff_s i_mul_dest_rdy (
	.din	(mul_req_sel),
	.clk	(rclk),
	.q	(mul_dest_rdy),
	.se	(se),
        .si	(),
        .so	()
);
dff_s i_div_dest_rdy (
	.din	(div_req_sel),
	.clk	(rclk),
	.q	(div_dest_rdy),
        .se	(se),
        .si	(),
        .so	()
);
endmodule
 
module fpu_out_dp (
	dest_rdy,
	req_thread,
	div_exc_out,
	d8stg_fdivd,
	d8stg_fdivs,
	div_sign_out,
	div_exp_out,
	div_frac_out,
	mul_exc_out,
	m6stg_fmul_dbl_dst,
	m6stg_fmuls,
	mul_sign_out,
	mul_exp_out,
	mul_frac_out,
	add_exc_out,
	a6stg_fcmpop,
	add_cc_out,
	add_fcc_out,
	a6stg_dbl_dst,
	a6stg_sng_dst,
	a6stg_long_dst,
	a6stg_int_dst,
	add_sign_out,
	add_exp_out,
	add_frac_out,
	rclk,
	
	fp_cpx_data_ca,
	se,
	si,
	so
);
input [2:0]	dest_rdy;		
input [1:0]	req_thread;		
input [4:0]	div_exc_out;		
input		d8stg_fdivd;		
input		d8stg_fdivs;		
input		div_sign_out;		
input [10:0]	div_exp_out;		
input [51:0]	div_frac_out;		
input [4:0]	mul_exc_out;		
input		m6stg_fmul_dbl_dst;	
input		m6stg_fmuls;		
input		mul_sign_out;		
input [10:0]	mul_exp_out;		
input [51:0]	mul_frac_out;		
input [4:0]	add_exc_out;		
input		a6stg_fcmpop;		
input [1:0]	add_cc_out;		
input [1:0]	add_fcc_out;		
input		a6stg_dbl_dst;		
input		a6stg_sng_dst;		
input		a6stg_long_dst;		
input		a6stg_int_dst;		
input		add_sign_out;		
input [10:0]	add_exp_out;		
input [63:0]	add_frac_out;		
input		rclk;		
output [144:0]	fp_cpx_data_ca;		
input           se;                     
input           si;                     
output          so;                     
wire [63:0]	add_out;
wire [63:0]	mul_out;
wire [63:0]	div_out;
wire [7:0]	fp_cpx_data_ca_84_77_in;
wire [76:0]	fp_cpx_data_ca_76_0_in;
wire [7:0]	fp_cpx_data_ca_84_77;
wire [76:0]	fp_cpx_data_ca_76_0;
wire [144:0]	fp_cpx_data_ca;
wire se_l;
wire        clk;
assign se_l = ~se;
clken_buf  ckbuf_out_dp (
  .clk(clk),
  .rclk(rclk),
  .enb_l(1'b0),
  .tmb_l(se_l)
  );
assign add_out[63:0]= ({64{a6stg_dbl_dst}}
			    & {add_sign_out, add_exp_out[10:0],
				add_frac_out[62:11]})
		| ({64{a6stg_sng_dst}}
			    & {add_sign_out, add_exp_out[7:0],
				add_frac_out[62:40], 32'b0})
		| ({64{a6stg_long_dst}}
			    & add_frac_out[63:0])
		| ({64{a6stg_int_dst}}
			    & {add_frac_out[63:32], 32'b0});
assign mul_out[63:0]= ({64{m6stg_fmul_dbl_dst}}
			    & {mul_sign_out, mul_exp_out[10:0],
				mul_frac_out[51:0]})
		| ({64{m6stg_fmuls}}
			    & {mul_sign_out, mul_exp_out[7:0],
				mul_frac_out[51:29], 32'b0});
assign div_out[63:0]= ({64{d8stg_fdivd}}
			    & {div_sign_out, div_exp_out[10:0],
				div_frac_out[51:0]})
		| ({64{d8stg_fdivs}}
			    & {div_sign_out, div_exp_out[7:0],
				div_frac_out[51:29], 32'b0});
assign fp_cpx_data_ca_84_77_in[7:0]= ({8{(|dest_rdy)}}
			    & {1'b1, 4'b1000, 1'b0, req_thread[1:0]});
assign fp_cpx_data_ca_76_0_in[76:0]= ({77{dest_rdy[2]}}
			    & {div_exc_out[4:0], 8'b0, div_out[63:0]})
		| ({77{dest_rdy[1]}}
			    & {mul_exc_out[4:0], 8'b0, mul_out[63:0]})
		| ({77{dest_rdy[0]}}
			    & {add_exc_out[4:0], 2'b0, a6stg_fcmpop,
				add_cc_out[1:0], add_fcc_out[1:0], 1'b0,
				add_out[63:0]});
dff_s #(8) i_fp_cpx_data_ca_84_77 (
	.din	(fp_cpx_data_ca_84_77_in[7:0]),
	.clk    (clk),
        .q      (fp_cpx_data_ca_84_77[7:0]),
	.se     (se),
        .si     (),
        .so     ()
);
dff_s #(77) i_fp_cpx_data_ca_76_0 (
	.din	(fp_cpx_data_ca_76_0_in[76:0]),
	.clk    (clk),
        .q      (fp_cpx_data_ca_76_0[76:0]),
	.se     (se),
        .si     (),
        .so     ()
);
assign fp_cpx_data_ca[144:0]= {fp_cpx_data_ca_84_77[7:3],
				3'b0,
				fp_cpx_data_ca_84_77[2:0],
				57'b0,
				fp_cpx_data_ca_76_0[76:0]};
endmodule
module fpu_bufrpt_grp64 (
	in,
	out
);
	
	input [63:0] in;
	output [63:0] out;
	assign out[63:0] = in[63:0];
endmodule
module fpu_bufrpt_grp32 (
	in,
	out
);
	input [31:0] in;
	output [31:0] out;
	assign out[31:0] = in[31:0];
endmodule
module fpu_rptr_groups (
	inq_in1,
	inq_in2,
	inq_id,
	inq_op,
	inq_rnd_mode,
	inq_in1_50_0_neq_0,
	inq_in1_53_0_neq_0,
	inq_in1_53_32_neq_0,
	inq_in1_exp_eq_0,
	inq_in1_exp_neq_ffs,
	inq_in2_50_0_neq_0,
	inq_in2_53_0_neq_0,
	inq_in2_53_32_neq_0,
	inq_in2_exp_eq_0,
	inq_in2_exp_neq_ffs,
	ctu_tst_macrotest,
	ctu_tst_pre_grst_l,
	ctu_tst_scan_disable,
	ctu_tst_scanmode,
	ctu_tst_short_chain,
	global_shift_enable,
	grst_l,
	cluster_cken,
	se,
	arst_l,
	fpu_grst_l,
	fmul_clken_l,
	fdiv_clken_l,
	scan_manual_6,
	si,
	so_unbuf,
	pcx_fpio_data_px2,
	pcx_fpio_data_rdy_px2,
	fp_cpx_req_cq,
	fp_cpx_data_ca,
	inq_sram_din_unbuf,
	inq_in1_add_buf1,
	inq_in1_mul_buf1,
	inq_in1_div_buf1,
	inq_in2_add_buf1,
	inq_in2_mul_buf1,
	inq_in2_div_buf1,
	inq_id_add_buf1,
	inq_id_mul_buf1,
	inq_id_div_buf1,
	inq_op_add_buf1,
	inq_op_div_buf1,
	inq_op_mul_buf1,
	inq_rnd_mode_add_buf1,
	inq_rnd_mode_div_buf1,
	inq_rnd_mode_mul_buf1,
	inq_in1_50_0_neq_0_add_buf1,
	inq_in1_50_0_neq_0_mul_buf1,
	inq_in1_50_0_neq_0_div_buf1,
	inq_in1_53_0_neq_0_add_buf1,
	inq_in1_53_0_neq_0_mul_buf1,
	inq_in1_53_0_neq_0_div_buf1,
	inq_in1_53_32_neq_0_add_buf1,
	inq_in1_53_32_neq_0_mul_buf1,
	inq_in1_53_32_neq_0_div_buf1,
	inq_in1_exp_eq_0_add_buf1,
	inq_in1_exp_eq_0_mul_buf1,
	inq_in1_exp_eq_0_div_buf1,
	inq_in1_exp_neq_ffs_add_buf1,
	inq_in1_exp_neq_ffs_mul_buf1,
	inq_in1_exp_neq_ffs_div_buf1,
	inq_in2_50_0_neq_0_add_buf1,
	inq_in2_50_0_neq_0_mul_buf1,
	inq_in2_50_0_neq_0_div_buf1,
	inq_in2_53_0_neq_0_add_buf1,
	inq_in2_53_0_neq_0_mul_buf1,
	inq_in2_53_0_neq_0_div_buf1,
	inq_in2_53_32_neq_0_add_buf1,
	inq_in2_53_32_neq_0_mul_buf1,
	inq_in2_53_32_neq_0_div_buf1,
	inq_in2_exp_eq_0_add_buf1,
	inq_in2_exp_eq_0_mul_buf1,
	inq_in2_exp_eq_0_div_buf1,
	inq_in2_exp_neq_ffs_add_buf1,
	inq_in2_exp_neq_ffs_mul_buf1,
	inq_in2_exp_neq_ffs_div_buf1,
	ctu_tst_macrotest_buf1,
	ctu_tst_pre_grst_l_buf1,
	ctu_tst_scan_disable_buf1,
	ctu_tst_scanmode_buf1,
	ctu_tst_short_chain_buf1,
	global_shift_enable_buf1,
	grst_l_buf1,
	cluster_cken_buf1,
	se_add_exp_buf2,
	se_add_frac_buf2,
	se_out_buf2,
	se_mul64_buf2,
	se_cluster_header_buf2,
	se_in_buf3,
	se_mul_buf4,
	se_div_buf5,
	arst_l_div_buf2,
	arst_l_mul_buf2,
	arst_l_cluster_header_buf2,
	arst_l_in_buf3,
	arst_l_out_buf3,
	arst_l_add_buf4,
	fpu_grst_l_mul_buf1,
	fpu_grst_l_in_buf2,
	fpu_grst_l_add_buf3,
	fmul_clken_l_buf1,
	fdiv_clken_l_div_exp_buf1,
	fdiv_clken_l_div_frac_buf1,
	scan_manual_6_buf1,
	si_buf1,
	so,
	pcx_fpio_data_px2_buf1,
	pcx_fpio_data_rdy_px2_buf1,
	fp_cpx_req_cq_buf1,
	fp_cpx_data_ca_buf1,
	inq_sram_din_buf1
);
	input [63:0] inq_in1;
	input [63:0] inq_in2;
	input [4:0] inq_id;
	input [7:0] inq_op;
	input [1:0] inq_rnd_mode;
	input inq_in1_50_0_neq_0;
	input inq_in1_53_0_neq_0;
	input inq_in1_53_32_neq_0;
	input inq_in1_exp_eq_0;
	input inq_in1_exp_neq_ffs;
	input inq_in2_50_0_neq_0;
	input inq_in2_53_0_neq_0;
	input inq_in2_53_32_neq_0;
	input inq_in2_exp_eq_0;
	input inq_in2_exp_neq_ffs;
	input ctu_tst_macrotest;
	input ctu_tst_pre_grst_l;
	input ctu_tst_scan_disable;
	input ctu_tst_scanmode;
	input ctu_tst_short_chain;
	input global_shift_enable;
	input grst_l;
	input cluster_cken;
	input se;
	input arst_l;
	input fpu_grst_l;
	input fmul_clken_l;
	input fdiv_clken_l;
	input scan_manual_6;
	input si;
	input so_unbuf;
	input [123:0] pcx_fpio_data_px2;
	input pcx_fpio_data_rdy_px2;
	input [7:0] fp_cpx_req_cq;
	input [144:0] fp_cpx_data_ca;
	input [155:0] inq_sram_din_unbuf;
	output [63:0] inq_in1_add_buf1;
	output [63:0] inq_in1_mul_buf1;
	output [63:0] inq_in1_div_buf1;
	output [63:0] inq_in2_add_buf1;
	output [63:0] inq_in2_mul_buf1;
	output [63:0] inq_in2_div_buf1;
	output [4:0] inq_id_add_buf1;
	output [4:0] inq_id_mul_buf1;
	output [4:0] inq_id_div_buf1;
	output [7:0] inq_op_add_buf1;
	output [7:0] inq_op_mul_buf1;
	output [7:0] inq_op_div_buf1;
	output [1:0] inq_rnd_mode_add_buf1;
	output [1:0] inq_rnd_mode_mul_buf1;
	output [1:0] inq_rnd_mode_div_buf1;
	output inq_in1_50_0_neq_0_add_buf1;
	output inq_in1_50_0_neq_0_mul_buf1;
	output inq_in1_50_0_neq_0_div_buf1;
	output inq_in1_53_0_neq_0_add_buf1;
	output inq_in1_53_0_neq_0_mul_buf1;
	output inq_in1_53_0_neq_0_div_buf1;
	output inq_in1_53_32_neq_0_add_buf1;
	output inq_in1_53_32_neq_0_mul_buf1;
	output inq_in1_53_32_neq_0_div_buf1;
	output inq_in1_exp_eq_0_add_buf1;
	output inq_in1_exp_eq_0_mul_buf1;
	output inq_in1_exp_eq_0_div_buf1;
	output inq_in1_exp_neq_ffs_add_buf1;
	output inq_in1_exp_neq_ffs_mul_buf1;
	output inq_in1_exp_neq_ffs_div_buf1;
	output inq_in2_50_0_neq_0_add_buf1;
	output inq_in2_50_0_neq_0_mul_buf1;
	output inq_in2_50_0_neq_0_div_buf1;
	output inq_in2_53_0_neq_0_add_buf1;
	output inq_in2_53_0_neq_0_mul_buf1;
	output inq_in2_53_0_neq_0_div_buf1;
	output inq_in2_53_32_neq_0_add_buf1;
	output inq_in2_53_32_neq_0_mul_buf1;
	output inq_in2_53_32_neq_0_div_buf1;
	output inq_in2_exp_eq_0_add_buf1;
	output inq_in2_exp_eq_0_mul_buf1;
	output inq_in2_exp_eq_0_div_buf1;
	output inq_in2_exp_neq_ffs_add_buf1;
	output inq_in2_exp_neq_ffs_mul_buf1;
	output inq_in2_exp_neq_ffs_div_buf1;
	output ctu_tst_macrotest_buf1;
	output ctu_tst_pre_grst_l_buf1;
	output ctu_tst_scan_disable_buf1;
	output ctu_tst_scanmode_buf1;
	output ctu_tst_short_chain_buf1;
	output global_shift_enable_buf1;
	output grst_l_buf1;
	output cluster_cken_buf1;
	output se_add_exp_buf2;
	output se_add_frac_buf2;
	output se_out_buf2;
	output se_mul64_buf2;
	output se_cluster_header_buf2;
	output se_in_buf3;
	output se_mul_buf4;
	output se_div_buf5;
	output arst_l_div_buf2;
	output arst_l_mul_buf2;
	output arst_l_cluster_header_buf2;
	output arst_l_in_buf3;
	output arst_l_out_buf3;
	output arst_l_add_buf4;
	output fpu_grst_l_mul_buf1;
	output fpu_grst_l_in_buf2;
	output fpu_grst_l_add_buf3;
	output fmul_clken_l_buf1;
	output fdiv_clken_l_div_exp_buf1;
	output fdiv_clken_l_div_frac_buf1;
	output scan_manual_6_buf1;
	output si_buf1;
	output so;
	output [123:0] pcx_fpio_data_px2_buf1;
	output pcx_fpio_data_rdy_px2_buf1;
	output [7:0] fp_cpx_req_cq_buf1;
	output [144:0] fp_cpx_data_ca_buf1;
	output [155:0] inq_sram_din_buf1;
	wire [3:0] inq_id_add_buf1_unused;
	wire [2:0] inq_id_mul_buf1_unused;
	wire [4:0] inq_id_div_buf1_unused;
	wire [1:0] ctu_tst_buf1_lo_unused;
	wire [1:0] cluster_cken_buf1_unused;
	wire [1:0] se_mul64_buf2_unused;
	wire [2:0] arst_l_buf1_unused;
	wire [1:0] fdiv_clken_l_buf1_unused;
	wire [2:0] so_cluster_header_buf1_unused;
	wire [2:0] si_buf1_unused;
	wire [2:0] pcx_fpio_data_px2_buf1_unused;
	wire [5:0] fp_cpx_buf1_9_unused;
    
    wire        se_add_buf1;
    wire        se_mul64_buf1;
    wire        so_buf1;
    wire        se_buf1_unused;
    wire        se_add_buf2_unused;
    wire        arst_l_buf1;
	
	fpu_bufrpt_grp32 i_inq_in1_add_buf1_hi (
		.in (inq_in1[63:32]),
		.out (inq_in1_add_buf1[63:32])
	);
	fpu_bufrpt_grp32 i_inq_in1_add_buf1_lo (
		.in (inq_in1[31:0]),
		.out (inq_in1_add_buf1[31:0])
	);
	fpu_bufrpt_grp32 i_inq_in1_mul_buf1_hi (
		.in (inq_in1[63:32]),
		.out (inq_in1_mul_buf1[63:32])
	);
	fpu_bufrpt_grp32 i_inq_in1_mul_buf1_lo (
		.in (inq_in1[31:0]),
		.out (inq_in1_mul_buf1[31:0])
	);
	fpu_bufrpt_grp64 i_inq_in1_div_buf1 (
		.in (inq_in1[63:0]),
		.out (inq_in1_div_buf1[63:0])
	);
	
	fpu_bufrpt_grp32 i_inq_in2_add_buf1_hi (
		.in (inq_in2[63:32]),
		.out (inq_in2_add_buf1[63:32])
	);
	fpu_bufrpt_grp32 i_inq_in2_add_buf1_lo (
		.in (inq_in2[31:0]),
		.out (inq_in2_add_buf1[31:0])
	);
	fpu_bufrpt_grp32 i_inq_in2_mul_buf1_hi (
		.in (inq_in2[63:32]),
		.out (inq_in2_mul_buf1[63:32])
	);
	fpu_bufrpt_grp32 i_inq_in2_mul_buf1_lo (
		.in (inq_in2[31:0]),
		.out (inq_in2_mul_buf1[31:0])
	);
	fpu_bufrpt_grp64 i_inq_in2_div_buf1 (
		.in (inq_in2[63:0]),
		.out (inq_in2_div_buf1[63:0])
	);
	
	fpu_bufrpt_grp32 i_inq_id_add_buf1 (
		.in ({4'h0,
			se_out_buf2,
			arst_l_out_buf3,
			fpu_grst_l_in_buf2,
			inq_id[4:0],
			inq_op[7:0],
			inq_rnd_mode[1:0],
			inq_in1_50_0_neq_0,
			inq_in1_53_0_neq_0,
			inq_in1_53_32_neq_0,
			inq_in1_exp_eq_0,
			inq_in1_exp_neq_ffs,
			inq_in2_50_0_neq_0,
			inq_in2_53_0_neq_0,
			inq_in2_53_32_neq_0,
			inq_in2_exp_eq_0,
			inq_in2_exp_neq_ffs}),
		.out ({inq_id_add_buf1_unused[3:0],
			se_in_buf3,
			arst_l_add_buf4,
			fpu_grst_l_add_buf3,
			inq_id_add_buf1[4:0],
			inq_op_add_buf1[7:0],
			inq_rnd_mode_add_buf1[1:0],
			inq_in1_50_0_neq_0_add_buf1,
			inq_in1_53_0_neq_0_add_buf1,
			inq_in1_53_32_neq_0_add_buf1,
			inq_in1_exp_eq_0_add_buf1,
			inq_in1_exp_neq_ffs_add_buf1,
			inq_in2_50_0_neq_0_add_buf1,
			inq_in2_53_0_neq_0_add_buf1,
			inq_in2_53_32_neq_0_add_buf1,
			inq_in2_exp_eq_0_add_buf1,
			inq_in2_exp_neq_ffs_add_buf1})
	);
	fpu_bufrpt_grp32 i_inq_id_mul_buf1 (
		.in ({3'h0,
			se_in_buf3,
			arst_l_mul_buf2,
			fpu_grst_l_mul_buf1,
			fmul_clken_l,
			inq_id[4:0],
			inq_op[7:0],
			inq_rnd_mode[1:0],
			inq_in1_50_0_neq_0,
			inq_in1_53_0_neq_0,
			inq_in1_53_32_neq_0,
			inq_in1_exp_eq_0,
			inq_in1_exp_neq_ffs,
			inq_in2_50_0_neq_0,
			inq_in2_53_0_neq_0,
			inq_in2_53_32_neq_0,
			inq_in2_exp_eq_0,
			inq_in2_exp_neq_ffs}),
		.out ({inq_id_mul_buf1_unused[2:0],
			se_mul_buf4,
			arst_l_out_buf3,
			fpu_grst_l_in_buf2,
			fmul_clken_l_buf1,
			inq_id_mul_buf1[4:0],
			inq_op_mul_buf1[7:0],
			inq_rnd_mode_mul_buf1[1:0],
			inq_in1_50_0_neq_0_mul_buf1,
			inq_in1_53_0_neq_0_mul_buf1,
			inq_in1_53_32_neq_0_mul_buf1,
			inq_in1_exp_eq_0_mul_buf1,
			inq_in1_exp_neq_ffs_mul_buf1,
			inq_in2_50_0_neq_0_mul_buf1,
			inq_in2_53_0_neq_0_mul_buf1,
			inq_in2_53_32_neq_0_mul_buf1,
			inq_in2_exp_eq_0_mul_buf1,
			inq_in2_exp_neq_ffs_mul_buf1})
	);
	fpu_bufrpt_grp32 i_inq_id_div_buf1 (
		.in ({5'h00,
			se_mul_buf4,
			arst_l_mul_buf2,
			inq_id[4:0],
			inq_op[7:0],
			inq_rnd_mode[1:0],
			inq_in1_50_0_neq_0,
			inq_in1_53_0_neq_0,
			inq_in1_53_32_neq_0,
			inq_in1_exp_eq_0,
			inq_in1_exp_neq_ffs,
			inq_in2_50_0_neq_0,
			inq_in2_53_0_neq_0,
			inq_in2_53_32_neq_0,
			inq_in2_exp_eq_0,
			inq_in2_exp_neq_ffs}),
		.out ({inq_id_div_buf1_unused[4:0],
			se_div_buf5,
			arst_l_in_buf3,
			inq_id_div_buf1[4:0],
			inq_op_div_buf1[7:0],
			inq_rnd_mode_div_buf1[1:0],
			inq_in1_50_0_neq_0_div_buf1,
			inq_in1_53_0_neq_0_div_buf1,
			inq_in1_53_32_neq_0_div_buf1,
			inq_in1_exp_eq_0_div_buf1,
			inq_in1_exp_neq_ffs_div_buf1,
			inq_in2_50_0_neq_0_div_buf1,
			inq_in2_53_0_neq_0_div_buf1,
			inq_in2_53_32_neq_0_div_buf1,
			inq_in2_exp_eq_0_div_buf1,
			inq_in2_exp_neq_ffs_div_buf1})
	);
	
	fpu_bufrpt_grp4 i_ctu_tst_buf1_hi (
		.in ({ctu_tst_short_chain,
			ctu_tst_macrotest,
			ctu_tst_scan_disable,
			ctu_tst_pre_grst_l}),
		.out ({ctu_tst_short_chain_buf1,
			ctu_tst_macrotest_buf1,
			ctu_tst_scan_disable_buf1,
			ctu_tst_pre_grst_l_buf1})
	);
	fpu_bufrpt_grp4 i_ctu_tst_buf1_lo (
		.in ({ctu_tst_scanmode,
			global_shift_enable,
			2'b00}),
		.out ({ctu_tst_scanmode_buf1,
			global_shift_enable_buf1,
			ctu_tst_buf1_lo_unused[1:0]})
	);
	
	fpu_bufrpt_grp4 i_cluster_cken_buf1 (
		.in ({cluster_cken,
			grst_l,
			2'b00}),
		.out ({cluster_cken_buf1,
			grst_l_buf1,
			cluster_cken_buf1_unused[1:0]})
	);
	
	fpu_bufrpt_grp4 i_se_buf1 (
		.in ({se,
			se,
			so_unbuf,
			1'b0}),
		.out ({se_add_buf1,
			se_mul64_buf1,
			so_buf1,
			se_buf1_unused})
	);
	fpu_bufrpt_grp4 i_se_add_buf2 (
		.in ({se_add_buf1,
			se_add_buf1,
			se_add_buf1,
			1'b0}),
		.out ({se_add_exp_buf2,
			se_add_frac_buf2,
			se_out_buf2,
			se_add_buf2_unused})
	);
	fpu_bufrpt_grp4 i_se_mul64_buf2 (
		.in ({se_mul64_buf1,
			se_mul64_buf1,
			2'b00}),
		.out ({se_mul64_buf2,
			se_cluster_header_buf2,
			se_mul64_buf2_unused[1:0]})
	);
	
	fpu_bufrpt_grp4 i_arst_l_buf1 (
		.in ({arst_l,
			3'b000}),
		.out ({arst_l_buf1,
			arst_l_buf1_unused[2:0]})
	);
	fpu_bufrpt_grp4 i_arst_l_buf2 (
		.in ({arst_l_buf1,
			arst_l_buf1,
			arst_l_buf1,
			fpu_grst_l}),
		.out ({arst_l_mul_buf2,
			arst_l_cluster_header_buf2,
			arst_l_div_buf2,
			fpu_grst_l_mul_buf1})
	);
	
	fpu_bufrpt_grp4 i_fdiv_clken_l_buf1 (
		.in ({fdiv_clken_l,
			fdiv_clken_l,
			2'b00}),
		.out ({fdiv_clken_l_div_exp_buf1,
			fdiv_clken_l_div_frac_buf1,
			fdiv_clken_l_buf1_unused[1:0]})
	);
	
	fpu_bufrpt_grp4 i_so_cluster_header_buf1 (
		.in ({scan_manual_6,
			3'b000}),
		.out ({scan_manual_6_buf1,
			so_cluster_header_buf1_unused[2:0]})
	);
	
	fpu_bufrpt_grp4 i_si_buf1 (
		.in ({si,
			3'b000}),
		.out ({si_buf1,
			si_buf1_unused[2:0]})
	);
	
	fpu_rptr_pcx_fpio_grp16 i_pcx_fpio_buf1_0 (
		.in ({pcx_fpio_data_px2[108],
			pcx_fpio_data_px2[109],
			pcx_fpio_data_px2[110],
			pcx_fpio_data_px2[111],
			pcx_fpio_data_px2[112],
			pcx_fpio_data_px2[113],
			pcx_fpio_data_px2[114],
			pcx_fpio_data_px2[115],
			pcx_fpio_data_px2[116],
			pcx_fpio_data_px2[117],
			pcx_fpio_data_px2[118],
			pcx_fpio_data_px2[119],
			pcx_fpio_data_px2[120],
			pcx_fpio_data_px2[121],
			pcx_fpio_data_px2[122],
			pcx_fpio_data_px2[123]}),
		.out ({pcx_fpio_data_px2_buf1[108],
			pcx_fpio_data_px2_buf1[109],
			pcx_fpio_data_px2_buf1[110],
			pcx_fpio_data_px2_buf1[111],
			pcx_fpio_data_px2_buf1[112],
			pcx_fpio_data_px2_buf1[113],
			pcx_fpio_data_px2_buf1[114],
			pcx_fpio_data_px2_buf1[115],
			pcx_fpio_data_px2_buf1[116],
			pcx_fpio_data_px2_buf1[117],
			pcx_fpio_data_px2_buf1[118],
			pcx_fpio_data_px2_buf1[119],
			pcx_fpio_data_px2_buf1[120],
			pcx_fpio_data_px2_buf1[121],
			pcx_fpio_data_px2_buf1[122],
			pcx_fpio_data_px2_buf1[123]})
	);
	fpu_rptr_pcx_fpio_grp16 i_pcx_fpio_buf1_1 (
		.in ({pcx_fpio_data_px2[92],
			pcx_fpio_data_px2[93],
			pcx_fpio_data_px2[94],
			pcx_fpio_data_px2[95],
			pcx_fpio_data_px2[96],
			pcx_fpio_data_px2[97],
			pcx_fpio_data_px2[98],
			pcx_fpio_data_px2[99],
			pcx_fpio_data_px2[100],
			pcx_fpio_data_px2[101],
			pcx_fpio_data_px2[102],
			pcx_fpio_data_px2[103],
			pcx_fpio_data_px2[104],
			pcx_fpio_data_px2[105],
			pcx_fpio_data_px2[106],
			pcx_fpio_data_px2[107]}),
		.out ({pcx_fpio_data_px2_buf1[92],
			pcx_fpio_data_px2_buf1[93],
			pcx_fpio_data_px2_buf1[94],
			pcx_fpio_data_px2_buf1[95],
			pcx_fpio_data_px2_buf1[96],
			pcx_fpio_data_px2_buf1[97],
			pcx_fpio_data_px2_buf1[98],
			pcx_fpio_data_px2_buf1[99],
			pcx_fpio_data_px2_buf1[100],
			pcx_fpio_data_px2_buf1[101],
			pcx_fpio_data_px2_buf1[102],
			pcx_fpio_data_px2_buf1[103],
			pcx_fpio_data_px2_buf1[104],
			pcx_fpio_data_px2_buf1[105],
			pcx_fpio_data_px2_buf1[106],
			pcx_fpio_data_px2_buf1[107]})
	);
	fpu_rptr_pcx_fpio_grp16 i_pcx_fpio_buf1_2 (
		.in ({pcx_fpio_data_px2[76],
			pcx_fpio_data_px2[77],
			pcx_fpio_data_px2[78],
			pcx_fpio_data_px2[79],
			pcx_fpio_data_px2[80],
			pcx_fpio_data_px2[81],
			pcx_fpio_data_px2[82],
			pcx_fpio_data_px2[83],
			pcx_fpio_data_px2[84],
			pcx_fpio_data_px2[85],
			pcx_fpio_data_px2[86],
			pcx_fpio_data_px2[87],
			pcx_fpio_data_px2[88],
			pcx_fpio_data_px2[89],
			pcx_fpio_data_px2[90],
			pcx_fpio_data_px2[91]}),
		.out ({pcx_fpio_data_px2_buf1[76],
			pcx_fpio_data_px2_buf1[77],
			pcx_fpio_data_px2_buf1[78],
			pcx_fpio_data_px2_buf1[79],
			pcx_fpio_data_px2_buf1[80],
			pcx_fpio_data_px2_buf1[81],
			pcx_fpio_data_px2_buf1[82],
			pcx_fpio_data_px2_buf1[83],
			pcx_fpio_data_px2_buf1[84],
			pcx_fpio_data_px2_buf1[85],
			pcx_fpio_data_px2_buf1[86],
			pcx_fpio_data_px2_buf1[87],
			pcx_fpio_data_px2_buf1[88],
			pcx_fpio_data_px2_buf1[89],
			pcx_fpio_data_px2_buf1[90],
			pcx_fpio_data_px2_buf1[91]})
	);
	fpu_rptr_pcx_fpio_grp16 i_pcx_fpio_buf1_3 (
		.in ({pcx_fpio_data_px2[3:0],
			pcx_fpio_data_px2[64],
			pcx_fpio_data_px2[65],
			pcx_fpio_data_px2[66],
			pcx_fpio_data_px2[67],
			pcx_fpio_data_px2[68],
			pcx_fpio_data_px2[69],
			pcx_fpio_data_px2[70],
			pcx_fpio_data_px2[71],
			pcx_fpio_data_px2[72],
			pcx_fpio_data_px2[73],
			pcx_fpio_data_px2[74],
			pcx_fpio_data_px2[75]}),
		.out ({pcx_fpio_data_px2_buf1[3:0],
			pcx_fpio_data_px2_buf1[64],
			pcx_fpio_data_px2_buf1[65],
			pcx_fpio_data_px2_buf1[66],
			pcx_fpio_data_px2_buf1[67],
			pcx_fpio_data_px2_buf1[68],
			pcx_fpio_data_px2_buf1[69],
			pcx_fpio_data_px2_buf1[70],
			pcx_fpio_data_px2_buf1[71],
			pcx_fpio_data_px2_buf1[72],
			pcx_fpio_data_px2_buf1[73],
			pcx_fpio_data_px2_buf1[74],
			pcx_fpio_data_px2_buf1[75]})
	);
	fpu_rptr_pcx_fpio_grp16 i_pcx_fpio_buf1_4 (
		.in (pcx_fpio_data_px2[19:4]),
		.out (pcx_fpio_data_px2_buf1[19:4])
	);
	fpu_rptr_pcx_fpio_grp16 i_pcx_fpio_buf1_5 (
		.in (pcx_fpio_data_px2[35:20]),
		.out (pcx_fpio_data_px2_buf1[35:20])
	);
	fpu_rptr_pcx_fpio_grp16 i_pcx_fpio_buf1_6 (
		.in ({pcx_fpio_data_rdy_px2,
			pcx_fpio_data_px2[50:36]}),
		.out ({pcx_fpio_data_rdy_px2_buf1,
			pcx_fpio_data_px2_buf1[50:36]})
	);
	fpu_rptr_pcx_fpio_grp16 i_pcx_fpio_buf1_7 (
		.in ({3'b000,
			pcx_fpio_data_px2[63:51]}),
		.out ({pcx_fpio_data_px2_buf1_unused[2:0],
			pcx_fpio_data_px2_buf1[63:51]})
	);
	
	fpu_rptr_fp_cpx_grp16 i_fp_cpx_buf1_0 (
		.in ({
			fp_cpx_data_ca[142],
			fp_cpx_data_ca[140],
			fp_cpx_data_ca[138],
			fp_cpx_data_ca[136],
			fp_cpx_data_ca[134],
			fp_cpx_data_ca[132],
			fp_cpx_data_ca[130],
			fp_cpx_data_ca[128],
			fp_cpx_req_cq[6],
			fp_cpx_req_cq[7],
			fp_cpx_req_cq[3],
			fp_cpx_req_cq[2],
			fp_cpx_req_cq[5],
			fp_cpx_req_cq[1],
			fp_cpx_req_cq[0],
			fp_cpx_req_cq[4]}),
		.out ({
			fp_cpx_data_ca_buf1[142],
			fp_cpx_data_ca_buf1[140],
			fp_cpx_data_ca_buf1[138],
			fp_cpx_data_ca_buf1[136],
			fp_cpx_data_ca_buf1[134],
			fp_cpx_data_ca_buf1[132],
			fp_cpx_data_ca_buf1[130],
			fp_cpx_data_ca_buf1[128],
			fp_cpx_req_cq_buf1[6],
			fp_cpx_req_cq_buf1[7],
			fp_cpx_req_cq_buf1[3],
			fp_cpx_req_cq_buf1[2],
			fp_cpx_req_cq_buf1[5],
			fp_cpx_req_cq_buf1[1],
			fp_cpx_req_cq_buf1[0],
			fp_cpx_req_cq_buf1[4]})
	);
	fpu_rptr_fp_cpx_grp16 i_fp_cpx_buf1_1 (
		.in ({
			fp_cpx_data_ca[34],
			fp_cpx_data_ca[36],
			fp_cpx_data_ca[38],
			fp_cpx_data_ca[40],
			fp_cpx_data_ca[42],
			fp_cpx_data_ca[44],
			fp_cpx_data_ca[46],
			fp_cpx_data_ca[48],
			fp_cpx_data_ca[50],
			fp_cpx_data_ca[52],
			fp_cpx_data_ca[54],
			fp_cpx_data_ca[56],
			fp_cpx_data_ca[58],
			fp_cpx_data_ca[60],
			fp_cpx_data_ca[62],
			fp_cpx_data_ca[144]}),
		.out ({
			fp_cpx_data_ca_buf1[34],
			fp_cpx_data_ca_buf1[36],
			fp_cpx_data_ca_buf1[38],
			fp_cpx_data_ca_buf1[40],
			fp_cpx_data_ca_buf1[42],
			fp_cpx_data_ca_buf1[44],
			fp_cpx_data_ca_buf1[46],
			fp_cpx_data_ca_buf1[48],
			fp_cpx_data_ca_buf1[50],
			fp_cpx_data_ca_buf1[52],
			fp_cpx_data_ca_buf1[54],
			fp_cpx_data_ca_buf1[56],
			fp_cpx_data_ca_buf1[58],
			fp_cpx_data_ca_buf1[60],
			fp_cpx_data_ca_buf1[62],
			fp_cpx_data_ca_buf1[144]})
	);
	fpu_rptr_fp_cpx_grp16 i_fp_cpx_buf1_2 (
		.in ({
			fp_cpx_data_ca[2],
			fp_cpx_data_ca[4],
			fp_cpx_data_ca[6],
			fp_cpx_data_ca[8],
			fp_cpx_data_ca[10],
			fp_cpx_data_ca[12],
			fp_cpx_data_ca[14],
			fp_cpx_data_ca[16],
			fp_cpx_data_ca[18],
			fp_cpx_data_ca[20],
			fp_cpx_data_ca[22],
			fp_cpx_data_ca[24],
			fp_cpx_data_ca[26],
			fp_cpx_data_ca[28],
			fp_cpx_data_ca[30],
			fp_cpx_data_ca[32]}),
		.out ({
			fp_cpx_data_ca_buf1[2],
			fp_cpx_data_ca_buf1[4],
			fp_cpx_data_ca_buf1[6],
			fp_cpx_data_ca_buf1[8],
			fp_cpx_data_ca_buf1[10],
			fp_cpx_data_ca_buf1[12],
			fp_cpx_data_ca_buf1[14],
			fp_cpx_data_ca_buf1[16],
			fp_cpx_data_ca_buf1[18],
			fp_cpx_data_ca_buf1[20],
			fp_cpx_data_ca_buf1[22],
			fp_cpx_data_ca_buf1[24],
			fp_cpx_data_ca_buf1[26],
			fp_cpx_data_ca_buf1[28],
			fp_cpx_data_ca_buf1[30],
			fp_cpx_data_ca_buf1[32]})
	);
	fpu_rptr_fp_cpx_grp16 i_fp_cpx_buf1_3 (
		.in ({
			fp_cpx_data_ca[31],
			fp_cpx_data_ca[27],
			fp_cpx_data_ca[23],
			fp_cpx_data_ca[25],
			fp_cpx_data_ca[21],
			fp_cpx_data_ca[17],
			fp_cpx_data_ca[19],
			fp_cpx_data_ca[15],
			fp_cpx_data_ca[11],
			fp_cpx_data_ca[13],
			fp_cpx_data_ca[9],
			fp_cpx_data_ca[5],
			fp_cpx_data_ca[7],
			fp_cpx_data_ca[3],
			fp_cpx_data_ca[0],
			fp_cpx_data_ca[1]}),
		.out ({
			fp_cpx_data_ca_buf1[31],
			fp_cpx_data_ca_buf1[27],
			fp_cpx_data_ca_buf1[23],
			fp_cpx_data_ca_buf1[25],
			fp_cpx_data_ca_buf1[21],
			fp_cpx_data_ca_buf1[17],
			fp_cpx_data_ca_buf1[19],
			fp_cpx_data_ca_buf1[15],
			fp_cpx_data_ca_buf1[11],
			fp_cpx_data_ca_buf1[13],
			fp_cpx_data_ca_buf1[9],
			fp_cpx_data_ca_buf1[5],
			fp_cpx_data_ca_buf1[7],
			fp_cpx_data_ca_buf1[3],
			fp_cpx_data_ca_buf1[0],
			fp_cpx_data_ca_buf1[1]})
	);
	fpu_rptr_fp_cpx_grp16 i_fp_cpx_buf1_4 (
		.in ({
			fp_cpx_data_ca[59],
			fp_cpx_data_ca[61],
			fp_cpx_data_ca[57],
			fp_cpx_data_ca[53],
			fp_cpx_data_ca[55],
			fp_cpx_data_ca[51],
			fp_cpx_data_ca[47],
			fp_cpx_data_ca[49],
			fp_cpx_data_ca[45],
			fp_cpx_data_ca[41],
			fp_cpx_data_ca[43],
			fp_cpx_data_ca[39],
			fp_cpx_data_ca[35],
			fp_cpx_data_ca[37],
			fp_cpx_data_ca[33],
			fp_cpx_data_ca[29]}),
		.out ({
			fp_cpx_data_ca_buf1[59],
			fp_cpx_data_ca_buf1[61],
			fp_cpx_data_ca_buf1[57],
			fp_cpx_data_ca_buf1[53],
			fp_cpx_data_ca_buf1[55],
			fp_cpx_data_ca_buf1[51],
			fp_cpx_data_ca_buf1[47],
			fp_cpx_data_ca_buf1[49],
			fp_cpx_data_ca_buf1[45],
			fp_cpx_data_ca_buf1[41],
			fp_cpx_data_ca_buf1[43],
			fp_cpx_data_ca_buf1[39],
			fp_cpx_data_ca_buf1[35],
			fp_cpx_data_ca_buf1[37],
			fp_cpx_data_ca_buf1[33],
			fp_cpx_data_ca_buf1[29]})
	);
	fpu_rptr_fp_cpx_grp16 i_fp_cpx_buf1_5 (
		.in ({
			fp_cpx_data_ca[113],
			fp_cpx_data_ca[117],
			fp_cpx_data_ca[121],
			fp_cpx_data_ca[119],
			fp_cpx_data_ca[123],
			fp_cpx_data_ca[127],
			fp_cpx_data_ca[125],
			fp_cpx_data_ca[129],
			fp_cpx_data_ca[133],
			fp_cpx_data_ca[131],
			fp_cpx_data_ca[135],
			fp_cpx_data_ca[139],
			fp_cpx_data_ca[137],
			fp_cpx_data_ca[141],
			fp_cpx_data_ca[143],
			fp_cpx_data_ca[63]}),
		.out ({
			fp_cpx_data_ca_buf1[113],
			fp_cpx_data_ca_buf1[117],
			fp_cpx_data_ca_buf1[121],
			fp_cpx_data_ca_buf1[119],
			fp_cpx_data_ca_buf1[123],
			fp_cpx_data_ca_buf1[127],
			fp_cpx_data_ca_buf1[125],
			fp_cpx_data_ca_buf1[129],
			fp_cpx_data_ca_buf1[133],
			fp_cpx_data_ca_buf1[131],
			fp_cpx_data_ca_buf1[135],
			fp_cpx_data_ca_buf1[139],
			fp_cpx_data_ca_buf1[137],
			fp_cpx_data_ca_buf1[141],
			fp_cpx_data_ca_buf1[143],
			fp_cpx_data_ca_buf1[63]})
	);
	fpu_rptr_fp_cpx_grp16 i_fp_cpx_buf1_6 (
		.in ({
			fp_cpx_data_ca[85],
			fp_cpx_data_ca[83],
			fp_cpx_data_ca[87],
			fp_cpx_data_ca[91],
			fp_cpx_data_ca[89],
			fp_cpx_data_ca[93],
			fp_cpx_data_ca[97],
			fp_cpx_data_ca[95],
			fp_cpx_data_ca[99],
			fp_cpx_data_ca[103],
			fp_cpx_data_ca[101],
			fp_cpx_data_ca[105],
			fp_cpx_data_ca[109],
			fp_cpx_data_ca[107],
			fp_cpx_data_ca[111],
			fp_cpx_data_ca[115]}),
		.out ({
			fp_cpx_data_ca_buf1[85],
			fp_cpx_data_ca_buf1[83],
			fp_cpx_data_ca_buf1[87],
			fp_cpx_data_ca_buf1[91],
			fp_cpx_data_ca_buf1[89],
			fp_cpx_data_ca_buf1[93],
			fp_cpx_data_ca_buf1[97],
			fp_cpx_data_ca_buf1[95],
			fp_cpx_data_ca_buf1[99],
			fp_cpx_data_ca_buf1[103],
			fp_cpx_data_ca_buf1[101],
			fp_cpx_data_ca_buf1[105],
			fp_cpx_data_ca_buf1[109],
			fp_cpx_data_ca_buf1[107],
			fp_cpx_data_ca_buf1[111],
			fp_cpx_data_ca_buf1[115]})
	);
	fpu_rptr_fp_cpx_grp16 i_fp_cpx_buf1_7 (
		.in ({
			fp_cpx_data_ca[114],
			fp_cpx_data_ca[116],
			fp_cpx_data_ca[118],
			fp_cpx_data_ca[120],
			fp_cpx_data_ca[122],
			fp_cpx_data_ca[124],
			fp_cpx_data_ca[126],
			fp_cpx_data_ca[65],
			fp_cpx_data_ca[67],
			fp_cpx_data_ca[69],
			fp_cpx_data_ca[73],
			fp_cpx_data_ca[71],
			fp_cpx_data_ca[75],
			fp_cpx_data_ca[79],
			fp_cpx_data_ca[77],
			fp_cpx_data_ca[81]}),
		.out ({
			fp_cpx_data_ca_buf1[114],
			fp_cpx_data_ca_buf1[116],
			fp_cpx_data_ca_buf1[118],
			fp_cpx_data_ca_buf1[120],
			fp_cpx_data_ca_buf1[122],
			fp_cpx_data_ca_buf1[124],
			fp_cpx_data_ca_buf1[126],
			fp_cpx_data_ca_buf1[65],
			fp_cpx_data_ca_buf1[67],
			fp_cpx_data_ca_buf1[69],
			fp_cpx_data_ca_buf1[73],
			fp_cpx_data_ca_buf1[71],
			fp_cpx_data_ca_buf1[75],
			fp_cpx_data_ca_buf1[79],
			fp_cpx_data_ca_buf1[77],
			fp_cpx_data_ca_buf1[81]})
	);
	fpu_rptr_fp_cpx_grp16 i_fp_cpx_buf1_8 (
		.in ({
			fp_cpx_data_ca[82],
			fp_cpx_data_ca[84],
			fp_cpx_data_ca[86],
			fp_cpx_data_ca[88],
			fp_cpx_data_ca[90],
			fp_cpx_data_ca[92],
			fp_cpx_data_ca[94],
			fp_cpx_data_ca[96],
			fp_cpx_data_ca[98],
			fp_cpx_data_ca[100],
			fp_cpx_data_ca[102],
			fp_cpx_data_ca[104],
			fp_cpx_data_ca[106],
			fp_cpx_data_ca[108],
			fp_cpx_data_ca[110],
			fp_cpx_data_ca[112]}),
		.out ({
			fp_cpx_data_ca_buf1[82],
			fp_cpx_data_ca_buf1[84],
			fp_cpx_data_ca_buf1[86],
			fp_cpx_data_ca_buf1[88],
			fp_cpx_data_ca_buf1[90],
			fp_cpx_data_ca_buf1[92],
			fp_cpx_data_ca_buf1[94],
			fp_cpx_data_ca_buf1[96],
			fp_cpx_data_ca_buf1[98],
			fp_cpx_data_ca_buf1[100],
			fp_cpx_data_ca_buf1[102],
			fp_cpx_data_ca_buf1[104],
			fp_cpx_data_ca_buf1[106],
			fp_cpx_data_ca_buf1[108],
			fp_cpx_data_ca_buf1[110],
			fp_cpx_data_ca_buf1[112]})
	);
	fpu_rptr_fp_cpx_grp16 i_fp_cpx_buf1_9 (
		.in ({
			6'b000000,
			so_buf1,
			fp_cpx_data_ca[64],
			fp_cpx_data_ca[66],
			fp_cpx_data_ca[68],
			fp_cpx_data_ca[70],
			fp_cpx_data_ca[72],
			fp_cpx_data_ca[74],
			fp_cpx_data_ca[76],
			fp_cpx_data_ca[78],
			fp_cpx_data_ca[80]}),
		.out ({
			fp_cpx_buf1_9_unused[5:0],
			so,
			fp_cpx_data_ca_buf1[64],
			fp_cpx_data_ca_buf1[66],
			fp_cpx_data_ca_buf1[68],
			fp_cpx_data_ca_buf1[70],
			fp_cpx_data_ca_buf1[72],
			fp_cpx_data_ca_buf1[74],
			fp_cpx_data_ca_buf1[76],
			fp_cpx_data_ca_buf1[78],
			fp_cpx_data_ca_buf1[80]})
	);
	
	fpu_rptr_inq i_inq_sram_din_buf1 (
		.in (inq_sram_din_unbuf[155:0]),
		.out (inq_sram_din_buf1[155:0])
	);
endmodule
module fpu_bufrpt_grp4 (
	in,
	out
);
	
	input [3:0] in;
	output [3:0] out;
	assign out[3:0] = in[3:0];
endmodule
module fpu_rptr_fp_cpx_grp16 (
	in,
	out
);
	input [15:0] in;
	output [15:0] out;
	assign out[15:0] = in[15:0];
endmodule
module fpu_rptr_pcx_fpio_grp16 (
	in,
	out
);
	input [15:0] in;
	output [15:0] out;
	assign out[15:0] = in[15:0];
endmodule
module fpu_rptr_inq (
	in,
	out
);
	
	input [155:0] in;
	output [155:0] out;
	assign out[155:0] = in[155:0];
endmodule
module io_xbar_top_wrap
(
    input clk,
    input reset_in,
    
    input [64-1:0] dataIn_0,
    input [64-1:0] dataIn_1,
    input [64-1:0] dataIn_2,
    input [64-1:0] dataIn_3,
    input [64-1:0] dataIn_4,
    input [64-1:0] dataIn_5,
    input validIn_0,
    input validIn_1,
    input validIn_2,
    input validIn_3,
    input validIn_4,
    input validIn_5,
    input yummyIn_0,
    input yummyIn_1,
    input yummyIn_2,
    input yummyIn_3,
    input yummyIn_4,
    input yummyIn_5,
       
    input [8-1:0] myLocX,       
    input [8-1:0] myLocY,
    input [14-1:0] myChipID,
    
    output [64-1:0] dataOut_0,
    output [64-1:0] dataOut_1,
    output [64-1:0] dataOut_2,
    output [64-1:0] dataOut_3,
    output [64-1:0] dataOut_4,
    output [64-1:0] dataOut_5,
    output validOut_0,
    output validOut_1,
    output validOut_2,
    output validOut_3,
    output validOut_4,
    output validOut_5,
    output yummyOut_0,
    output yummyOut_1,
    output yummyOut_2,
    output yummyOut_3,
    output yummyOut_4,
    output yummyOut_5,
    
    
    output thanksIn_5      
);
    io_xbar_top io_xbar_top
    (
        .clk(clk),
        .reset_in(reset_in),
        
        .dataIn_0(dataIn_0),
        .dataIn_1(dataIn_1),
        .dataIn_2(dataIn_2),
        .dataIn_3(dataIn_3),
        .dataIn_4(dataIn_4),
        .dataIn_5(dataIn_5),
        .validIn_0(validIn_0),
        .validIn_1(validIn_1),
        .validIn_2(validIn_2),
        .validIn_3(validIn_3),
        .validIn_4(validIn_4),
        .validIn_5(validIn_5),
        .yummyIn_0(yummyIn_0),
        .yummyIn_1(yummyIn_1),
        .yummyIn_2(yummyIn_2),
        .yummyIn_3(yummyIn_3),
        .yummyIn_4(yummyIn_4),
        .yummyIn_5(yummyIn_5),
        .myLocX(myLocX),
        .myLocY(myLocY),
        .myChipID(myChipID),
        .ec_cfg(24'b0),
        .store_meter_partner_address_X(5'b0),
        .store_meter_partner_address_Y(5'b0),
        
        .dataOut_0(dataOut_0),
        .dataOut_1(dataOut_1),
        .dataOut_2(dataOut_2),
        .dataOut_3(dataOut_3),
        .dataOut_4(dataOut_4),
        .dataOut_5(dataOut_5),
        .validOut_0(validOut_0),
        .validOut_1(validOut_1),
        .validOut_2(validOut_2),
        .validOut_3(validOut_3),
        .validOut_4(validOut_4),
        .validOut_5(validOut_5),
        .yummyOut_0(yummyOut_0),
        .yummyOut_1(yummyOut_1),
        .yummyOut_2(yummyOut_2),
        .yummyOut_3(yummyOut_3),
        .yummyOut_4(yummyOut_4),
        .yummyOut_5(yummyOut_5),
        .thanksIn_5(thanksIn_5),
        .external_interrupt(),
        .store_meter_ack_partner(),
        .store_meter_ack_non_partner(),
        .ec_out()
    ); 
endmodule
module io_xbar_top(clk,
		    reset_in,
        dataIn_0, dataIn_1, dataIn_2, dataIn_3, dataIn_4, dataIn_5, 
        validIn_0, validIn_1, validIn_2, validIn_3, validIn_4, validIn_5, 
        yummyIn_0,yummyIn_1,yummyIn_2,yummyIn_3,yummyIn_4,yummyIn_5,
		    myLocX,
		    myLocY,
            myChipID,
		    store_meter_partner_address_X,
		    store_meter_partner_address_Y,
		    ec_cfg,
        dataOut_0, dataOut_1, dataOut_2, dataOut_3, dataOut_4, dataOut_5, 
        validOut_0, validOut_1, validOut_2, validOut_3, validOut_4, validOut_5, 
        yummyOut_0,yummyOut_1,yummyOut_2,yummyOut_3,yummyOut_4,yummyOut_5,
		    thanksIn_5,
		    external_interrupt,
		    store_meter_ack_partner,
		    store_meter_ack_non_partner,
		    ec_out);
input clk;
input reset_in;
input [64-1:0] dataIn_0;
input [64-1:0] dataIn_1;
input [64-1:0] dataIn_2;
input [64-1:0] dataIn_3;
input [64-1:0] dataIn_4;
input [64-1:0] dataIn_5;
input validIn_0;
input validIn_1;
input validIn_2;
input validIn_3;
input validIn_4;
input validIn_5;
input yummyIn_0;
input yummyIn_1;
input yummyIn_2;
input yummyIn_3;
input yummyIn_4;
input yummyIn_5;
   
input [8-1:0] myLocX;		
input [8-1:0] myLocY;
input [14-1:0] myChipID;
input [4:0] store_meter_partner_address_X;
input [4:0] store_meter_partner_address_Y;
input [23:0] ec_cfg;            
output [64-1:0] dataOut_0;
output [64-1:0] dataOut_1;
output [64-1:0] dataOut_2;
output [64-1:0] dataOut_3;
output [64-1:0] dataOut_4;
output [64-1:0] dataOut_5;
output validOut_0;
output validOut_1;
output validOut_2;
output validOut_3;
output validOut_4;
output validOut_5;
output yummyOut_0;
output yummyOut_1;
output yummyOut_2;
output yummyOut_3;
output yummyOut_4;
output yummyOut_5;
output thanksIn_5;		
output external_interrupt;	
				
output store_meter_ack_partner;      
                                     
output store_meter_ack_non_partner;  
                                     
output [5:0] ec_out;
wire   ec_wants_to_send_but_cannot_0;
wire   ec_wants_to_send_but_cannot_1;
wire   ec_wants_to_send_but_cannot_2;
wire   ec_wants_to_send_but_cannot_3;
wire   ec_wants_to_send_but_cannot_4;
wire   ec_wants_to_send_but_cannot_5;
   wire store_ack_received;
   wire store_ack_received_r;
   wire [9:0] store_ack_addr;
   wire [9:0] store_ack_addr_r;
wire node_0_input_tail;
wire node_1_input_tail;
wire node_2_input_tail;
wire node_3_input_tail;
wire node_4_input_tail;
wire node_5_input_tail;
wire [64-1:0] node_0_input_data;
wire [64-1:0] node_1_input_data;
wire [64-1:0] node_2_input_data;
wire [64-1:0] node_3_input_data;
wire [64-1:0] node_4_input_data;
wire [64-1:0] node_5_input_data;
wire node_0_input_valid;
wire node_1_input_valid;
wire node_2_input_valid;
wire node_3_input_valid;
wire node_4_input_valid;
wire node_5_input_valid;
wire thanks_0_to_0;
wire thanks_0_to_1;
wire thanks_0_to_2;
wire thanks_0_to_3;
wire thanks_0_to_4;
wire thanks_0_to_5;
wire thanks_1_to_0;
wire thanks_1_to_1;
wire thanks_1_to_2;
wire thanks_1_to_3;
wire thanks_1_to_4;
wire thanks_1_to_5;
wire thanks_2_to_0;
wire thanks_2_to_1;
wire thanks_2_to_2;
wire thanks_2_to_3;
wire thanks_2_to_4;
wire thanks_2_to_5;
wire thanks_3_to_0;
wire thanks_3_to_1;
wire thanks_3_to_2;
wire thanks_3_to_3;
wire thanks_3_to_4;
wire thanks_3_to_5;
wire thanks_4_to_0;
wire thanks_4_to_1;
wire thanks_4_to_2;
wire thanks_4_to_3;
wire thanks_4_to_4;
wire thanks_4_to_5;
wire thanks_5_to_0;
wire thanks_5_to_1;
wire thanks_5_to_2;
wire thanks_5_to_3;
wire thanks_5_to_4;
wire thanks_5_to_5;
wire route_req_0_to_0;
wire route_req_0_to_1;
wire route_req_0_to_2;
wire route_req_0_to_3;
wire route_req_0_to_4;
wire route_req_0_to_5;
wire route_req_1_to_0;
wire route_req_1_to_1;
wire route_req_1_to_2;
wire route_req_1_to_3;
wire route_req_1_to_4;
wire route_req_1_to_5;
wire route_req_2_to_0;
wire route_req_2_to_1;
wire route_req_2_to_2;
wire route_req_2_to_3;
wire route_req_2_to_4;
wire route_req_2_to_5;
wire route_req_3_to_0;
wire route_req_3_to_1;
wire route_req_3_to_2;
wire route_req_3_to_3;
wire route_req_3_to_4;
wire route_req_3_to_5;
wire route_req_4_to_0;
wire route_req_4_to_1;
wire route_req_4_to_2;
wire route_req_4_to_3;
wire route_req_4_to_4;
wire route_req_4_to_5;
wire route_req_5_to_0;
wire route_req_5_to_1;
wire route_req_5_to_2;
wire route_req_5_to_3;
wire route_req_5_to_4;
wire route_req_5_to_5;
wire default_ready_2_to_0;
wire default_ready_3_to_1;
wire default_ready_4_to_2;
wire default_ready_0_to_3;
wire default_ready_1_to_4;
wire default_ready_2_to_5;
wire yummyOut_0_internal;
wire yummyOut_1_internal;
wire yummyOut_2_internal;
wire yummyOut_3_internal;
wire yummyOut_4_internal;
wire yummyOut_5_internal;
wire validOut_0_internal;
wire validOut_1_internal;
wire validOut_2_internal;
wire validOut_3_internal;
wire validOut_4_internal;
wire validOut_5_internal;
wire [64-1:0] dataOut_0_internal;
wire [64-1:0] dataOut_1_internal;
wire [64-1:0] dataOut_2_internal;
wire [64-1:0] dataOut_3_internal;
wire [64-1:0] dataOut_4_internal;
wire [64-1:0] dataOut_5_internal;
wire yummyOut_0_flip1_out;
wire yummyOut_1_flip1_out;
wire yummyOut_2_flip1_out;
wire yummyOut_3_flip1_out;
wire yummyOut_4_flip1_out;
wire validOut_0_flip1_out;
wire validOut_1_flip1_out;
wire validOut_2_flip1_out;
wire validOut_3_flip1_out;
wire validOut_4_flip1_out;
wire [64-1:0] dataOut_0_flip1_out;
wire [64-1:0] dataOut_1_flip1_out;
wire [64-1:0] dataOut_2_flip1_out;
wire [64-1:0] dataOut_3_flip1_out;
wire [64-1:0] dataOut_4_flip1_out;
wire yummyIn_0_internal;
wire yummyIn_1_internal;
wire yummyIn_2_internal;
wire yummyIn_3_internal;
wire yummyIn_4_internal;
wire yummyIn_5_internal;
wire validIn_0_internal;
wire validIn_1_internal;
wire validIn_2_internal;
wire validIn_3_internal;
wire validIn_4_internal;
wire [64-1:0] dataIn_0_internal;
wire [64-1:0] dataIn_1_internal;
wire [64-1:0] dataIn_2_internal;
wire [64-1:0] dataIn_3_internal;
wire [64-1:0] dataIn_4_internal;
wire yummyIn_0_flip1_out;
wire yummyIn_1_flip1_out;
wire yummyIn_2_flip1_out;
wire yummyIn_3_flip1_out;
wire yummyIn_4_flip1_out;
wire validIn_0_flip1_out;
wire validIn_1_flip1_out;
wire validIn_2_flip1_out;
wire validIn_3_flip1_out;
wire validIn_4_flip1_out;
wire [64-1:0] dataIn_0_flip1_out;
wire [64-1:0] dataIn_1_flip1_out;
wire [64-1:0] dataIn_2_flip1_out;
wire [64-1:0] dataIn_3_flip1_out;
wire [64-1:0] dataIn_4_flip1_out;
reg [8-1:0] myLocX_f;
reg [8-1:0] myLocY_f;
reg [14-1:0] myChipID_f;
wire   reset;
reg ec_thanks_0_to_0_reg, ec_thanks_0_to_1_reg, ec_thanks_0_to_2_reg, ec_thanks_0_to_3_reg, ec_thanks_0_to_4_reg, ec_thanks_0_to_5_reg;
reg ec_thanks_1_to_0_reg, ec_thanks_1_to_1_reg, ec_thanks_1_to_2_reg, ec_thanks_1_to_3_reg, ec_thanks_1_to_4_reg, ec_thanks_1_to_5_reg;
reg ec_thanks_2_to_0_reg, ec_thanks_2_to_1_reg, ec_thanks_2_to_2_reg, ec_thanks_2_to_3_reg, ec_thanks_2_to_4_reg, ec_thanks_2_to_5_reg;
reg ec_thanks_3_to_0_reg, ec_thanks_3_to_1_reg, ec_thanks_3_to_2_reg, ec_thanks_3_to_3_reg, ec_thanks_3_to_4_reg, ec_thanks_3_to_5_reg;
reg ec_thanks_4_to_0_reg, ec_thanks_4_to_1_reg, ec_thanks_4_to_2_reg, ec_thanks_4_to_3_reg, ec_thanks_4_to_4_reg, ec_thanks_4_to_5_reg;
reg ec_thanks_5_to_0_reg, ec_thanks_5_to_1_reg, ec_thanks_5_to_2_reg, ec_thanks_5_to_3_reg, ec_thanks_5_to_4_reg, ec_thanks_5_to_5_reg;
reg ec_wants_to_send_but_cannot_0_reg, ec_wants_to_send_but_cannot_1_reg, ec_wants_to_send_but_cannot_2_reg, ec_wants_to_send_but_cannot_3_reg, ec_wants_to_send_but_cannot_4_reg, ec_wants_to_send_but_cannot_5_reg;
reg ec_0_input_valid_reg, ec_1_input_valid_reg, ec_2_input_valid_reg, ec_3_input_valid_reg, ec_4_input_valid_reg, ec_5_input_valid_reg;
always @(posedge clk)
  begin
    
    ec_thanks_0_to_0_reg <= thanks_0_to_0; ec_thanks_0_to_1_reg <= thanks_0_to_1; ec_thanks_0_to_2_reg <= thanks_0_to_2; ec_thanks_0_to_3_reg <= thanks_0_to_3; ec_thanks_0_to_4_reg <= thanks_0_to_4; ec_thanks_0_to_5_reg <= thanks_0_to_5;
    ec_thanks_1_to_0_reg <= thanks_1_to_0; ec_thanks_1_to_1_reg <= thanks_1_to_1; ec_thanks_1_to_2_reg <= thanks_1_to_2; ec_thanks_1_to_3_reg <= thanks_1_to_3; ec_thanks_1_to_4_reg <= thanks_1_to_4; ec_thanks_1_to_5_reg <= thanks_1_to_5;
    ec_thanks_2_to_0_reg <= thanks_2_to_0; ec_thanks_2_to_1_reg <= thanks_2_to_1; ec_thanks_2_to_2_reg <= thanks_2_to_2; ec_thanks_2_to_3_reg <= thanks_2_to_3; ec_thanks_2_to_4_reg <= thanks_2_to_4; ec_thanks_2_to_5_reg <= thanks_2_to_5;
    ec_thanks_3_to_0_reg <= thanks_3_to_0; ec_thanks_3_to_1_reg <= thanks_3_to_1; ec_thanks_3_to_2_reg <= thanks_3_to_2; ec_thanks_3_to_3_reg <= thanks_3_to_3; ec_thanks_3_to_4_reg <= thanks_3_to_4; ec_thanks_3_to_5_reg <= thanks_3_to_5;
    ec_thanks_4_to_0_reg <= thanks_4_to_0; ec_thanks_4_to_1_reg <= thanks_4_to_1; ec_thanks_4_to_2_reg <= thanks_4_to_2; ec_thanks_4_to_3_reg <= thanks_4_to_3; ec_thanks_4_to_4_reg <= thanks_4_to_4; ec_thanks_4_to_5_reg <= thanks_4_to_5;
    ec_thanks_5_to_0_reg <= thanks_5_to_0; ec_thanks_5_to_1_reg <= thanks_5_to_1; ec_thanks_5_to_2_reg <= thanks_5_to_2; ec_thanks_5_to_3_reg <= thanks_5_to_3; ec_thanks_5_to_4_reg <= thanks_5_to_4; ec_thanks_5_to_5_reg <= thanks_5_to_5;
    ec_wants_to_send_but_cannot_0_reg <= ec_wants_to_send_but_cannot_0;
    ec_wants_to_send_but_cannot_1_reg <= ec_wants_to_send_but_cannot_1;
    ec_wants_to_send_but_cannot_2_reg <= ec_wants_to_send_but_cannot_2;
    ec_wants_to_send_but_cannot_3_reg <= ec_wants_to_send_but_cannot_3;
    ec_wants_to_send_but_cannot_4_reg <= ec_wants_to_send_but_cannot_4;
    ec_wants_to_send_but_cannot_5_reg <= ec_wants_to_send_but_cannot_5;
    ec_0_input_valid_reg <= node_0_input_valid;
    ec_1_input_valid_reg <= node_1_input_valid;
    ec_2_input_valid_reg <= node_2_input_valid;
    ec_3_input_valid_reg <= node_3_input_valid;
    ec_4_input_valid_reg <= node_4_input_valid;
    ec_5_input_valid_reg <= node_5_input_valid;
    
  end
wire ec_thanks_to_0= ec_thanks_0_to_0_reg | ec_thanks_1_to_0_reg | ec_thanks_2_to_0_reg | ec_thanks_3_to_0_reg | ec_thanks_4_to_0_reg | ec_thanks_5_to_0_reg ;
wire ec_thanks_to_1= ec_thanks_0_to_1_reg | ec_thanks_1_to_1_reg | ec_thanks_2_to_1_reg | ec_thanks_3_to_1_reg | ec_thanks_4_to_1_reg | ec_thanks_5_to_1_reg ;
wire ec_thanks_to_2= ec_thanks_0_to_2_reg | ec_thanks_1_to_2_reg | ec_thanks_2_to_2_reg | ec_thanks_3_to_2_reg | ec_thanks_4_to_2_reg | ec_thanks_5_to_2_reg ;
wire ec_thanks_to_3= ec_thanks_0_to_3_reg | ec_thanks_1_to_3_reg | ec_thanks_2_to_3_reg | ec_thanks_3_to_3_reg | ec_thanks_4_to_3_reg | ec_thanks_5_to_3_reg ;
wire ec_thanks_to_4= ec_thanks_0_to_4_reg | ec_thanks_1_to_4_reg | ec_thanks_2_to_4_reg | ec_thanks_3_to_4_reg | ec_thanks_4_to_4_reg | ec_thanks_5_to_4_reg ;
wire ec_thanks_to_5= ec_thanks_0_to_5_reg | ec_thanks_1_to_5_reg | ec_thanks_2_to_5_reg | ec_thanks_3_to_5_reg | ec_thanks_4_to_5_reg | ec_thanks_5_to_5_reg ;
io_xbar_one_of_n_plus_3 #(1) ec_mux_0(.in0(ec_wants_to_send_but_cannot_0),
                        .in1(ec_thanks_5_to_0_reg),
                        .in2(ec_thanks_4_to_0_reg),
                        .in3(ec_thanks_3_to_0_reg),
                        .in4(ec_thanks_2_to_0_reg),
                        .in5(ec_thanks_1_to_0_reg),
                        .in6(ec_thanks_0_to_0_reg),
                        .in7(ec_thanks_to_0),
                        .in8(ec_0_input_valid_reg & ~ec_thanks_to_0),
                        .sel(ec_cfg[23:20]),
                        .out(ec_out[5]));
io_xbar_one_of_n_plus_3 #(1) ec_mux_1(.in0(ec_wants_to_send_but_cannot_1),
                        .in1(ec_thanks_5_to_1_reg),
                        .in2(ec_thanks_4_to_1_reg),
                        .in3(ec_thanks_3_to_1_reg),
                        .in4(ec_thanks_2_to_1_reg),
                        .in5(ec_thanks_1_to_1_reg),
                        .in6(ec_thanks_0_to_1_reg),
                        .in7(ec_thanks_to_1),
                        .in8(ec_1_input_valid_reg & ~ec_thanks_to_1),
                        .sel(ec_cfg[19:16]),
                        .out(ec_out[4]));
io_xbar_one_of_n_plus_3 #(1) ec_mux_2(.in0(ec_wants_to_send_but_cannot_2),
                        .in1(ec_thanks_5_to_2_reg),
                        .in2(ec_thanks_4_to_2_reg),
                        .in3(ec_thanks_3_to_2_reg),
                        .in4(ec_thanks_2_to_2_reg),
                        .in5(ec_thanks_1_to_2_reg),
                        .in6(ec_thanks_0_to_2_reg),
                        .in7(ec_thanks_to_2),
                        .in8(ec_2_input_valid_reg & ~ec_thanks_to_2),
                        .sel(ec_cfg[15:12]),
                        .out(ec_out[3]));
io_xbar_one_of_n_plus_3 #(1) ec_mux_3(.in0(ec_wants_to_send_but_cannot_3),
                        .in1(ec_thanks_5_to_3_reg),
                        .in2(ec_thanks_4_to_3_reg),
                        .in3(ec_thanks_3_to_3_reg),
                        .in4(ec_thanks_2_to_3_reg),
                        .in5(ec_thanks_1_to_3_reg),
                        .in6(ec_thanks_0_to_3_reg),
                        .in7(ec_thanks_to_3),
                        .in8(ec_3_input_valid_reg & ~ec_thanks_to_3),
                        .sel(ec_cfg[11:8]),
                        .out(ec_out[2]));
io_xbar_one_of_n_plus_3 #(1) ec_mux_4(.in0(ec_wants_to_send_but_cannot_4),
                        .in1(ec_thanks_5_to_4_reg),
                        .in2(ec_thanks_4_to_4_reg),
                        .in3(ec_thanks_3_to_4_reg),
                        .in4(ec_thanks_2_to_4_reg),
                        .in5(ec_thanks_1_to_4_reg),
                        .in6(ec_thanks_0_to_4_reg),
                        .in7(ec_thanks_to_4),
                        .in8(ec_4_input_valid_reg & ~ec_thanks_to_4),
                        .sel(ec_cfg[7:4]),
                        .out(ec_out[1]));
io_xbar_one_of_n_plus_3 #(1) ec_mux_5(.in0(ec_wants_to_send_but_cannot_5),
                        .in1(ec_thanks_5_to_5_reg),
                        .in2(ec_thanks_4_to_5_reg),
                        .in3(ec_thanks_3_to_5_reg),
                        .in4(ec_thanks_2_to_5_reg),
                        .in5(ec_thanks_1_to_5_reg),
                        .in6(ec_thanks_0_to_5_reg),
                        .in7(ec_thanks_to_5),
                        .in8(ec_5_input_valid_reg & ~ec_thanks_to_5),
                        .sel(ec_cfg[3:0]),
                        .out(ec_out[0]));
io_xbar_net_dff #(1) REG_reset_fin(.d(reset_in), .q(reset), .clk(clk));
io_xbar_net_dff #(10) REG_store_ack_addr(   .d(store_ack_addr),     .q(store_ack_addr_r),     .clk(clk));
io_xbar_net_dff #(1) REG_store_ack_received(.d(store_ack_received), .q(store_ack_received_r), .clk(clk));
   wire is_partner_address_v_r;
   io_xbar_bus_compare_equal #(10) CMP_partner_address (.a(store_ack_addr_r),
                                        .b({ store_meter_partner_address_Y, store_meter_partner_address_X } ),
                                        .bus_equal(is_partner_address_v_r));
   assign store_meter_ack_partner     = is_partner_address_v_r & store_ack_received_r;
   assign store_meter_ack_non_partner = ~is_partner_address_v_r & store_ack_received_r;
always @ (posedge clk)
begin
        if(reset)
        begin
                myLocY_f <= 8'd0;
                myLocX_f <= 8'd0;
                myChipID_f <= 14'd0;
        end
        else
        begin
                myLocY_f <= myLocY;
                myLocX_f <= myLocX;
                myChipID_f <= myChipID;
        end
end
assign thanksIn_5 = thanks_0_to_5 | thanks_1_to_5 | thanks_2_to_5 | thanks_3_to_5 | thanks_4_to_5 | thanks_5_to_5 ;
assign validOut_5 = validOut_5_internal;
assign dataOut_5 = dataOut_5_internal;
assign yummyIn_5_internal = yummyIn_5;
assign yummyOut_5 = yummyOut_5_internal;
io_xbar_flip_bus #(1, 14) yummyOut_0_flip1(yummyOut_0_internal, yummyOut_0_flip1_out);
io_xbar_flip_bus #(1, 14) yummyOut_1_flip1(yummyOut_1_internal, yummyOut_1_flip1_out);
io_xbar_flip_bus #(1, 14) yummyOut_2_flip1(yummyOut_2_internal, yummyOut_2_flip1_out);
io_xbar_flip_bus #(1, 14) yummyOut_3_flip1(yummyOut_3_internal, yummyOut_3_flip1_out);
io_xbar_flip_bus #(1, 14) yummyOut_4_flip1(yummyOut_4_internal, yummyOut_4_flip1_out);
io_xbar_flip_bus #(1, 21) yummyOut_0_flip2(yummyOut_0_flip1_out, yummyOut_0);
io_xbar_flip_bus #(1, 21) yummyOut_1_flip2(yummyOut_1_flip1_out, yummyOut_1);
io_xbar_flip_bus #(1, 21) yummyOut_2_flip2(yummyOut_2_flip1_out, yummyOut_2);
io_xbar_flip_bus #(1, 21) yummyOut_3_flip2(yummyOut_3_flip1_out, yummyOut_3);
io_xbar_flip_bus #(1, 21) yummyOut_4_flip2(yummyOut_4_flip1_out, yummyOut_4);
io_xbar_flip_bus #(1, 14) validOut_0_flip1(validOut_0_internal, validOut_0_flip1_out);
io_xbar_flip_bus #(1, 14) validOut_1_flip1(validOut_1_internal, validOut_1_flip1_out);
io_xbar_flip_bus #(1, 14) validOut_2_flip1(validOut_2_internal, validOut_2_flip1_out);
io_xbar_flip_bus #(1, 14) validOut_3_flip1(validOut_3_internal, validOut_3_flip1_out);
io_xbar_flip_bus #(1, 14) validOut_4_flip1(validOut_4_internal, validOut_4_flip1_out);
io_xbar_flip_bus #(1, 21) validOut_0_flip2(validOut_0_flip1_out, validOut_0);
io_xbar_flip_bus #(1, 21) validOut_1_flip2(validOut_1_flip1_out, validOut_1);
io_xbar_flip_bus #(1, 21) validOut_2_flip2(validOut_2_flip1_out, validOut_2);
io_xbar_flip_bus #(1, 21) validOut_3_flip2(validOut_3_flip1_out, validOut_3);
io_xbar_flip_bus #(1, 21) validOut_4_flip2(validOut_4_flip1_out, validOut_4);
io_xbar_flip_bus #(64, 14) dataOut_0_flip1(dataOut_0_internal, dataOut_0_flip1_out);
io_xbar_flip_bus #(64, 14) dataOut_1_flip1(dataOut_1_internal, dataOut_1_flip1_out);
io_xbar_flip_bus #(64, 14) dataOut_2_flip1(dataOut_2_internal, dataOut_2_flip1_out);
io_xbar_flip_bus #(64, 14) dataOut_3_flip1(dataOut_3_internal, dataOut_3_flip1_out);
io_xbar_flip_bus #(64, 14) dataOut_4_flip1(dataOut_4_internal, dataOut_4_flip1_out);
io_xbar_flip_bus #(64, 21) dataOut_0_flip2(dataOut_0_flip1_out, dataOut_0);
io_xbar_flip_bus #(64, 21) dataOut_1_flip2(dataOut_1_flip1_out, dataOut_1);
io_xbar_flip_bus #(64, 21) dataOut_2_flip2(dataOut_2_flip1_out, dataOut_2);
io_xbar_flip_bus #(64, 21) dataOut_3_flip2(dataOut_3_flip1_out, dataOut_3);
io_xbar_flip_bus #(64, 21) dataOut_4_flip2(dataOut_4_flip1_out, dataOut_4);
io_xbar_flip_bus #(1, 14) yummyIn_0_flip1(yummyIn_0, yummyIn_0_flip1_out);
io_xbar_flip_bus #(1, 14) yummyIn_1_flip1(yummyIn_1, yummyIn_1_flip1_out);
io_xbar_flip_bus #(1, 14) yummyIn_2_flip1(yummyIn_2, yummyIn_2_flip1_out);
io_xbar_flip_bus #(1, 14) yummyIn_3_flip1(yummyIn_3, yummyIn_3_flip1_out);
io_xbar_flip_bus #(1, 14) yummyIn_4_flip1(yummyIn_4, yummyIn_4_flip1_out);
io_xbar_flip_bus #(1, 10) yummyIn_0_flip2(yummyIn_0_flip1_out, yummyIn_0_internal);
io_xbar_flip_bus #(1, 10) yummyIn_1_flip2(yummyIn_1_flip1_out, yummyIn_1_internal);
io_xbar_flip_bus #(1, 10) yummyIn_2_flip2(yummyIn_2_flip1_out, yummyIn_2_internal);
io_xbar_flip_bus #(1, 10) yummyIn_3_flip2(yummyIn_3_flip1_out, yummyIn_3_internal);
io_xbar_flip_bus #(1, 10) yummyIn_4_flip2(yummyIn_4_flip1_out, yummyIn_4_internal);
io_xbar_flip_bus #(1, 14) validIn_0_flip1(validIn_0, validIn_0_flip1_out);
io_xbar_flip_bus #(1, 14) validIn_1_flip1(validIn_1, validIn_1_flip1_out);
io_xbar_flip_bus #(1, 14) validIn_2_flip1(validIn_2, validIn_2_flip1_out);
io_xbar_flip_bus #(1, 14) validIn_3_flip1(validIn_3, validIn_3_flip1_out);
io_xbar_flip_bus #(1, 14) validIn_4_flip1(validIn_4, validIn_4_flip1_out);
io_xbar_flip_bus #(1, 10) validIn_0_flip2(validIn_0_flip1_out, validIn_0_internal);
io_xbar_flip_bus #(1, 10) validIn_1_flip2(validIn_1_flip1_out, validIn_1_internal);
io_xbar_flip_bus #(1, 10) validIn_2_flip2(validIn_2_flip1_out, validIn_2_internal);
io_xbar_flip_bus #(1, 10) validIn_3_flip2(validIn_3_flip1_out, validIn_3_internal);
io_xbar_flip_bus #(1, 10) validIn_4_flip2(validIn_4_flip1_out, validIn_4_internal);
io_xbar_flip_bus #(64, 14) dataIn_0_flip1(dataIn_0, dataIn_0_flip1_out);
io_xbar_flip_bus #(64, 14) dataIn_1_flip1(dataIn_1, dataIn_1_flip1_out);
io_xbar_flip_bus #(64, 14) dataIn_2_flip1(dataIn_2, dataIn_2_flip1_out);
io_xbar_flip_bus #(64, 14) dataIn_3_flip1(dataIn_3, dataIn_3_flip1_out);
io_xbar_flip_bus #(64, 14) dataIn_4_flip1(dataIn_4, dataIn_4_flip1_out);
io_xbar_flip_bus #(64, 10) dataIn_0_flip2(dataIn_0_flip1_out, dataIn_0_internal);
io_xbar_flip_bus #(64, 10) dataIn_1_flip2(dataIn_1_flip1_out, dataIn_1_internal);
io_xbar_flip_bus #(64, 10) dataIn_2_flip2(dataIn_2_flip1_out, dataIn_2_internal);
io_xbar_flip_bus #(64, 10) dataIn_3_flip2(dataIn_3_flip1_out, dataIn_3_internal);
io_xbar_flip_bus #(64, 10) dataIn_4_flip2(dataIn_4_flip1_out, dataIn_4_internal);
io_xbar_input_top_4 node_0_input(.route_req_0_out(route_req_0_to_0), .route_req_1_out(route_req_0_to_1), .route_req_2_out(route_req_0_to_2), .route_req_3_out(route_req_0_to_3), .route_req_4_out(route_req_0_to_4), .route_req_5_out(route_req_0_to_5), .default_ready_0_out(), .default_ready_1_out(), .default_ready_2_out(), .default_ready_3_out(default_ready_0_to_3), .default_ready_4_out(), .default_ready_5_out(), .tail_out(node_0_input_tail), .yummy_out(yummyOut_0_internal), .data_out(node_0_input_data), .valid_out(node_0_input_valid), .clk(clk), .reset(reset), .my_loc_x_in(myLocX_f), .my_loc_y_in(myLocY_f), .my_chip_id_in(myChipID_f), .valid_in(validIn_0_internal), .data_in(dataIn_0_internal), .thanks_0(thanks_0_to_0), .thanks_1(thanks_1_to_0), .thanks_2(thanks_2_to_0), .thanks_3(thanks_3_to_0), .thanks_4(thanks_4_to_0), .thanks_5(thanks_5_to_0));
io_xbar_input_top_4 node_1_input(.route_req_0_out(route_req_1_to_0), .route_req_1_out(route_req_1_to_1), .route_req_2_out(route_req_1_to_2), .route_req_3_out(route_req_1_to_3), .route_req_4_out(route_req_1_to_4), .route_req_5_out(route_req_1_to_5), .default_ready_0_out(), .default_ready_1_out(), .default_ready_2_out(), .default_ready_3_out(), .default_ready_4_out(default_ready_1_to_4), .default_ready_5_out(), .tail_out(node_1_input_tail), .yummy_out(yummyOut_1_internal), .data_out(node_1_input_data), .valid_out(node_1_input_valid), .clk(clk), .reset(reset), .my_loc_x_in(myLocX_f), .my_loc_y_in(myLocY_f), .my_chip_id_in(myChipID_f), .valid_in(validIn_1_internal), .data_in(dataIn_1_internal), .thanks_0(thanks_0_to_1), .thanks_1(thanks_1_to_1), .thanks_2(thanks_2_to_1), .thanks_3(thanks_3_to_1), .thanks_4(thanks_4_to_1), .thanks_5(thanks_5_to_1));
io_xbar_input_top_4 node_2_input(.route_req_0_out(route_req_2_to_0), .route_req_1_out(route_req_2_to_1), .route_req_2_out(route_req_2_to_2), .route_req_3_out(route_req_2_to_3), .route_req_4_out(route_req_2_to_4), .route_req_5_out(route_req_2_to_5), .default_ready_0_out(default_ready_2_to_0), .default_ready_1_out(), .default_ready_2_out(), .default_ready_3_out(), .default_ready_4_out(), .default_ready_5_out(default_ready_2_to_5), .tail_out(node_2_input_tail), .yummy_out(yummyOut_2_internal), .data_out(node_2_input_data), .valid_out(node_2_input_valid), .clk(clk), .reset(reset), .my_loc_x_in(myLocX_f), .my_loc_y_in(myLocY_f), .my_chip_id_in(myChipID_f), .valid_in(validIn_2_internal), .data_in(dataIn_2_internal), .thanks_0(thanks_0_to_2), .thanks_1(thanks_1_to_2), .thanks_2(thanks_2_to_2), .thanks_3(thanks_3_to_2), .thanks_4(thanks_4_to_2), .thanks_5(thanks_5_to_2));
io_xbar_input_top_4 node_3_input(.route_req_0_out(route_req_3_to_0), .route_req_1_out(route_req_3_to_1), .route_req_2_out(route_req_3_to_2), .route_req_3_out(route_req_3_to_3), .route_req_4_out(route_req_3_to_4), .route_req_5_out(route_req_3_to_5), .default_ready_0_out(), .default_ready_1_out(default_ready_3_to_1), .default_ready_2_out(), .default_ready_3_out(), .default_ready_4_out(), .default_ready_5_out(), .tail_out(node_3_input_tail), .yummy_out(yummyOut_3_internal), .data_out(node_3_input_data), .valid_out(node_3_input_valid), .clk(clk), .reset(reset), .my_loc_x_in(myLocX_f), .my_loc_y_in(myLocY_f), .my_chip_id_in(myChipID_f), .valid_in(validIn_3_internal), .data_in(dataIn_3_internal), .thanks_0(thanks_0_to_3), .thanks_1(thanks_1_to_3), .thanks_2(thanks_2_to_3), .thanks_3(thanks_3_to_3), .thanks_4(thanks_4_to_3), .thanks_5(thanks_5_to_3));
io_xbar_input_top_4 node_4_input(.route_req_0_out(route_req_4_to_0), .route_req_1_out(route_req_4_to_1), .route_req_2_out(route_req_4_to_2), .route_req_3_out(route_req_4_to_3), .route_req_4_out(route_req_4_to_4), .route_req_5_out(route_req_4_to_5), .default_ready_0_out(), .default_ready_1_out(), .default_ready_2_out(default_ready_4_to_2), .default_ready_3_out(), .default_ready_4_out(), .default_ready_5_out(), .tail_out(node_4_input_tail), .yummy_out(yummyOut_4_internal), .data_out(node_4_input_data), .valid_out(node_4_input_valid), .clk(clk), .reset(reset), .my_loc_x_in(myLocX_f), .my_loc_y_in(myLocY_f), .my_chip_id_in(myChipID_f), .valid_in(validIn_4_internal), .data_in(dataIn_4_internal), .thanks_0(thanks_0_to_4), .thanks_1(thanks_1_to_4), .thanks_2(thanks_2_to_4), .thanks_3(thanks_3_to_4), .thanks_4(thanks_4_to_4), .thanks_5(thanks_5_to_4));
io_xbar_input_top_4 node_5_input(.route_req_0_out(route_req_5_to_0), .route_req_1_out(route_req_5_to_1), .route_req_2_out(route_req_5_to_2), .route_req_3_out(route_req_5_to_3), .route_req_4_out(route_req_5_to_4), .route_req_5_out(route_req_5_to_5), .default_ready_0_out(), .default_ready_1_out(), .default_ready_2_out(), .default_ready_3_out(), .default_ready_4_out(), .default_ready_5_out(), .tail_out(node_5_input_tail), .yummy_out(yummyOut_5_internal), .data_out(node_5_input_data), .valid_out(node_5_input_valid), .clk(clk), .reset(reset), .my_loc_x_in(myLocX_f), .my_loc_y_in(myLocY_f), .my_chip_id_in(myChipID_f), .valid_in(validIn_5), .data_in(dataIn_5), .thanks_0(thanks_0_to_5), .thanks_1(thanks_1_to_5), .thanks_2(thanks_2_to_5), .thanks_3(thanks_3_to_5), .thanks_4(thanks_4_to_5), .thanks_5(thanks_5_to_5));
io_xbar_output_top node_0_output(.data_out(dataOut_0_internal), .thanks_0_out(thanks_0_to_2), .thanks_1_out(thanks_0_to_3), .thanks_2_out(thanks_0_to_4), .thanks_3_out(thanks_0_to_5), .thanks_4_out(thanks_0_to_1), .thanks_5_out(thanks_0_to_0), .valid_out(validOut_0_internal), .popped_interrupt_mesg_out(), .popped_memory_ack_mesg_out(), .popped_memory_ack_mesg_out_sender(), .ec_wants_to_send_but_cannot(ec_wants_to_send_but_cannot_0), .clk(clk), .reset(reset), .route_req_0_in(route_req_2_to_0), .route_req_1_in(route_req_3_to_0), .route_req_2_in(route_req_4_to_0), .route_req_3_in(route_req_5_to_0), .route_req_4_in(route_req_1_to_0), .route_req_5_in(route_req_0_to_0), .tail_0_in(node_2_input_tail), .tail_1_in(node_3_input_tail), .tail_2_in(node_4_input_tail), .tail_3_in(node_5_input_tail), .tail_4_in(node_1_input_tail), .tail_5_in(node_0_input_tail), .data_0_in(node_2_input_data), .data_1_in(node_3_input_data), .data_2_in(node_4_input_data), .data_3_in(node_5_input_data), .data_4_in(node_1_input_data), .data_5_in(node_0_input_data), .valid_0_in(node_2_input_valid), .valid_1_in(node_3_input_valid), .valid_2_in(node_4_input_valid), .valid_3_in(node_5_input_valid), .valid_4_in(node_1_input_valid), .valid_5_in(node_0_input_valid), .default_ready_in(default_ready_2_to_0),.yummy_in(yummyIn_0_internal));
io_xbar_output_top node_1_output(.data_out(dataOut_1_internal), .thanks_0_out(thanks_1_to_3), .thanks_1_out(thanks_1_to_4), .thanks_2_out(thanks_1_to_5), .thanks_3_out(thanks_1_to_0), .thanks_4_out(thanks_1_to_2), .thanks_5_out(thanks_1_to_1), .valid_out(validOut_1_internal), .popped_interrupt_mesg_out(), .popped_memory_ack_mesg_out(), .popped_memory_ack_mesg_out_sender(), .ec_wants_to_send_but_cannot(ec_wants_to_send_but_cannot_1), .clk(clk), .reset(reset), .route_req_0_in(route_req_3_to_1), .route_req_1_in(route_req_4_to_1), .route_req_2_in(route_req_5_to_1), .route_req_3_in(route_req_0_to_1), .route_req_4_in(route_req_2_to_1), .route_req_5_in(route_req_1_to_1), .tail_0_in(node_3_input_tail), .tail_1_in(node_4_input_tail), .tail_2_in(node_5_input_tail), .tail_3_in(node_0_input_tail), .tail_4_in(node_2_input_tail), .tail_5_in(node_1_input_tail), .data_0_in(node_3_input_data), .data_1_in(node_4_input_data), .data_2_in(node_5_input_data), .data_3_in(node_0_input_data), .data_4_in(node_2_input_data), .data_5_in(node_1_input_data), .valid_0_in(node_3_input_valid), .valid_1_in(node_4_input_valid), .valid_2_in(node_5_input_valid), .valid_3_in(node_0_input_valid), .valid_4_in(node_2_input_valid), .valid_5_in(node_1_input_valid), .default_ready_in(default_ready_3_to_1),.yummy_in(yummyIn_1_internal));
io_xbar_output_top node_2_output(.data_out(dataOut_2_internal), .thanks_0_out(thanks_2_to_4), .thanks_1_out(thanks_2_to_5), .thanks_2_out(thanks_2_to_0), .thanks_3_out(thanks_2_to_1), .thanks_4_out(thanks_2_to_3), .thanks_5_out(thanks_2_to_2), .valid_out(validOut_2_internal), .popped_interrupt_mesg_out(), .popped_memory_ack_mesg_out(), .popped_memory_ack_mesg_out_sender(), .ec_wants_to_send_but_cannot(ec_wants_to_send_but_cannot_2), .clk(clk), .reset(reset), .route_req_0_in(route_req_4_to_2), .route_req_1_in(route_req_5_to_2), .route_req_2_in(route_req_0_to_2), .route_req_3_in(route_req_1_to_2), .route_req_4_in(route_req_3_to_2), .route_req_5_in(route_req_2_to_2), .tail_0_in(node_4_input_tail), .tail_1_in(node_5_input_tail), .tail_2_in(node_0_input_tail), .tail_3_in(node_1_input_tail), .tail_4_in(node_3_input_tail), .tail_5_in(node_2_input_tail), .data_0_in(node_4_input_data), .data_1_in(node_5_input_data), .data_2_in(node_0_input_data), .data_3_in(node_1_input_data), .data_4_in(node_3_input_data), .data_5_in(node_2_input_data), .valid_0_in(node_4_input_valid), .valid_1_in(node_5_input_valid), .valid_2_in(node_0_input_valid), .valid_3_in(node_1_input_valid), .valid_4_in(node_3_input_valid), .valid_5_in(node_2_input_valid), .default_ready_in(default_ready_4_to_2),.yummy_in(yummyIn_2_internal));
io_xbar_output_top node_3_output(.data_out(dataOut_3_internal), .thanks_0_out(thanks_3_to_0), .thanks_1_out(thanks_3_to_1), .thanks_2_out(thanks_3_to_2), .thanks_3_out(thanks_3_to_4), .thanks_4_out(thanks_3_to_5), .thanks_5_out(thanks_3_to_3), .valid_out(validOut_3_internal), .popped_interrupt_mesg_out(), .popped_memory_ack_mesg_out(), .popped_memory_ack_mesg_out_sender(), .ec_wants_to_send_but_cannot(ec_wants_to_send_but_cannot_3), .clk(clk), .reset(reset), .route_req_0_in(route_req_0_to_3), .route_req_1_in(route_req_1_to_3), .route_req_2_in(route_req_2_to_3), .route_req_3_in(route_req_4_to_3), .route_req_4_in(route_req_5_to_3), .route_req_5_in(route_req_3_to_3), .tail_0_in(node_0_input_tail), .tail_1_in(node_1_input_tail), .tail_2_in(node_2_input_tail), .tail_3_in(node_4_input_tail), .tail_4_in(node_5_input_tail), .tail_5_in(node_3_input_tail), .data_0_in(node_0_input_data), .data_1_in(node_1_input_data), .data_2_in(node_2_input_data), .data_3_in(node_4_input_data), .data_4_in(node_5_input_data), .data_5_in(node_3_input_data), .valid_0_in(node_0_input_valid), .valid_1_in(node_1_input_valid), .valid_2_in(node_2_input_valid), .valid_3_in(node_4_input_valid), .valid_4_in(node_5_input_valid), .valid_5_in(node_3_input_valid), .default_ready_in(default_ready_0_to_3),.yummy_in(yummyIn_3_internal));
io_xbar_output_top node_4_output(.data_out(dataOut_4_internal), .thanks_0_out(thanks_4_to_1), .thanks_1_out(thanks_4_to_2), .thanks_2_out(thanks_4_to_3), .thanks_3_out(thanks_4_to_5), .thanks_4_out(thanks_4_to_0), .thanks_5_out(thanks_4_to_4), .valid_out(validOut_4_internal), .popped_interrupt_mesg_out(), .popped_memory_ack_mesg_out(), .popped_memory_ack_mesg_out_sender(), .ec_wants_to_send_but_cannot(ec_wants_to_send_but_cannot_4), .clk(clk), .reset(reset), .route_req_0_in(route_req_1_to_4), .route_req_1_in(route_req_2_to_4), .route_req_2_in(route_req_3_to_4), .route_req_3_in(route_req_5_to_4), .route_req_4_in(route_req_0_to_4), .route_req_5_in(route_req_4_to_4), .tail_0_in(node_1_input_tail), .tail_1_in(node_2_input_tail), .tail_2_in(node_3_input_tail), .tail_3_in(node_5_input_tail), .tail_4_in(node_0_input_tail), .tail_5_in(node_4_input_tail), .data_0_in(node_1_input_data), .data_1_in(node_2_input_data), .data_2_in(node_3_input_data), .data_3_in(node_5_input_data), .data_4_in(node_0_input_data), .data_5_in(node_4_input_data), .valid_0_in(node_1_input_valid), .valid_1_in(node_2_input_valid), .valid_2_in(node_3_input_valid), .valid_3_in(node_5_input_valid), .valid_4_in(node_0_input_valid), .valid_5_in(node_4_input_valid), .default_ready_in(default_ready_1_to_4),.yummy_in(yummyIn_4_internal));
io_xbar_output_top #(1'b0) node_5_output(.data_out(dataOut_5_internal), .thanks_0_out(thanks_5_to_2), .thanks_1_out(thanks_5_to_3), .thanks_2_out(thanks_5_to_4), .thanks_3_out(thanks_5_to_0), .thanks_4_out(thanks_5_to_1), .thanks_5_out(thanks_5_to_5), .valid_out(validOut_5_internal), .popped_interrupt_mesg_out(external_interrupt), .popped_memory_ack_mesg_out(store_ack_received), .popped_memory_ack_mesg_out_sender(store_ack_addr), .ec_wants_to_send_but_cannot(ec_wants_to_send_but_cannot_5), .clk(clk), .reset(reset), .route_req_0_in(route_req_2_to_5), .route_req_1_in(route_req_3_to_5), .route_req_2_in(route_req_4_to_5), .route_req_3_in(route_req_0_to_5), .route_req_4_in(route_req_1_to_5), .route_req_5_in(route_req_5_to_5), .tail_0_in(node_2_input_tail), .tail_1_in(node_3_input_tail), .tail_2_in(node_4_input_tail), .tail_3_in(node_0_input_tail), .tail_4_in(node_1_input_tail), .tail_5_in(node_5_input_tail), .data_0_in(node_2_input_data), .data_1_in(node_3_input_data), .data_2_in(node_4_input_data), .data_3_in(node_0_input_data), .data_4_in(node_1_input_data), .data_5_in(node_5_input_data), .valid_0_in(node_2_input_valid), .valid_1_in(node_3_input_valid), .valid_2_in(node_4_input_valid), .valid_3_in(node_0_input_valid), .valid_4_in(node_1_input_valid), .valid_5_in(node_5_input_valid), .default_ready_in(default_ready_2_to_5),.yummy_in(yummyIn_5_internal));
endmodule 
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
module sram_l15_data
(
input wire MEMCLK,
input wire RESET_N,
input wire CE,
input wire [9-1:0] A,
input wire RDWEN,
input wire [128-1:0] BW,
input wire [128-1:0] DIN,
output wire [128-1:0] DOUT,
input wire [4-1:0] BIST_COMMAND,
input wire [4-1:0] BIST_DIN,
output reg [4-1:0] BIST_DOUT,
input wire [8-1:0] SRAMID
);
wire [128-1:0] DOUT_bram;
assign DOUT = DOUT_bram;
bram_1rw_wrapper #(
   .NAME          (""             ),
   .DEPTH         (512),
   .ADDR_WIDTH    (9),
   .BITMASK_WIDTH (128),
   .DATA_WIDTH    (128)
)   sram_l15_data (
   .MEMCLK        (MEMCLK     ),
   .RESET_N        (RESET_N     ),
   .CE            (CE         ),
   .A             (A          ),
   .RDWEN         (RDWEN      ),
   .BW            (BW         ),
   .DIN           (DIN        ),
   .DOUT          (DOUT_bram       )
);
      
 
 endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
module sram_l15_hmt
(
input wire MEMCLK,
input wire RESET_N,
input wire CE,
input wire [9-1:0] A,
input wire RDWEN,
input wire [32-1:0] BW,
input wire [32-1:0] DIN,
output wire [32-1:0] DOUT,
input wire [4-1:0] BIST_COMMAND,
input wire [4-1:0] BIST_DIN,
output reg [4-1:0] BIST_DOUT,
input wire [8-1:0] SRAMID
);
wire [32-1:0] DOUT_bram;
assign DOUT = DOUT_bram;
bram_1rw_wrapper #(
   .NAME          (""             ),
   .DEPTH         (512),
   .ADDR_WIDTH    (9),
   .BITMASK_WIDTH (32),
   .DATA_WIDTH    (32)
)   sram_l15_hmt (
   .MEMCLK        (MEMCLK     ),
   .RESET_N        (RESET_N     ),
   .CE            (CE         ),
   .A             (A          ),
   .RDWEN         (RDWEN      ),
   .BW            (BW         ),
   .DIN           (DIN        ),
   .DOUT          (DOUT_bram       )
);
      
 
 endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
module sram_l15_tag
(
input wire MEMCLK,
input wire RESET_N,
input wire CE,
input wire [((9-2))-1:0] A,
input wire RDWEN,
input wire [33*4-1:0] BW,
input wire [33*4-1:0] DIN,
output wire [33*4-1:0] DOUT,
input wire [4-1:0] BIST_COMMAND,
input wire [4-1:0] BIST_DIN,
output reg [4-1:0] BIST_DOUT,
input wire [8-1:0] SRAMID
);
wire [33*4-1:0] DOUT_bram;
assign DOUT = DOUT_bram;
bram_1rw_wrapper #(
   .NAME          (""             ),
   .DEPTH         ((512/4)),
   .ADDR_WIDTH    (((9-2))),
   .BITMASK_WIDTH (33*4),
   .DATA_WIDTH    (33*4)
)   sram_l15_tag (
   .MEMCLK        (MEMCLK     ),
   .RESET_N        (RESET_N     ),
   .CE            (CE         ),
   .A             (A          ),
   .RDWEN         (RDWEN      ),
   .BW            (BW         ),
   .DIN           (DIN        ),
   .DOUT          (DOUT_bram       )
);
      
 
 endmodule
      
 
module sram_l2_data
(
input wire MEMCLK,
input wire RESET_N,
input wire CE,
input wire [12-1:0] A,
input wire RDWEN,
input wire [144-1:0] BW,
input wire [144-1:0] DIN,
output wire [144-1:0] DOUT,
input wire [4-1:0] BIST_COMMAND,
input wire [4-1:0] BIST_DIN,
output reg [4-1:0] BIST_DOUT,
input wire [8-1:0] SRAMID
);
wire [144-1:0] DOUT_bram;
assign DOUT = DOUT_bram;
bram_1rw_wrapper #(
   .NAME          (""             ),
   .DEPTH         (4096),
   .ADDR_WIDTH    (12),
   .BITMASK_WIDTH (144),
   .DATA_WIDTH    (144)
)   sram_l2_data (
   .MEMCLK        (MEMCLK     ),
   .RESET_N        (RESET_N     ),
   .CE            (CE         ),
   .A             (A          ),
   .RDWEN         (RDWEN      ),
   .BW            (BW         ),
   .DIN           (DIN        ),
   .DOUT          (DOUT_bram       )
);
      
 
 endmodule
      
 
module sram_l2_dir
(
input wire MEMCLK,
input wire RESET_N,
input wire CE,
input wire [10-1:0] A,
input wire RDWEN,
input wire [64-1:0] BW,
input wire [64-1:0] DIN,
output wire [64-1:0] DOUT,
input wire [4-1:0] BIST_COMMAND,
input wire [4-1:0] BIST_DIN,
output reg [4-1:0] BIST_DOUT,
input wire [8-1:0] SRAMID
);
wire [64-1:0] DOUT_bram;
assign DOUT = DOUT_bram;
bram_1rw_wrapper #(
   .NAME          (""             ),
   .DEPTH         (1024),
   .ADDR_WIDTH    (10),
   .BITMASK_WIDTH (64),
   .DATA_WIDTH    (64)
)   sram_l2_dir (
   .MEMCLK        (MEMCLK     ),
   .RESET_N        (RESET_N     ),
   .CE            (CE         ),
   .A             (A          ),
   .RDWEN         (RDWEN      ),
   .BW            (BW         ),
   .DIN           (DIN        ),
   .DOUT          (DOUT_bram       )
);
      
 
 endmodule
      
 
module sram_l2_state
(
input wire MEMCLK,
input wire RESET_N,
input wire CEA,
input wire [8-1:0] AA,
input wire RDWENA,
input wire CEB,
input wire [8-1:0] AB,
input wire RDWENB,
input wire [15*4+2+4-1:0] BWA,
input wire [15*4+2+4-1:0] DINA,
output wire [15*4+2+4-1:0] DOUTA,
input wire [15*4+2+4-1:0] BWB,
input wire [15*4+2+4-1:0] DINB,
output wire [15*4+2+4-1:0] DOUTB,
input wire [4-1:0] BIST_COMMAND,
input wire [4-1:0] BIST_DIN,
output reg [4-1:0] BIST_DOUT,
input wire [8-1:0] SRAMID
);
  
wire [15*4+2+4-1:0] DOUTA_bram;
wire [15*4+2+4-1:0] DOUTB_bram;
assign DOUTA = DOUTA_bram;
assign DOUTB = DOUTB_bram;
bram_1r1w_wrapper #(
   .NAME          (""             ),
   .DEPTH         (256),
   .ADDR_WIDTH    (8),
   .BITMASK_WIDTH (15*4+2+4),
   .DATA_WIDTH    (15*4+2+4)
)   sram_l2_state (
   .MEMCLK        (MEMCLK     ),
   .RESET_N        (RESET_N     ),
   .CEA        (CEA     ),
   .AA        (AA     ),
   .AB        (AB     ),
   .RDWENA        (RDWENA     ),
   .CEB        (CEB     ),
   .RDWENB        (RDWENB     ),
   .BWA        (BWA     ),
   .DINA        (DINA     ),
   .DOUTA        (DOUTA_bram     ),
   .BWB        (BWB     ),
   .DINB        (DINB     ),
   .DOUTB        (DOUTB_bram     )
);
      
  
 
 endmodule
      
 
module sram_l2_tag
(
input wire MEMCLK,
input wire RESET_N,
input wire CE,
input wire [8-1:0] A,
input wire RDWEN,
input wire [104-1:0] BW,
input wire [104-1:0] DIN,
output wire [104-1:0] DOUT,
input wire [4-1:0] BIST_COMMAND,
input wire [4-1:0] BIST_DIN,
output reg [4-1:0] BIST_DOUT,
input wire [8-1:0] SRAMID
);
wire [104-1:0] DOUT_bram;
assign DOUT = DOUT_bram;
bram_1rw_wrapper #(
   .NAME          (""             ),
   .DEPTH         (256),
   .ADDR_WIDTH    (8),
   .BITMASK_WIDTH (104),
   .DATA_WIDTH    (104)
)   sram_l2_tag (
   .MEMCLK        (MEMCLK     ),
   .RESET_N        (RESET_N     ),
   .CE            (CE         ),
   .A             (A          ),
   .RDWEN         (RDWEN      ),
   .BW            (BW         ),
   .DIN           (DIN        ),
   .DOUT          (DOUT_bram       )
);
      
 
 endmodule
module noc_axilite_bridge #(
    
    
    
    parameter SLAVE_RESP_BYTEWIDTH = 4,
    
    parameter SWAP_ENDIANESS       = 0,
    
    parameter ALIGN_RDATA          = 1
) (
    
    input  wire                                   clk,
    input  wire                                   rst,
    
    input  wire                                   splitter_bridge_val,
    input  wire [64-1:0]             splitter_bridge_data,
    output wire                                   bridge_splitter_rdy,
    
    output  reg                                   bridge_splitter_val,
    output  reg  [64-1:0]            bridge_splitter_data,
    input  wire                                   splitter_bridge_rdy,
    
    output  reg  [64-1:0]   m_axi_awaddr,
    output  reg                                   m_axi_awvalid,
    input  wire                                   m_axi_awready,
    
    output wire  [64-1:0]   m_axi_wdata,
    output  reg  [64/8-1:0] m_axi_wstrb,
    output  reg                                   m_axi_wvalid,
    input  wire                                   m_axi_wready,
    
    output  reg  [64-1:0]   m_axi_araddr,
    output  reg                                   m_axi_arvalid,
    input                                         m_axi_arready,
    
    input  wire [64-1:0]    m_axi_rdata,
    input  wire [2-1:0]    m_axi_rresp,
    input  wire                                   m_axi_rvalid,
    output  reg                                   m_axi_rready,
    
    input  wire [2-1:0]    m_axi_bresp,
    input  wire                                   m_axi_bvalid,
    output reg                                    m_axi_bready,
    
    output  reg  [3-1:0]   w_reqbuf_size,
    output  reg  [3-1:0]   r_reqbuf_size
);
localparam MSG_STATE_INVAL      = 3'd0; 
localparam MSG_STATE_HEADER_0   = 3'd1; 
localparam MSG_STATE_HEADER_1   = 3'd2; 
localparam MSG_STATE_HEADER_2   = 3'd3; 
localparam MSG_STATE_DATA       = 3'd4; 
localparam MSG_TYPE_INVAL       = 2'd0; 
localparam MSG_TYPE_LOAD        = 2'd1; 
localparam MSG_TYPE_STORE       = 2'd2; 
localparam BUF_STATUS_INCOMP    = 2'd0; 
localparam BUF_STATUS_COMP      = 2'd1; 
localparam BUF_STATUS_WAITRESP  = 2'd2; 
localparam BUF_STATUS_RESPSEND  = 2'd3; 
localparam LOAD_ACK = 1'd0;
localparam STORE_ACK = 1'd1;
 reg  [2:0]                          splitter_io_msg_state_f;
 reg  [1:0]                          splitter_io_msg_type_f;
 reg  [8-1:0]        splitter_io_msg_counter_f;
 reg  [64-1:0]          r_req_buf_header0_f;
 reg  [64-1:0]          r_req_buf_header1_f;
 reg  [64-1:0]          r_req_buf_header2_f;
 reg  [1:0]                          r_req_buf_status_f;
 reg  [64-1:0]          w_req_buf_header0_f;
 reg  [64-1:0]          w_req_buf_header1_f;
 reg  [64-1:0]          w_req_buf_header2_f;
 reg  [64-1:0]          w_req_buf_data0_f;
 wire [1:0]                          w_req_buf_status;
 reg  [1:0]                          w_addr_req_buf_status_f;
 reg  [1:0]                          w_data_req_buf_status_f;
 reg  [64-1:0]          r_resp_buf_header0_f;
 reg  [64-1:0] r_resp_buf_data0_f;
 reg  [2-1:0] r_resp_buf_rresp_f;
 reg  [1:0]                          r_resp_buf_status_f;
 reg  [64-1:0]          w_resp_buf_header0_f;
 reg  [2-1:0] w_resp_buf_bresp_f;
 wire [1:0]                          w_resp_buf_status;
 reg  [1:0]                          w_addr_resp_buf_status_f;
 reg  [1:0]                          w_data_resp_buf_status_f;
 wire                         splitter_io_go;
 wire                         splitter_io_load_go;
 wire                         splitter_io_store_go;
 wire                         splitter_io_msg_is_load;
 wire                         splitter_io_msg_is_store;
 wire                         splitter_io_msg_is_load_next;
 wire                         splitter_io_msg_is_store_next;
 wire [2:0]                   splitter_io_msg_state_next;
 wire [2:0]                   splitter_io_msg_type_mux_out;
 wire [2:0]                   splitter_io_msg_type_next;
 wire [8-1:0] splitter_io_msg_counter_next;
 wire                         m_axi_ar_go;
 wire                         m_axi_w_go;
 wire                         m_axi_aw_go;
 wire                         m_axi_b_go;
 wire                         m_axi_r_go;
 reg  [64-1:0]   a_axi_rdata_shifted;
 wire [64-1:0]   a_axi_rdata_masked;
 wire [64-1:0]   r_resp_buf_header0_next;
 wire [64-1:0]   w_resp_buf_header0_next;
 reg  [8-1:0] io_splitter_ack_load_counter_f;
 reg                          io_splitter_arb_f;
 reg                          io_splitter_ack_mux_sel;
 wire                         r_resp_buf_val;
 wire                         w_resp_buf_val;
 wire [64-1:0]   io_splitter_ack_store;
 wire [64-1:0]   io_splitter_ack_load;
 wire                         io_splitter_ack_load_go;
 wire                         io_splitter_ack_store_go;
    
    assign splitter_io_msg_type_mux_out =
        (!splitter_bridge_val) ? MSG_TYPE_INVAL :
        (((splitter_bridge_data[21:14] == 8'd31   )  ||
          (splitter_bridge_data[21:14] == 8'd14)  ||
          (splitter_bridge_data[21:14] == 8'd19   )     ) ? MSG_TYPE_LOAD  :
         ((splitter_bridge_data[21:14] == 8'd2   ) ||
          (splitter_bridge_data[21:14] == 8'd15) ||
          (splitter_bridge_data[21:14] == 8'd20   )    ) ? MSG_TYPE_STORE :
                                                                            MSG_TYPE_INVAL );
    
    assign splitter_io_msg_type_next =
        (splitter_io_msg_state_next == MSG_STATE_INVAL   ) ? MSG_TYPE_INVAL               :
        (splitter_io_msg_state_next == MSG_STATE_HEADER_0) ? splitter_io_msg_type_mux_out :
                                                             splitter_io_msg_type_f       ;
    
    assign splitter_io_msg_is_load       = (splitter_io_msg_type_f    == MSG_TYPE_LOAD );
    assign splitter_io_msg_is_store      = (splitter_io_msg_type_f    == MSG_TYPE_STORE);
    
    assign splitter_io_msg_is_load_next  = (splitter_io_msg_type_next == MSG_TYPE_LOAD );
    assign splitter_io_msg_is_store_next = (splitter_io_msg_type_next == MSG_TYPE_STORE);
    
    assign splitter_io_go = splitter_bridge_val && bridge_splitter_rdy;
    
    assign splitter_io_load_go  = splitter_io_msg_is_load_next  && splitter_io_go && (r_req_buf_status_f == BUF_STATUS_INCOMP);
    assign splitter_io_store_go = splitter_io_msg_is_store_next && splitter_io_go && (w_req_buf_status   == BUF_STATUS_INCOMP);
    
    assign splitter_io_msg_state_next =
        (splitter_io_msg_state_f == MSG_STATE_INVAL   ) ? MSG_STATE_HEADER_0  :
        (splitter_io_msg_state_f == MSG_STATE_HEADER_0) ? MSG_STATE_HEADER_1  :
        (splitter_io_msg_state_f == MSG_STATE_HEADER_1) ? MSG_STATE_HEADER_2  :
        (splitter_io_msg_counter_f == 0               ) ? MSG_STATE_HEADER_0  :
        (splitter_io_msg_state_f == MSG_STATE_HEADER_2) ? MSG_STATE_DATA      :
        (splitter_io_msg_state_f == MSG_STATE_DATA    ) ? MSG_STATE_DATA      :
                                                          MSG_STATE_INVAL     ;
    
    assign splitter_io_msg_counter_next =
        (splitter_io_msg_state_next == MSG_STATE_HEADER_0) ? splitter_bridge_data[29:22] :
                                                             splitter_io_msg_counter_f - 1'b1  ;
    
    
    
    always @(posedge clk) begin
        if (rst) begin
            splitter_io_msg_state_f   <= MSG_STATE_INVAL;
            splitter_io_msg_type_f    <= MSG_TYPE_INVAL;
            splitter_io_msg_counter_f <= {8{1'b0}};
        end
        else begin
            splitter_io_msg_state_f   <= splitter_io_go ? splitter_io_msg_state_next
                                                        : splitter_io_msg_state_f;
            splitter_io_msg_type_f    <= splitter_io_go ? splitter_io_msg_type_next
                                                        : splitter_io_msg_type_f;
            splitter_io_msg_counter_f <= splitter_io_go ? splitter_io_msg_counter_next
                                                        : splitter_io_msg_counter_f;
        end
    end
    
    
    
    always @(posedge clk) begin
        if (rst) begin
            r_req_buf_header0_f <= {64{1'b0}};
            r_req_buf_header1_f <= {64{1'b0}};
            r_req_buf_header2_f <= {64{1'b0}};
            r_req_buf_status_f  <= BUF_STATUS_INCOMP;
        end
        else begin
            r_req_buf_header0_f <= (splitter_io_load_go &
                                    (splitter_io_msg_state_next == MSG_STATE_HEADER_0)) ? splitter_bridge_data :
                                                                                          r_req_buf_header0_f  ;
            r_req_buf_header1_f <= (splitter_io_load_go &
                                    (splitter_io_msg_state_next == MSG_STATE_HEADER_1)) ? splitter_bridge_data :
                                                                                          r_req_buf_header1_f  ;
            r_req_buf_header2_f <= (splitter_io_load_go &
                                    (splitter_io_msg_state_next == MSG_STATE_HEADER_2)) ? splitter_bridge_data :
                                                                                          r_req_buf_header2_f  ;
            r_req_buf_status_f  <= (splitter_io_load_go &
                                    (splitter_io_msg_state_next == MSG_STATE_HEADER_2)) ? BUF_STATUS_COMP      :
                                   (m_axi_ar_go)                                        ? BUF_STATUS_INCOMP    :
                                                                                          r_req_buf_status_f   ;
        end
    end
    
    
    
    wire    w_status_update;
    assign  w_status_update =   splitter_io_store_go &
                                (splitter_io_msg_state_next == MSG_STATE_DATA) &
                                (splitter_io_msg_counter_f == 8'd1);
    always @(posedge clk) begin
        if (rst) begin
            w_req_buf_header0_f     <= {64{1'b0}};
            w_req_buf_header1_f     <= {64{1'b0}};
            w_req_buf_header2_f     <= {64{1'b0}};
            w_req_buf_data0_f       <= {64{1'b0}};
            w_addr_req_buf_status_f <= BUF_STATUS_INCOMP;
            w_data_req_buf_status_f <= BUF_STATUS_INCOMP;
        end
        else begin
            w_req_buf_header0_f     <= (splitter_io_store_go &
                                        (splitter_io_msg_state_next == MSG_STATE_HEADER_0)) ? splitter_bridge_data    :
                                                                                              w_req_buf_header0_f     ;
            w_req_buf_header1_f     <= (splitter_io_store_go &
                                        (splitter_io_msg_state_next == MSG_STATE_HEADER_1)) ? splitter_bridge_data    :
                                                                                              w_req_buf_header1_f     ;
            w_req_buf_header2_f     <= (splitter_io_store_go &
                                        (splitter_io_msg_state_next == MSG_STATE_HEADER_2)) ? splitter_bridge_data    :
                                                                                              w_req_buf_header2_f     ;
            w_req_buf_data0_f       <= (splitter_io_store_go &
                                        (splitter_io_msg_state_next == MSG_STATE_DATA))     ? splitter_bridge_data    :
                                                                                              w_req_buf_data0_f       ;
            w_addr_req_buf_status_f <= w_status_update                                      ? BUF_STATUS_COMP         :
                                       m_axi_aw_go                                          ? BUF_STATUS_INCOMP       :
                                                                                              w_addr_req_buf_status_f ;
            w_data_req_buf_status_f <= w_status_update                                      ? BUF_STATUS_COMP         :
                                       m_axi_w_go                                           ? BUF_STATUS_INCOMP       :
                                                                                              w_data_req_buf_status_f ;
        end
    end
    
    assign w_req_buf_status =
        ((w_addr_req_buf_status_f == BUF_STATUS_INCOMP) &&
         (w_data_req_buf_status_f == BUF_STATUS_INCOMP)    ) ? BUF_STATUS_INCOMP :
                                                               BUF_STATUS_COMP   ;
    wire [64-1:0]          paddings;
    reg  [64-1:0] m_axi_wdata_tmp;
    assign paddings = 0;
    
    always @ (*) begin
        
        m_axi_awvalid = (w_req_buf_status == BUF_STATUS_COMP) && (w_addr_resp_buf_status_f == BUF_STATUS_INCOMP);
        m_axi_awaddr = {paddings[64-1:40], w_req_buf_header1_f[(16 + 40 - 1):(16 + 40 - 1)-39]};
        
        m_axi_wvalid    = (w_req_buf_status == BUF_STATUS_COMP) && (w_data_resp_buf_status_f == BUF_STATUS_INCOMP);
        m_axi_wdata_tmp = w_req_buf_data0_f[64-1:0];
        
        m_axi_arvalid = (r_req_buf_status_f == BUF_STATUS_COMP) && (r_resp_buf_status_f == BUF_STATUS_INCOMP);
        m_axi_araddr = {paddings[64-1:40], r_req_buf_header1_f[(16 + 40 - 1):(16 + 40 - 1)-39]};
    end
    
    always @ (*) begin
        if (w_req_buf_header1_f[10:8] == 3'b000) begin
            m_axi_wstrb   = 8'b00000000;
            w_reqbuf_size = 3'b00;
        end
        else if (w_req_buf_header1_f[10:8] == 3'b001) begin
            m_axi_wstrb   = 8'b00000001;
            w_reqbuf_size = 3'b00;
        end
        else if (w_req_buf_header1_f[10:8] == 3'b010) begin
            m_axi_wstrb   = 8'b00000011;
            w_reqbuf_size = 3'b01;
        end
        else if (w_req_buf_header1_f[10:8] == 3'b011) begin
            m_axi_wstrb   = 8'b00001111;
            w_reqbuf_size = 3'b10;
        end
        else if (w_req_buf_header1_f[10:8] == 3'b100) begin
            m_axi_wstrb   = 8'b11111111;
            w_reqbuf_size = 3'b11;
        end
        else begin
            m_axi_wstrb   = 8'b11111111;
            w_reqbuf_size = 3'b11;
        end
    end
    generate
        if (SWAP_ENDIANESS) begin
            initial begin : p_endianess_check
              if (!(64 == 64 && 64 == 64))
                  $fatal(1,"swapped endianess only works for 64bit NOC and AXI bus");
            end
            
            
            assign m_axi_wdata[56 +: 8] = m_axi_wdata_tmp[ 0 +: 8];
            assign m_axi_wdata[48 +: 8] = m_axi_wdata_tmp[ 8 +: 8];
            assign m_axi_wdata[40 +: 8] = m_axi_wdata_tmp[16 +: 8];
            assign m_axi_wdata[32 +: 8] = m_axi_wdata_tmp[24 +: 8];
            assign m_axi_wdata[24 +: 8] = m_axi_wdata_tmp[32 +: 8];
            assign m_axi_wdata[16 +: 8] = m_axi_wdata_tmp[40 +: 8];
            assign m_axi_wdata[ 8 +: 8] = m_axi_wdata_tmp[48 +: 8];
            assign m_axi_wdata[ 0 +: 8] = m_axi_wdata_tmp[56 +: 8];
        end else begin
            assign m_axi_wdata = m_axi_wdata_tmp;
        end
    endgenerate
    assign m_axi_ar_go = m_axi_arvalid && m_axi_arready;
    assign m_axi_w_go  = m_axi_wvalid & m_axi_wready;
    assign m_axi_aw_go = m_axi_awvalid & m_axi_awready;
    
    always @( * ) begin
        m_axi_rready = (r_resp_buf_status_f == BUF_STATUS_WAITRESP);
        m_axi_bready = (w_resp_buf_status == BUF_STATUS_WAITRESP);
    end
    
    assign r_resp_buf_header0_next[63:50] = r_req_buf_header2_f[63:50];
    assign r_resp_buf_header0_next[49:42]      = r_req_buf_header2_f[49:42];
    assign r_resp_buf_header0_next[41:34]      = r_req_buf_header2_f[41:34];
    assign r_resp_buf_header0_next[33:30]  = r_req_buf_header2_f[33:30]; 
    assign r_resp_buf_header0_next[29:22]     = (r_req_buf_header0_f[21:14] == 8'd14 &&
                                                       r_req_buf_header1_f[10:8] <= 3'b100) ? 8'd1 :
                                                       8'd8; 
    assign r_resp_buf_header0_next[21:14]       = (r_req_buf_header0_f[21:14] == 8'd14) ? 8'd26 :
                                                      (r_req_buf_header0_f[21:14] == 8'd19) ? 8'd24 :
                                                      8'dx;
    assign r_resp_buf_header0_next[13:6]     = r_req_buf_header0_f[13:6];
    assign r_resp_buf_header0_next[5:0]  = 6'd0; 
    assign w_resp_buf_header0_next[63:50] = w_req_buf_header2_f[63:50];
    assign w_resp_buf_header0_next[49:42]      = w_req_buf_header2_f[49:42];
    assign w_resp_buf_header0_next[41:34]      = w_req_buf_header2_f[41:34];
    assign w_resp_buf_header0_next[33:30]  = w_req_buf_header2_f[33:30]; 
    assign w_resp_buf_header0_next[29:22]     = 8'd0;
    assign w_resp_buf_header0_next[21:14]       = (w_req_buf_header0_f[21:14] == 8'd15) ? 8'd27 :
                                                      (w_req_buf_header0_f[21:14] == 8'd20) ? 8'd25 :
                                                      8'dx;
    assign w_resp_buf_header0_next[13:6]     = w_req_buf_header0_f[13:6];
    assign w_resp_buf_header0_next[5:0]  = 6'd0; 
    
    assign m_axi_b_go = m_axi_bready && m_axi_bvalid;
    assign m_axi_r_go = m_axi_rready && m_axi_rvalid;
    
    generate
      if (ALIGN_RDATA) begin
        always @( * ) begin
            a_axi_rdata_shifted = (m_axi_rdata >> {m_axi_araddr[2:0], 3'b000});
        end
      end else begin
        always @( * ) begin
            a_axi_rdata_shifted = m_axi_rdata;
        end
      end
    endgenerate
    
    reg  [64-1:0]   a_axi_rdata_masked_tmp;
    generate
      if (SLAVE_RESP_BYTEWIDTH <= 0) begin
        
        always @( * ) begin
            case (r_req_buf_header1_f[10:8])
                3'b000: begin
                    a_axi_rdata_masked_tmp = {8{8'd0}};
                    r_reqbuf_size          = 3'b00;
                end
                3'b001: begin
                    a_axi_rdata_masked_tmp = {8{a_axi_rdata_shifted[7:0]}};
                    r_reqbuf_size          = 3'b00;
                end
                3'b010: begin
                    a_axi_rdata_masked_tmp = {4{a_axi_rdata_shifted[15:0]}};
                    r_reqbuf_size          = 3'b01;
                end
                3'b011: begin
                    a_axi_rdata_masked_tmp = {2{a_axi_rdata_shifted[31:0]}};
                    r_reqbuf_size          = 3'b10;
                end
                3'b100: begin
                    a_axi_rdata_masked_tmp = a_axi_rdata_shifted;
                    r_reqbuf_size          = 3'b11;
                end
                default: begin
                    a_axi_rdata_masked_tmp = a_axi_rdata_shifted;
                    r_reqbuf_size          = 3'b11;
                end
            endcase
        end
      end else if (SLAVE_RESP_BYTEWIDTH == 1) begin
          always @( * ) begin
              a_axi_rdata_masked_tmp = {8{m_axi_rdata[7:0]}};
              r_reqbuf_size          = 3'b00;
          end
      end else if (SLAVE_RESP_BYTEWIDTH == 2) begin
          always @( * ) begin
              a_axi_rdata_masked_tmp = {4{m_axi_rdata[15:0]}};
              r_reqbuf_size          = 3'b01;
          end
      end else if (SLAVE_RESP_BYTEWIDTH == 4) begin
          always @( * ) begin
              a_axi_rdata_masked_tmp = {2{m_axi_rdata[31:0]}};
              r_reqbuf_size          = 3'b10;
          end
      end else if (SLAVE_RESP_BYTEWIDTH == 8) begin
          always @( * ) begin
              a_axi_rdata_masked_tmp = m_axi_rdata;
              r_reqbuf_size          = 3'b11;
          end
      end else begin
          always @( * ) begin
              a_axi_rdata_masked_tmp = m_axi_rdata;
              r_reqbuf_size          = 3'b11;
          end
      end
    endgenerate
    generate
        if (SWAP_ENDIANESS) begin
            assign a_axi_rdata_masked[56 +: 8] = a_axi_rdata_masked_tmp[ 0 +: 8];
            assign a_axi_rdata_masked[48 +: 8] = a_axi_rdata_masked_tmp[ 8 +: 8];
            assign a_axi_rdata_masked[40 +: 8] = a_axi_rdata_masked_tmp[16 +: 8];
            assign a_axi_rdata_masked[32 +: 8] = a_axi_rdata_masked_tmp[24 +: 8];
            assign a_axi_rdata_masked[24 +: 8] = a_axi_rdata_masked_tmp[32 +: 8];
            assign a_axi_rdata_masked[16 +: 8] = a_axi_rdata_masked_tmp[40 +: 8];
            assign a_axi_rdata_masked[ 8 +: 8] = a_axi_rdata_masked_tmp[48 +: 8];
            assign a_axi_rdata_masked[ 0 +: 8] = a_axi_rdata_masked_tmp[56 +: 8];
        end else begin
            assign a_axi_rdata_masked = a_axi_rdata_masked_tmp;
        end
    endgenerate
    
    
    
    always @(posedge clk) begin
        if (rst) begin
            w_resp_buf_header0_f     <=  {64{1'b0}};
            w_resp_buf_bresp_f       <=  {2{1'b0}};
            w_addr_resp_buf_status_f <=  BUF_STATUS_INCOMP;
            w_data_resp_buf_status_f <=  BUF_STATUS_INCOMP;
        end
        else begin
            w_resp_buf_header0_f     <=  m_axi_aw_go              ? w_resp_buf_header0_next  :
                                                                    w_resp_buf_header0_f     ;
            w_resp_buf_bresp_f       <=  m_axi_b_go               ? m_axi_bresp              :
                                                                    w_resp_buf_bresp_f       ;
            w_addr_resp_buf_status_f <=  m_axi_aw_go              ? BUF_STATUS_WAITRESP      :
                                         m_axi_b_go               ? BUF_STATUS_RESPSEND      :
                                         io_splitter_ack_store_go ? BUF_STATUS_INCOMP        :
                                                                    w_addr_resp_buf_status_f ;
            w_data_resp_buf_status_f <=  m_axi_w_go               ? BUF_STATUS_WAITRESP      :
                                         m_axi_b_go               ? BUF_STATUS_RESPSEND      :
                                         io_splitter_ack_store_go ? BUF_STATUS_INCOMP        :
                                                                    w_data_resp_buf_status_f ;
        end
    end
    
    assign w_resp_buf_status =
        ((w_addr_resp_buf_status_f == BUF_STATUS_INCOMP  ) ||
         (w_data_resp_buf_status_f == BUF_STATUS_INCOMP  )    ) ? BUF_STATUS_INCOMP   :
        ((w_addr_resp_buf_status_f == BUF_STATUS_COMP    ) ||
         (w_data_resp_buf_status_f == BUF_STATUS_COMP    )    ) ? BUF_STATUS_COMP     :
        ((w_addr_resp_buf_status_f == BUF_STATUS_WAITRESP) ||
         (w_data_resp_buf_status_f == BUF_STATUS_WAITRESP)    ) ? BUF_STATUS_WAITRESP :
                                                                  BUF_STATUS_RESPSEND ;
    
    
    
    always @(posedge clk) begin
        if (rst) begin
            r_resp_buf_header0_f <= {64{1'b0}};
            r_resp_buf_data0_f   <= {64{1'b0}};
            r_resp_buf_rresp_f   <= {2{1'b0}};
            r_resp_buf_status_f  <= BUF_STATUS_INCOMP;
        end
        else begin
            r_resp_buf_header0_f <= m_axi_ar_go                                        ? r_resp_buf_header0_next :
                                                                                         r_resp_buf_header0_f    ;
            r_resp_buf_data0_f   <= m_axi_r_go                                         ? a_axi_rdata_masked      :
                                                                                         r_resp_buf_data0_f      ;
            r_resp_buf_rresp_f   <= m_axi_r_go                                         ? m_axi_rresp             :
                                                                                         r_resp_buf_rresp_f      ;
            r_resp_buf_status_f  <= m_axi_ar_go                                        ? BUF_STATUS_WAITRESP     :
                                    m_axi_r_go                                         ? BUF_STATUS_RESPSEND     :
                                    (io_splitter_ack_load_go                       &
                                     (io_splitter_ack_load_counter_f == 0)         &
                                     ~(r_resp_buf_status_f == BUF_STATUS_WAITRESP)   ) ? BUF_STATUS_INCOMP       :
                                                                                         r_resp_buf_status_f     ;
        end
    end
    assign  r_resp_buf_val = (r_resp_buf_status_f == BUF_STATUS_RESPSEND);
    assign  w_resp_buf_val = (w_resp_buf_status == BUF_STATUS_RESPSEND);
    assign  io_splitter_ack_store = w_resp_buf_header0_f;
    assign  io_splitter_ack_load = (io_splitter_ack_load_counter_f == r_resp_buf_header0_f[29:22]) ? r_resp_buf_header0_f
                                                       : r_resp_buf_data0_f;
    assign  io_splitter_ack_load_go = (io_splitter_ack_mux_sel == LOAD_ACK) && (r_resp_buf_val) && splitter_bridge_rdy;
    assign  io_splitter_ack_store_go = (io_splitter_ack_mux_sel == STORE_ACK) && (w_resp_buf_val) && splitter_bridge_rdy;
    always @( * ) begin
        
        if (io_splitter_ack_mux_sel == LOAD_ACK) begin
            bridge_splitter_val = r_resp_buf_val;
            bridge_splitter_data = io_splitter_ack_load;
        end
        else begin
            bridge_splitter_val = w_resp_buf_val;
            bridge_splitter_data = io_splitter_ack_store;
        end
    end
    
    always @( * ) begin
        if (r_resp_buf_val && (!w_resp_buf_val)) begin
            io_splitter_ack_mux_sel = LOAD_ACK;
        end
        else if (w_resp_buf_val && (!r_resp_buf_val)) begin
            io_splitter_ack_mux_sel = STORE_ACK;
        end
        else if (w_resp_buf_val && r_resp_buf_val) begin
            if(io_splitter_ack_load_counter_f == r_resp_buf_header0_f[29:22]) begin
                io_splitter_ack_mux_sel = io_splitter_arb_f;
            end
            else begin
                io_splitter_ack_mux_sel = LOAD_ACK;
            end
        end
        else begin
            io_splitter_ack_mux_sel = LOAD_ACK;
        end
    end
    
    always @(posedge clk) begin
        if (rst) begin
                io_splitter_arb_f <= 0;
                io_splitter_ack_load_counter_f <= 0;
        end
        else begin
            
            if (w_resp_buf_val && r_resp_buf_val && io_splitter_ack_load_go) begin
                io_splitter_arb_f <= STORE_ACK;
            end
            else if (w_resp_buf_val && r_resp_buf_val && io_splitter_ack_store_go) begin
                io_splitter_arb_f <= LOAD_ACK;
            end
            
            if (r_resp_buf_status_f == BUF_STATUS_WAITRESP) begin
                io_splitter_ack_load_counter_f <= r_resp_buf_header0_f[29:22];
            end
            else if(io_splitter_ack_load_go) begin
                if (io_splitter_ack_load_counter_f != 0) begin
                    io_splitter_ack_load_counter_f <= io_splitter_ack_load_counter_f - 1;
                end
            end
        end
    end
    assign bridge_splitter_rdy =
        ((splitter_io_msg_type_next == MSG_TYPE_INVAL) ||
         (splitter_io_msg_is_load_next && (r_req_buf_status_f == BUF_STATUS_INCOMP)) ||
         (splitter_io_msg_is_store_next && (w_req_buf_status == BUF_STATUS_INCOMP)));
endmodule
module blinker (
    input           clk,
    input           rst_n,
    output reg      GPIO_LED_0,
    output reg      GPIO_LED_1,
    output reg      GPIO_LED_2,
    output reg      GPIO_LED_3,
    output reg      GPIO_LED_4,
    output reg      GPIO_LED_5,
    output reg      GPIO_LED_6
 );
reg [31:0]              cnt;
reg                     out_val;
wire                    flag_0, flag_1, flag_2, flag_3;
always @(posedge clk) begin
        if (~rst_n)
                cnt <= 32'b0;
        else
                cnt <= cnt + 1;
end
always @(posedge clk) begin
        if (~rst_n) begin
                GPIO_LED_0 <= 1'b0;
                     GPIO_LED_1 <= 1'b0;
                     GPIO_LED_2 <= 1'b0;
                     GPIO_LED_3 <= 1'b0;
          end
        else begin
                GPIO_LED_0 <= flag_0 ? ~GPIO_LED_0 : GPIO_LED_0;
                     GPIO_LED_1 <= flag_1 ? ~GPIO_LED_1 : GPIO_LED_1;
                     GPIO_LED_2 <= flag_2 ? ~GPIO_LED_2 : GPIO_LED_2;
                     GPIO_LED_3 <= flag_3 ? ~GPIO_LED_3 : GPIO_LED_3;
          end
end
assign flag_0 = (cnt % 32'h100000)  == 32'b0;
assign flag_1 = (cnt % 32'h200000)  == 32'b0;
assign flag_2 = (cnt % 32'h300000)  == 32'b0;
assign flag_3 = (cnt % 32'h400000)  == 32'b0;
always @(*) begin
    GPIO_LED_4 = 1'b1;
    GPIO_LED_5 = 1'b0;
    GPIO_LED_6 = 1'b1;
end
endmodule
    
    
 
    
    
    
    
    
    
 
 
 
  
    
 
 
    
    
    
    
    
    
    
 
 
    
    
    
     
    
    
    
    
    
    
    
    
    
    
    
    
   
    
   
    
       
        
        
    
  
   
     
    
   
   
    
    
module chipset(
    input sys_clk,
    
    
    
     
    
    
     
    
    
     
     
    
     
 
 
  
 
    
    
        input                                   io_clk,
     
     
 
    
    input                                       rst_n,
    
    input                                       piton_ready_n,
    input                                       piton_prsnt_n,
    output                                      chipset_prsnt_n,
  
    
    
    
    
    
    
    
    
 
    
    output [31:0]                               intf_chip_data,
    output [1:0]                                intf_chip_channel,
    input  [2:0]                                intf_chip_credit_back,
    input  [31:0]                               chip_intf_data,
    input  [1:0]                                chip_intf_channel,
    output [2:0]                                chip_intf_credit_back,
 
    
    
    
 
 
 
    input                                        mc_clk,
    
    output wire [6     -1:0]    m_axi_awid,
    output wire [64   -1:0]    m_axi_awaddr,
    output wire [8    -1:0]    m_axi_awlen,
    output wire [3   -1:0]    m_axi_awsize,
    output wire [2  -1:0]    m_axi_awburst,
    output wire                                  m_axi_awlock,
    output wire [4  -1:0]    m_axi_awcache,
    output wire [3   -1:0]    m_axi_awprot,
    output wire [4    -1:0]    m_axi_awqos,
    output wire [4 -1:0]    m_axi_awregion,
    output wire [11   -1:0]    m_axi_awuser,
    output wire                                  m_axi_awvalid,
    input  wire                                  m_axi_awready,
    
    output wire  [6     -1:0]    m_axi_wid,
    output wire  [512   -1:0]    m_axi_wdata,
    output wire  [64   -1:0]    m_axi_wstrb,
    output wire                                   m_axi_wlast,
    output wire  [11   -1:0]    m_axi_wuser,
    output wire                                   m_axi_wvalid,
    input  wire                                   m_axi_wready,
    
    output wire  [6     -1:0]    m_axi_arid,
    output wire  [64   -1:0]    m_axi_araddr,
    output wire  [8    -1:0]    m_axi_arlen,
    output wire  [3   -1:0]    m_axi_arsize,
    output wire  [2  -1:0]    m_axi_arburst,
    output wire                                   m_axi_arlock,
    output wire  [4  -1:0]    m_axi_arcache,
    output wire  [3   -1:0]    m_axi_arprot,
    output wire  [4    -1:0]    m_axi_arqos,
    output wire  [4 -1:0]    m_axi_arregion,
    output wire  [11   -1:0]    m_axi_aruser,
    output wire                                   m_axi_arvalid,
    input  wire                                   m_axi_arready,
    
    input  wire  [6     -1:0]    m_axi_rid,
    input  wire  [512   -1:0]    m_axi_rdata,
    input  wire  [2   -1:0]    m_axi_rresp,
    input  wire                                   m_axi_rlast,
    input  wire  [11   -1:0]    m_axi_ruser,
    input  wire                                   m_axi_rvalid,
    output wire                                   m_axi_rready,
    
    input  wire  [6     -1:0]    m_axi_bid,
    input  wire  [2   -1:0]    m_axi_bresp,
    input  wire  [11   -1:0]    m_axi_buser,
    input  wire                                   m_axi_bvalid,
    output wire                                   m_axi_bready,
    input  wire                                   ddr_ready,
 
 
 
    
        
            
            
         
        
        
     
    
        
        
        
        
     
    
     
 
 
   
    
    
               
    
    
    
    
    
    
        
    
    
    
    
    
     
    
        input [31:0]  ext_irq,
        input [31:0] ext_irq_trigger
     
  
    ,
    
    output                                      ndmreset_o,    
    output                                      dmactive_o,    
    output  [1-1:0]                    debug_req_o,   
    input   [1-1:0]                    unavailable_i, 
    
    input                                       tck_i,
    input                                       tms_i,
    input                                       trst_ni,
    input                                       td_i,
    output                                      td_o,
    output                                      tdo_oe_o,
    
    input                                       rtc_i,         
    output  [1-1:0]                    timer_irq_o,   
    output  [1-1:0]                    ipi_o,         
    
    output  [1*2-1:0]                  irq_o          
);
  
 
wire                                            clk_locked;
reg                                             rst_n_rect;
reg                                             chipset_rst_n;
reg                                             chipset_rst_n_f;
reg                                             chipset_rst_n_ff;
wire                                            uart_boot_en;
wire                                            uart_timeout_en;
wire  [3:0]                                     noc_power_test_hop_count;
wire  [64-1:0]                     fpga_intf_data_noc1;
wire  [64-1:0]                     fpga_intf_data_noc2;
wire  [64-1:0]                     fpga_intf_data_noc3;
wire                                            fpga_intf_val_noc1;
wire                                            fpga_intf_val_noc2;
wire                                            fpga_intf_val_noc3;
wire                                            fpga_intf_rdy_noc1;
wire                                            fpga_intf_rdy_noc2;
wire                                            fpga_intf_rdy_noc3;
wire  [64-1:0]                     intf_fpga_data_noc1;
wire  [64-1:0]                     intf_fpga_data_noc2;
wire  [64-1:0]                     intf_fpga_data_noc3;
wire                                            intf_fpga_val_noc1;
wire                                            intf_fpga_val_noc2;
wire                                            intf_fpga_val_noc3;
wire                                            intf_fpga_rdy_noc1;
wire                                            intf_fpga_rdy_noc2;
wire                                            intf_fpga_rdy_noc3;
wire                                            processor_offchip_noc1_valid;
wire  [64-1:0]                     processor_offchip_noc1_data;
wire                                            processor_offchip_noc1_yummy;
wire                                            processor_offchip_noc2_valid;
wire  [64-1:0]                     processor_offchip_noc2_data;
wire                                            processor_offchip_noc2_yummy;
wire                                            processor_offchip_noc3_valid;
wire  [64-1:0]                     processor_offchip_noc3_data;
wire                                            processor_offchip_noc3_yummy;
wire                                            offchip_processor_noc1_valid;
wire  [64-1:0]                     offchip_processor_noc1_data;
wire                                            offchip_processor_noc1_yummy;
wire                                            offchip_processor_noc2_valid;
wire  [64-1:0]                     offchip_processor_noc2_data;
wire                                            offchip_processor_noc2_yummy;
wire                                            offchip_processor_noc3_valid;
wire  [64-1:0]                     offchip_processor_noc3_data;
wire                                            offchip_processor_noc3_yummy;
 
wire  [64-1:0]                     chipset_intf_data_noc1;
wire  [64-1:0]                     chipset_intf_data_noc2;
wire  [64-1:0]                     chipset_intf_data_noc3;
wire                                            chipset_intf_val_noc1;
wire                                            chipset_intf_val_noc2;
wire                                            chipset_intf_val_noc3;
wire                                            chipset_intf_rdy_noc1;
wire                                            chipset_intf_rdy_noc2;
wire                                            chipset_intf_rdy_noc3;
wire  [64-1:0]                     intf_chipset_data_noc1;
wire  [64-1:0]                     intf_chipset_data_noc2;
wire  [64-1:0]                     intf_chipset_data_noc3;
wire                                            intf_chipset_val_noc1;
wire                                            intf_chipset_val_noc2;
wire                                            intf_chipset_val_noc3;
wire                                            intf_chipset_rdy_noc1;
wire                                            intf_chipset_rdy_noc2;
wire                                            intf_chipset_rdy_noc3;
wire                                            init_calib_complete;
wire                                        test_start;
wire            net_phy_clk_inter;
wire            net_axi_clk;
wire            net_phy_txctl_inter;
wire    [3:0]   net_phy_txd_inter;
wire            net_phy_rxc_ibufg_out;
wire            net_phy_rxc_inter;
wire            net_phy_rxc_delayed;
reg             net_phy_rx_dv_f;
reg             net_phy_rx_err_f;
reg             net_phy_rx_dv_ff;
reg             net_phy_rx_err_ff;
wire            net_phy_rx_dv_inter;
wire            net_phy_rx_err_inter;
reg     [3:0]   net_phy_rxd_f;
reg     [3:0]   net_phy_rxd_ff;
wire    [3:0]   net_phy_rxd_inter;
wire            sd_clk_out_internal;
wire            invalid_access;
always @ (posedge chipset_clk)
begin
    chipset_rst_n_f <= chipset_rst_n;
    chipset_rst_n_ff <= chipset_rst_n_f;
end
  
    
        assign io_clk_loopback = io_clk;
    
    
     
 
always @ *
begin
 
    rst_n_rect = rst_n;
 
    
    chipset_rst_n = rst_n_rect & clk_locked & (~piton_prsnt_n);
 
  
end
    assign clk_locked = 1'b1;
 
    assign chipset_prsnt_n = ~rst_n_rect | ~clk_locked | ~test_start;
  
    
        
            
            
            
            
                
         
     
 
    
    
    
    
        
 
    
        
            
            
             
        
         
    
     
  
 
    assign uart_boot_en = 1'b0;
    assign uart_timeout_en = 1'b0;
    assign noc_power_test_hop_count = 4'b0;
 
    
        
            
            
            
            
            
             
             
            
             
            
            
             
            
            
         
     
        assign clk_locked = 1'b1;
        assign chipset_clk = sys_clk;
     
 
    
    
    
    
 
  
fpga_bridge
#(.SEND_CREDIT_THRESHOLD(9'd7))
 
fpga_bridge(
    
    .rst_n              (chipset_rst_n          ),
    .fpga_out_clk       (chipset_clk            ),
    .fpga_in_clk        (chipset_clk            ),
    
     
        .intf_out_clk   (io_clk_loopback        ),
        .intf_in_clk    (io_clk_loopback        ),
     
    .fpga_intf_data_noc1(fpga_intf_data_noc1),
    .fpga_intf_data_noc2(fpga_intf_data_noc2),
    .fpga_intf_data_noc3(fpga_intf_data_noc3),
    .fpga_intf_val_noc1(fpga_intf_val_noc1),
    .fpga_intf_val_noc2(fpga_intf_val_noc2),
    .fpga_intf_val_noc3(fpga_intf_val_noc3),
    .fpga_intf_rdy_noc1(fpga_intf_rdy_noc1),
    .fpga_intf_rdy_noc2(fpga_intf_rdy_noc2),
    .fpga_intf_rdy_noc3(fpga_intf_rdy_noc3),
    .fpga_intf_data(intf_chip_data),
    .fpga_intf_channel(intf_chip_channel),
    .fpga_intf_credit_back(intf_chip_credit_back),
    .intf_fpga_data_noc1(intf_fpga_data_noc1),
    .intf_fpga_data_noc2(intf_fpga_data_noc2),
    .intf_fpga_data_noc3(intf_fpga_data_noc3),
    .intf_fpga_val_noc1(intf_fpga_val_noc1),
    .intf_fpga_val_noc2(intf_fpga_val_noc2),
    .intf_fpga_val_noc3(intf_fpga_val_noc3),
    .intf_fpga_rdy_noc1(intf_fpga_rdy_noc1),
    .intf_fpga_rdy_noc2(intf_fpga_rdy_noc2),
    .intf_fpga_rdy_noc3(intf_fpga_rdy_noc3),
    .intf_fpga_data(chip_intf_data),
    .intf_fpga_channel(chip_intf_channel),
    .intf_fpga_credit_back(chip_intf_credit_back)
);
credit_to_valrdy offchip_processor_noc1_c2v(
    .clk(chipset_clk),
    .reset(~chipset_rst_n_ff),
    .data_in(offchip_processor_noc1_data),
    .valid_in(offchip_processor_noc1_valid),
    .yummy_in(offchip_processor_noc1_yummy),
    .data_out(fpga_intf_data_noc1),
    .valid_out(fpga_intf_val_noc1),
    .ready_out(fpga_intf_rdy_noc1)
);
credit_to_valrdy offchip_processor_noc2_c2v(
    .clk(chipset_clk),
    .reset(~chipset_rst_n_ff),
    .data_in(offchip_processor_noc2_data),
    .valid_in(offchip_processor_noc2_valid),
    .yummy_in(offchip_processor_noc2_yummy),
    .data_out(fpga_intf_data_noc2),
    .valid_out(fpga_intf_val_noc2),
    .ready_out(fpga_intf_rdy_noc2)
);
credit_to_valrdy offchip_processor_noc3_c2v(
    .clk(chipset_clk),
    .reset(~chipset_rst_n_ff),
    .data_in(offchip_processor_noc3_data),
    .valid_in(offchip_processor_noc3_valid),
    .yummy_in(offchip_processor_noc3_yummy),
    .data_out(fpga_intf_data_noc3),
    .valid_out(fpga_intf_val_noc3),
    .ready_out(fpga_intf_rdy_noc3)
);
valrdy_to_credit #(4, 3) processor_offchip_noc1_v2c(
    .clk(chipset_clk),
    .reset(~chipset_rst_n_ff),
    .data_in(intf_fpga_data_noc1),
    .valid_in(intf_fpga_val_noc1),
    .ready_in(intf_fpga_rdy_noc1),
    .data_out(processor_offchip_noc1_data),
    .valid_out(processor_offchip_noc1_valid),
    .yummy_out(processor_offchip_noc1_yummy)
);
valrdy_to_credit #(4, 3) processor_offchip_noc2_v2c(
    .clk(chipset_clk),
    .reset(~chipset_rst_n_ff),
    .data_in(intf_fpga_data_noc2),
    .valid_in(intf_fpga_val_noc2),
    .ready_in(intf_fpga_rdy_noc2),
    .data_out(processor_offchip_noc2_data),
    .valid_out(processor_offchip_noc2_valid),
    .yummy_out(processor_offchip_noc2_yummy)
);
valrdy_to_credit #(4, 3) processor_offchip_noc3_v2c(
    .clk(chipset_clk),
    .reset(~chipset_rst_n_ff),
    .data_in(intf_fpga_data_noc3),
    .valid_in(intf_fpga_val_noc3),
    .ready_in(intf_fpga_rdy_noc3),
    .data_out(processor_offchip_noc3_data),
    .valid_out(processor_offchip_noc3_valid),
    .yummy_out(processor_offchip_noc3_yummy)
);
 
valrdy_to_credit #(4, 3) offchip_processor_noc1_v2c(
    .clk(chipset_clk),
    .reset(~chipset_rst_n_ff),
    .data_in(chipset_intf_data_noc1),
    .valid_in(chipset_intf_val_noc1),
    .ready_in(chipset_intf_rdy_noc1),
    .data_out(offchip_processor_noc1_data),
    .valid_out(offchip_processor_noc1_valid),
    .yummy_out(offchip_processor_noc1_yummy)
);
valrdy_to_credit #(4, 3) offchip_processor_noc2_v2c(
    .clk(chipset_clk),
    .reset(~chipset_rst_n_ff),
    .data_in(chipset_intf_data_noc2),
    .valid_in(chipset_intf_val_noc2),
    .ready_in(chipset_intf_rdy_noc2),
    .data_out(offchip_processor_noc2_data),
    .valid_out(offchip_processor_noc2_valid),
    .yummy_out(offchip_processor_noc2_yummy)
);
valrdy_to_credit #(4, 3) offchip_processor_noc3_v2c(
    .clk(chipset_clk),
    .reset(~chipset_rst_n_ff),
    .data_in(chipset_intf_data_noc3),
    .valid_in(chipset_intf_val_noc3),
    .ready_in(chipset_intf_rdy_noc3),
    .data_out(offchip_processor_noc3_data),
    .valid_out(offchip_processor_noc3_valid),
    .yummy_out(offchip_processor_noc3_yummy)
);
credit_to_valrdy processor_offchip_noc1_c2v(
    .clk(chipset_clk),
    .reset(~chipset_rst_n_ff),
    .data_in(processor_offchip_noc1_data),
    .valid_in(processor_offchip_noc1_valid),
    .yummy_in(processor_offchip_noc1_yummy),
    .data_out(intf_chipset_data_noc1),
    .valid_out(intf_chipset_val_noc1),
    .ready_out(intf_chipset_rdy_noc1)
);
credit_to_valrdy processor_offchip_noc2_c2v(
    .clk(chipset_clk),
    .reset(~chipset_rst_n_ff),
    .data_in(processor_offchip_noc2_data),
    .valid_in(processor_offchip_noc2_valid),
    .yummy_in(processor_offchip_noc2_yummy),
    .data_out(intf_chipset_data_noc2),
    .valid_out(intf_chipset_val_noc2),
    .ready_out(intf_chipset_rdy_noc2)
);
credit_to_valrdy processor_offchip_noc3_c2v(
    .clk(chipset_clk),
    .reset(~chipset_rst_n_ff),
    .data_in(processor_offchip_noc3_data),
    .valid_in(processor_offchip_noc3_valid),
    .yummy_in(processor_offchip_noc3_yummy),
    .data_out(intf_chipset_data_noc3),
    .valid_out(intf_chipset_val_noc3),
    .ready_out(intf_chipset_rdy_noc3)
);
  
chipset_impl    chipset_impl    (
    .chipset_clk        (chipset_clk        ),
    .chipset_rst_n      (chipset_rst_n_ff   ),
    .piton_ready_n      (piton_ready_n      ),
    .test_start         (test_start         ),
    .uart_rst_out_n     (uart_rst_out_n     ),
    .invalid_access_o   (invalid_access     ),
    
    
    
        
        
        
          
     
     
     
    .chipset_intf_data_noc1(chipset_intf_data_noc1),
    .chipset_intf_data_noc2(chipset_intf_data_noc2),
    .chipset_intf_data_noc3(chipset_intf_data_noc3),
    .chipset_intf_val_noc1(chipset_intf_val_noc1),
    .chipset_intf_val_noc2(chipset_intf_val_noc2),
    .chipset_intf_val_noc3(chipset_intf_val_noc3),
    .chipset_intf_rdy_noc1(chipset_intf_rdy_noc1),
    .chipset_intf_rdy_noc2(chipset_intf_rdy_noc2),
    .chipset_intf_rdy_noc3(chipset_intf_rdy_noc3),
    .intf_chipset_data_noc1(intf_chipset_data_noc1),
    .intf_chipset_data_noc2(intf_chipset_data_noc2),
    .intf_chipset_data_noc3(intf_chipset_data_noc3),
    .intf_chipset_val_noc1(intf_chipset_val_noc1),
    .intf_chipset_val_noc2(intf_chipset_val_noc2),
    .intf_chipset_val_noc3(intf_chipset_val_noc3),
    .intf_chipset_rdy_noc1(intf_chipset_rdy_noc1),
    .intf_chipset_rdy_noc2(intf_chipset_rdy_noc2),
    .intf_chipset_rdy_noc3(intf_chipset_rdy_noc3)
    
    
         
            ,
            .init_calib_complete(init_calib_complete),
            
                 
                
                
                
                 
            
                
                
                
             
                .mc_clk(mc_clk),
                
                .m_axi_awid(m_axi_awid),
                .m_axi_awaddr(m_axi_awaddr),
                .m_axi_awlen(m_axi_awlen),
                .m_axi_awsize(m_axi_awsize),
                .m_axi_awburst(m_axi_awburst),
                .m_axi_awlock(m_axi_awlock),
                .m_axi_awcache(m_axi_awcache),
                .m_axi_awprot(m_axi_awprot),
                .m_axi_awqos(m_axi_awqos),
                .m_axi_awregion(m_axi_awregion),
                .m_axi_awuser(m_axi_awuser),
                .m_axi_awvalid(m_axi_awvalid),
                .m_axi_awready(m_axi_awready),
                
                .m_axi_wid(m_axi_wid),
                .m_axi_wdata(m_axi_wdata),
                .m_axi_wstrb(m_axi_wstrb),
                .m_axi_wlast(m_axi_wlast),
                .m_axi_wuser(m_axi_wuser),
                .m_axi_wvalid(m_axi_wvalid),
                .m_axi_wready(m_axi_wready),
                
                .m_axi_arid(m_axi_arid),
                .m_axi_araddr(m_axi_araddr),
                .m_axi_arlen(m_axi_arlen),
                .m_axi_arsize(m_axi_arsize),
                .m_axi_arburst(m_axi_arburst),
                .m_axi_arlock(m_axi_arlock),
                .m_axi_arcache(m_axi_arcache),
                .m_axi_arprot(m_axi_arprot),
                .m_axi_arqos(m_axi_arqos),
                .m_axi_arregion(m_axi_arregion),
                .m_axi_aruser(m_axi_aruser),
                .m_axi_arvalid(m_axi_arvalid),
                .m_axi_arready(m_axi_arready),
                
                .m_axi_rid(m_axi_rid),
                .m_axi_rdata(m_axi_rdata),
                .m_axi_rresp(m_axi_rresp),
                .m_axi_rlast(m_axi_rlast),
                .m_axi_ruser(m_axi_ruser),
                .m_axi_rvalid(m_axi_rvalid),
                .m_axi_rready(m_axi_rready),
                
                .m_axi_bid(m_axi_bid),
                .m_axi_bresp(m_axi_bresp),
                .m_axi_buser(m_axi_buser),
                .m_axi_bvalid(m_axi_bvalid),
                .m_axi_bready(m_axi_bready), 
                .ddr_ready(ddr_ready)
             
         
     
    
        
            
             
         
        
            
            
            
            
            
            
         
            
             
     
    
        ,
        .ext_irq(ext_irq),
        .ext_irq_trigger(ext_irq_trigger)
     
    
        ,
        .ndmreset_o             ( ndmreset_o    ),
        .dmactive_o             ( dmactive_o    ),
        .debug_req_o            ( debug_req_o   ),
        .unavailable_i          ( unavailable_i ),
        .tck_i                  ( tck_i         ),
        .tms_i                  ( tms_i         ),
        .trst_ni                ( trst_ni       ),
        .td_i                   ( td_i          ),
        .td_o                   ( td_o          ),
        .tdo_oe_o               ( tdo_oe_o      ),
        .rtc_i                  ( rtc_i         ),
        .timer_irq_o            ( timer_irq_o   ),
        .ipi_o                  ( ipi_o         ),
        .irq_o                  ( irq_o         )
    
);
                    
     
    
    
    
    
    
    
  
endmodule
   
    
   
    
       
        
        
    
  
   
     
    
   
   
    
    
module test_end_checker(
    input clk,
    input rst_n,
    
    
    
    input                       src_checker_noc2_val,
    input [64-1:0] src_checker_noc2_data,
    input                       src_checker_noc2_rdy,
    input                       uart_boot_en,
    output                      test_good_end,
    output                      test_bad_end
);
    localparam IDLE = 2'b00;
    localparam TWOFLITS = 2'b01;
    localparam COUNTDOWN = 2'b10;
    reg [1:0] state_reg;
    reg [1:0] state_next;
    reg [8-1:0] num_flits_reg;
    reg [8-1:0] num_flits_next;
    reg test_good_end_reg;
    reg test_good_end_next;
    reg test_bad_end_reg;
    reg test_bad_end_next;
    reg future_good_end_reg;
    reg future_good_end_next;
    reg future_bad_end_reg;
    reg future_bad_end_next;
    assign test_good_end = test_good_end_reg;
    assign test_bad_end  = test_bad_end_reg;
    always @* begin
        case (state_reg)
        IDLE: begin
            test_good_end_next   = 1'b0;
            test_bad_end_next    = 1'b0;
            future_good_end_next = 1'b0;
            future_bad_end_next  = 1'b0;
            if (src_checker_noc2_val & src_checker_noc2_rdy) begin
                num_flits_next = src_checker_noc2_data[29:22];
                
                if (src_checker_noc2_data[29:22] == 8'b0) begin
                    state_next = IDLE;
                end
                else begin
                    state_next = TWOFLITS;
                end
            end
            else begin
                num_flits_next = num_flits_reg;
                state_next = IDLE;
            end
        end
        TWOFLITS: begin
            test_good_end_next   = 1'b0;
            test_bad_end_next    = 1'b0;
            future_good_end_next = 1'b0;
            future_bad_end_next  = 1'b0;
            
            if (src_checker_noc2_val & src_checker_noc2_rdy) begin
                num_flits_next = num_flits_reg - 8'b1;
                
                if (num_flits_reg == 8'b1) begin
                    
                    test_good_end_next = (src_checker_noc2_data[((16 + 40 - 1)):(16)] == 40'h8100000000) & uart_boot_en;
                    test_bad_end_next  = (src_checker_noc2_data[((16 + 40 - 1)):(16)] == 40'h8200000000) & uart_boot_en;
                    state_next = IDLE;
                end
                else begin
                    
                    future_good_end_next = (src_checker_noc2_data[((16 + 40 - 1)):(16)] == 40'h8100000000) & uart_boot_en;
                    future_bad_end_next  = (src_checker_noc2_data[((16 + 40 - 1)):(16)] == 40'h8200000000) & uart_boot_en;
                    state_next = COUNTDOWN;
                end
            end
            else begin
                num_flits_next = num_flits_reg;
                state_next = TWOFLITS;
            end
        end
        COUNTDOWN: begin
            test_good_end_next   = 1'b0;
            test_bad_end_next    = 1'b0;
            future_good_end_next = future_good_end_reg;
            future_bad_end_next  = future_bad_end_reg;
            if (src_checker_noc2_val & src_checker_noc2_rdy) begin
                num_flits_next = num_flits_reg - 8'b1;
                if (num_flits_reg == 8'b1) begin
                    test_good_end_next = future_good_end_reg;
                    test_bad_end_next  = future_bad_end_reg;
                    state_next = IDLE;
                end
                else begin
                    state_next = COUNTDOWN;
                end
            end
            else begin
                num_flits_next = num_flits_reg;
                state_next = COUNTDOWN;
            end
        end
        default: begin
            test_good_end_next   = 1'bx;
            test_bad_end_next    = 1'bx;
            future_good_end_next = 1'bx;
            future_bad_end_next  = 1'bx;
            num_flits_next = {8{1'bx}};
            state_next = 2'bxx;
        end
        endcase
    end
    always @(posedge clk) begin
        if (!rst_n) begin
            state_reg           <= 2'b0;
            num_flits_reg       <= 8'b0;
            test_good_end_reg   <= 1'b0;
            test_bad_end_reg    <= 1'b0;
            future_good_end_reg <= 1'b0;
            future_bad_end_reg  <= 1'b0;
        end
        else begin
            state_reg           <= state_next;
            num_flits_reg       <= num_flits_next;
            test_good_end_reg   <= test_good_end_next;
            test_bad_end_reg    <= test_bad_end_next;
            future_good_end_reg <= future_good_end_next;
            future_bad_end_reg  <= future_bad_end_next;
        end
    end
endmodule
module noc_bidir_afifo (
    input wire          clk_1,
    input wire          rst_1,
    
    input wire          clk_2,
    input wire          rst_2,
    
    
    input wire          flit_in_val_1,
    input wire [63:0]   flit_in_data_1,
    output wire         flit_in_rdy_1,
    output wire         flit_out_val_2,
    output wire [63:0]  flit_out_data_2,
    input wire          flit_out_rdy_2,
    
    
    input wire          flit_in_val_2,
    input wire [63:0]   flit_in_data_2,
    output wire         flit_in_rdy_2,
    output wire         flit_out_val_1,
    output wire [63:0]  flit_out_data_1,
    input wire          flit_out_rdy_1
);
wire fifo_recv_full;
wire fifo_recv_empty;
reg  fifo_recv_empty_reg;
wire fifo_send_full;
wire fifo_send_empty;
reg  fifo_send_empty_reg;
wire    [63:0]  fifo_data_to_splitter;
wire            fifo_recv_rd_en;
reg             outreg_empty;
 
assign flit_out_data_2 = flit_in_data_1;
assign flit_data_to_splitter = flit_in_data_2;
 
assign flit_in_rdy_1 = ~fifo_send_full;
assign flit_in_rdy_2 = ~fifo_recv_full;
always @ (posedge clk_1)
    fifo_recv_empty_reg <= fifo_recv_empty;
always @ (posedge clk_2)
begin
    if (rst_2)
    begin
        fifo_send_empty_reg <= 1'b1;
    end
    else
    begin
        if (flit_out_rdy_2)
        begin
            fifo_send_empty_reg <= fifo_send_empty;  
        end
        else
        begin
            fifo_send_empty_reg <= fifo_send_empty_reg;  
        end
    end
end
always @(posedge clk_1) begin
    if (rst_1)
        outreg_empty <= 1'b1;
    else
        outreg_empty <= fifo_recv_rd_en                                     ? 1'b0 :
                        ~outreg_empty & flit_out_rdy_1 & ~fifo_recv_rd_en   ? 1'b1 : outreg_empty;
end
assign fifo_recv_rd_en = ~fifo_recv_empty & (outreg_empty | (~outreg_empty & flit_out_rdy_1));
assign flit_out_val_1 = ~outreg_empty;
assign flit_out_data_1 = fifo_data_to_splitter;
assign flit_out_val_2 = ~fifo_send_empty_reg;
endmodule
    
    
 
    
    
    
    
    
    
 
 
 
  
    
 
 
    
    
    
    
    
    
    
 
 
    
    
    
     
    
    
    
    
    
    
    
    
    
    
    
    
         
         
   
    
   
    
       
        
        
    
  
   
     
    
   
   
    
    
module chipset_impl(
    
    input                                       chipset_clk,
    input                                       chipset_rst_n,
    input                                       piton_ready_n,
    output                                      test_start,
    output                                      uart_rst_out_n,
    
    output                                      invalid_access_o,
 
 
 
 
    
    output [64-1:0]                chipset_intf_data_noc1,
    output [64-1:0]                chipset_intf_data_noc2,
    output [64-1:0]                chipset_intf_data_noc3,
    output                                      chipset_intf_val_noc1,
    output                                      chipset_intf_val_noc2,
    output                                      chipset_intf_val_noc3,
    input                                       chipset_intf_rdy_noc1,
    input                                       chipset_intf_rdy_noc2,
    input                                       chipset_intf_rdy_noc3,
    input  [64-1:0]                intf_chipset_data_noc1,
    input  [64-1:0]                intf_chipset_data_noc2,
    input  [64-1:0]                intf_chipset_data_noc3,
    input                                       intf_chipset_val_noc1,
    input                                       intf_chipset_val_noc2,
    input                                       intf_chipset_val_noc3,
    output                                      intf_chipset_rdy_noc1,
    output                                      intf_chipset_rdy_noc2,
    output                                      intf_chipset_rdy_noc3
    
    ,
    output                                      init_calib_complete
    
    
 
 
 
    
    ,
    input                                        mc_clk,
    output wire [6     -1:0]    m_axi_awid,
    output wire [64   -1:0]    m_axi_awaddr,
    output wire [8    -1:0]    m_axi_awlen,
    output wire [3   -1:0]    m_axi_awsize,
    output wire [2  -1:0]    m_axi_awburst,
    output wire                                  m_axi_awlock,
    output wire [4  -1:0]    m_axi_awcache,
    output wire [3   -1:0]    m_axi_awprot,
    output wire [4    -1:0]    m_axi_awqos,
    output wire [4 -1:0]    m_axi_awregion,
    output wire [11   -1:0]    m_axi_awuser,
    output wire                                  m_axi_awvalid,
    input  wire                                  m_axi_awready,
    
    output wire  [6     -1:0]    m_axi_wid,
    output wire  [512   -1:0]    m_axi_wdata,
    output wire  [64   -1:0]    m_axi_wstrb,
    output wire                                   m_axi_wlast,
    output wire  [11   -1:0]    m_axi_wuser,
    output wire                                   m_axi_wvalid,
    input  wire                                   m_axi_wready,
    
    output wire  [6     -1:0]    m_axi_arid,
    output wire  [64   -1:0]    m_axi_araddr,
    output wire  [8    -1:0]    m_axi_arlen,
    output wire  [3   -1:0]    m_axi_arsize,
    output wire  [2  -1:0]    m_axi_arburst,
    output wire                                   m_axi_arlock,
    output wire  [4  -1:0]    m_axi_arcache,
    output wire  [3   -1:0]    m_axi_arprot,
    output wire  [4    -1:0]    m_axi_arqos,
    output wire  [4 -1:0]    m_axi_arregion,
    output wire  [11   -1:0]    m_axi_aruser,
    output wire                                   m_axi_arvalid,
    input  wire                                   m_axi_arready,
    
    input  wire  [6     -1:0]    m_axi_rid,
    input  wire  [512   -1:0]    m_axi_rdata,
    input  wire  [2   -1:0]    m_axi_rresp,
    input  wire                                   m_axi_rlast,
    input  wire  [11   -1:0]    m_axi_ruser,
    input  wire                                   m_axi_rvalid,
    output wire                                   m_axi_rready,
    
    input  wire  [6     -1:0]    m_axi_bid,
    input  wire  [2   -1:0]    m_axi_bresp,
    input  wire  [11   -1:0]    m_axi_buser,
    input  wire                                   m_axi_bvalid,
    output wire                                   m_axi_bready, 
    input  wire                                   ddr_ready
 
 
 
 
 
 
 
 
    
        ,
        input [31:0]  ext_irq,
        input [31:0] ext_irq_trigger
     
    ,
    
    output                                      ndmreset_o,    
    output                                      dmactive_o,    
    output [1-1:0]                     debug_req_o,   
    input  [1-1:0]                     unavailable_i, 
    
    input                                       tck_i,
    input                                       tms_i,
    input                                       trst_ni,
    input                                       td_i,
    output                                      td_o,
    output                                      tdo_oe_o,
    
    input                                       rtc_i,         
    output [1-1:0]                     timer_irq_o,   
    output [1-1:0]                     ipi_o,         
    
    output [1*2-1:0]                   irq_o          
);
wire                                            mc_ui_clk_sync_rst;
reg                                             init_calib_complete_f;
reg                                             init_calib_complete_ff;
reg                                             io_ctrl_rst_n;
 
wire                                            uart_boot_en;
wire                                            uart_timeout_en;
 
 
 
 
wire                                            cpu_mem_traffic;
wire                                            chip_filter_noc2_valid;
wire    [64-1:0]                   chip_filter_noc2_data;
wire                                            filter_chip_noc2_ready;
wire                                            filter_chip_noc3_valid;
wire    [64-1:0]                   filter_chip_noc3_data;
wire                                            chip_filter_noc3_ready;
wire                                            test_good_end;
wire                                            test_bad_end;
wire [64-1:0] chip_buf_xbar_noc2_data;
wire                   chip_buf_xbar_noc2_valid;
wire                   chip_buf_xbar_noc2_yummy;
wire [64-1:0] xbar_buf_chip_noc2_data;
wire                   xbar_buf_chip_noc2_valid;
wire                   xbar_buf_chip_noc2_yummy;
wire [64-1:0] buf_chip_noc2_data;
wire                   buf_chip_noc2_valid;
wire                   chip_buf_noc2_ready;
wire [64-1:0] chip_buf_noc2_data;
wire                   chip_buf_noc2_valid;
wire                   buf_chip_noc2_ready;
wire [64-1:0] chip_buf_xbar_noc3_data;
wire                   chip_buf_xbar_noc3_valid;
wire                   chip_buf_xbar_noc3_yummy;
wire [64-1:0] xbar_buf_chip_noc3_data;
wire                   xbar_buf_chip_noc3_valid;
wire                   xbar_buf_chip_noc3_yummy;
wire [64-1:0] buf_chip_noc3_data;
wire                   buf_chip_noc3_valid;
wire                   chip_buf_noc3_ready;
wire [64-1:0] chip_buf_noc3_data;
wire                   chip_buf_noc3_valid;
wire                   buf_chip_noc3_ready;
wire [64-1:0] mem_buf_xbar_noc2_data;
wire                   mem_buf_xbar_noc2_valid;
wire                   mem_buf_xbar_noc2_yummy;
wire [64-1:0] xbar_buf_mem_noc2_data;
wire                   xbar_buf_mem_noc2_valid;
wire                   xbar_buf_mem_noc2_yummy;
wire [64-1:0] buf_mem_noc2_data;
wire                   buf_mem_noc2_valid;
wire                   mem_buf_noc2_ready;
wire [64-1:0] mem_buf_noc2_data;
wire                   mem_buf_noc2_valid;
wire                   buf_mem_noc2_ready;
wire [64-1:0] mem_buf_xbar_noc3_data;
wire                   mem_buf_xbar_noc3_valid;
wire                   mem_buf_xbar_noc3_yummy;
wire [64-1:0] xbar_buf_mem_noc3_data;
wire                   xbar_buf_mem_noc3_valid;
wire                   xbar_buf_mem_noc3_yummy;
wire [64-1:0] buf_mem_noc3_data;
wire                   buf_mem_noc3_valid;
wire                   mem_buf_noc3_ready;
wire [64-1:0] mem_buf_noc3_data;
wire                   mem_buf_noc3_valid;
wire                   buf_mem_noc3_ready;
assign mem_buf_noc2_data = 64'b0;
assign mem_buf_noc2_valid = 1'b0;
assign mem_buf_noc3_ready = 1'b0;
wire [64-1:0] iob_buf_xbar_noc2_data;
wire                   iob_buf_xbar_noc2_valid;
wire                   iob_buf_xbar_noc2_yummy;
wire [64-1:0] xbar_buf_iob_noc2_data;
wire                   xbar_buf_iob_noc2_valid;
wire                   xbar_buf_iob_noc2_yummy;
wire [64-1:0] buf_iob_noc2_data;
wire                   buf_iob_noc2_valid;
wire                   iob_buf_noc2_ready;
wire [64-1:0] iob_buf_noc2_data;
wire                   iob_buf_noc2_valid;
wire                   buf_iob_noc2_ready;
wire [64-1:0] iob_buf_xbar_noc3_data;
wire                   iob_buf_xbar_noc3_valid;
wire                   iob_buf_xbar_noc3_yummy;
wire [64-1:0] xbar_buf_iob_noc3_data;
wire                   xbar_buf_iob_noc3_valid;
wire                   xbar_buf_iob_noc3_yummy;
wire [64-1:0] buf_iob_noc3_data;
wire                   buf_iob_noc3_valid;
wire                   iob_buf_noc3_ready;
wire [64-1:0] iob_buf_noc3_data;
wire                   iob_buf_noc3_valid;
wire                   buf_iob_noc3_ready;
wire [64-1:0]            iob_filter_noc2_data;
wire                              iob_filter_noc2_valid;
wire                              filter_iob_noc2_ready;
wire [64-1:0]             filter_iob_noc3_data;
wire                               filter_iob_noc3_valid;
wire                               iob_filter_noc3_ready;
wire [64-1:0] sd_buf_xbar_noc2_data;
wire                   sd_buf_xbar_noc2_valid;
wire                   sd_buf_xbar_noc2_yummy;
wire [64-1:0] xbar_buf_sd_noc2_data;
wire                   xbar_buf_sd_noc2_valid;
wire                   xbar_buf_sd_noc2_yummy;
wire [64-1:0] buf_sd_noc2_data;
wire                   buf_sd_noc2_valid;
wire                   sd_buf_noc2_ready;
wire [64-1:0] sd_buf_noc2_data;
wire                   sd_buf_noc2_valid;
wire                   buf_sd_noc2_ready;
wire [64-1:0] sd_buf_xbar_noc3_data;
wire                   sd_buf_xbar_noc3_valid;
wire                   sd_buf_xbar_noc3_yummy;
wire [64-1:0] xbar_buf_sd_noc3_data;
wire                   xbar_buf_sd_noc3_valid;
wire                   xbar_buf_sd_noc3_yummy;
wire [64-1:0] buf_sd_noc3_data;
wire                   buf_sd_noc3_valid;
wire                   sd_buf_noc3_ready;
wire [64-1:0] sd_buf_noc3_data;
wire                   sd_buf_noc3_valid;
wire                   buf_sd_noc3_ready;
assign sd_buf_noc2_data = 64'b0;
assign sd_buf_noc2_valid = 1'b0;
assign sd_buf_noc3_ready = 1'b0;
wire [64-1:0] uart_buf_xbar_noc2_data;
wire                   uart_buf_xbar_noc2_valid;
wire                   uart_buf_xbar_noc2_yummy;
wire [64-1:0] xbar_buf_uart_noc2_data;
wire                   xbar_buf_uart_noc2_valid;
wire                   xbar_buf_uart_noc2_yummy;
wire [64-1:0] buf_uart_noc2_data;
wire                   buf_uart_noc2_valid;
wire                   uart_buf_noc2_ready;
wire [64-1:0] uart_buf_noc2_data;
wire                   uart_buf_noc2_valid;
wire                   buf_uart_noc2_ready;
wire [64-1:0] uart_buf_xbar_noc3_data;
wire                   uart_buf_xbar_noc3_valid;
wire                   uart_buf_xbar_noc3_yummy;
wire [64-1:0] xbar_buf_uart_noc3_data;
wire                   xbar_buf_uart_noc3_valid;
wire                   xbar_buf_uart_noc3_yummy;
wire [64-1:0] buf_uart_noc3_data;
wire                   buf_uart_noc3_valid;
wire                   uart_buf_noc3_ready;
wire [64-1:0] uart_buf_noc3_data;
wire                   uart_buf_noc3_valid;
wire                   buf_uart_noc3_ready;
wire [64-1:0]            uart_filter_noc2_data;
wire                              uart_filter_noc2_valid;
wire                              filter_uart_noc2_ready;
wire [64-1:0]             filter_uart_noc3_data;
wire                               filter_uart_noc3_valid;
wire                               uart_filter_noc3_ready;
wire [64-1:0] net_buf_xbar_noc2_data;
wire                   net_buf_xbar_noc2_valid;
wire                   net_buf_xbar_noc2_yummy;
wire [64-1:0] xbar_buf_net_noc2_data;
wire                   xbar_buf_net_noc2_valid;
wire                   xbar_buf_net_noc2_yummy;
wire [64-1:0] buf_net_noc2_data;
wire                   buf_net_noc2_valid;
wire                   net_buf_noc2_ready;
wire [64-1:0] net_buf_noc2_data;
wire                   net_buf_noc2_valid;
wire                   buf_net_noc2_ready;
wire [64-1:0] net_buf_xbar_noc3_data;
wire                   net_buf_xbar_noc3_valid;
wire                   net_buf_xbar_noc3_yummy;
wire [64-1:0] xbar_buf_net_noc3_data;
wire                   xbar_buf_net_noc3_valid;
wire                   xbar_buf_net_noc3_yummy;
wire [64-1:0] buf_net_noc3_data;
wire                   buf_net_noc3_valid;
wire                   net_buf_noc3_ready;
wire [64-1:0] net_buf_noc3_data;
wire                   net_buf_noc3_valid;
wire                   buf_net_noc3_ready;
assign net_buf_noc2_data = 64'b0;
assign net_buf_noc2_valid = 1'b0;
assign net_buf_noc3_ready = 1'b0;
always @ (posedge chipset_clk)
begin
    init_calib_complete_f <= init_calib_complete;
    init_calib_complete_ff <= init_calib_complete_f;
end
 
 
 
assign chipset_intf_data_noc1 = {64{1'b0}};
assign chipset_intf_val_noc1 = 1'b0;
assign intf_chipset_rdy_noc3 = 1'b0;
assign chip_buf_noc3_valid = 1'b0;
assign chip_buf_noc3_data = {64{1'b0}};
 
 
    always @ *
    begin
    
    
        
        
        io_ctrl_rst_n = ~mc_ui_clk_sync_rst & init_calib_complete_ff;
    
     
    
     
    end
 
 
    
        assign uart_boot_en = 1'b0;
        assign uart_timeout_en = 1'b0;
     
        
         
     
 
    assign cpu_mem_traffic = test_start | (~uart_boot_en);
assign chipset_intf_val_noc2 = buf_chip_noc2_valid;
assign chipset_intf_data_noc2 = buf_chip_noc2_data;
assign chip_buf_noc2_ready = chipset_intf_rdy_noc2;
assign chip_filter_noc2_valid = intf_chipset_val_noc2;
assign chip_filter_noc2_data = intf_chipset_data_noc2;
assign intf_chipset_rdy_noc2    = filter_chip_noc2_ready & cpu_mem_traffic;
assign chipset_intf_val_noc3    = cpu_mem_traffic & filter_chip_noc3_valid;
assign chipset_intf_data_noc3   = filter_chip_noc3_data;
assign chip_filter_noc3_ready  = cpu_mem_traffic ? chipset_intf_rdy_noc3 : 1'b1;
    assign test_good_end = 1'b0;
    assign test_bad_end = 1'b0;
wire [3-1:0] invalid_access;
assign invalid_access_o = |invalid_access;
packet_filter chip_packet_filter(
    .clk(chipset_clk),
    .rst_n(chipset_rst_n),
    
    .invalid_access_o(invalid_access[0]),
    
    .noc2_filter_val(chip_filter_noc2_valid),
    .noc2_filter_data(chip_filter_noc2_data),
    .filter_noc2_rdy(filter_chip_noc2_ready),
    
    .filter_noc3_val(filter_chip_noc3_valid),
    .filter_noc3_data(filter_chip_noc3_data),
    .noc3_filter_rdy(chip_filter_noc3_ready),
    
    .filter_xbar_val(chip_buf_noc2_valid),
    .filter_xbar_data(chip_buf_noc2_data),
    .xbar_filter_rdy(buf_chip_noc2_ready),
    
    .xbar_filter_val(buf_chip_noc3_valid),
    .xbar_filter_data(buf_chip_noc3_data),
    .filter_xbar_rdy(chip_buf_noc3_ready),
    .uart_boot_en(uart_boot_en)
);
packet_filter iob_packet_filter(
    .clk(chipset_clk),
    .rst_n(chipset_rst_n),
    
    .invalid_access_o(invalid_access[1]),
    
    .noc2_filter_val(iob_filter_noc2_valid),
    .noc2_filter_data(iob_filter_noc2_data),
    .filter_noc2_rdy(filter_iob_noc2_ready),
    
    .filter_noc3_val(filter_iob_noc3_valid),
    .filter_noc3_data(filter_iob_noc3_data),
    .noc3_filter_rdy(iob_filter_noc3_ready),
    
    .filter_xbar_val(iob_buf_noc2_valid),
    .filter_xbar_data(iob_buf_noc2_data),
    .xbar_filter_rdy(buf_iob_noc2_ready),
    
    .xbar_filter_val(buf_iob_noc3_valid),
    .xbar_filter_data(buf_iob_noc3_data),
    .filter_xbar_rdy(iob_buf_noc3_ready),
    .uart_boot_en(uart_boot_en)
);
packet_filter uart_packet_filter(
    .clk(chipset_clk),
    .rst_n(chipset_rst_n),
    
    .invalid_access_o(invalid_access[2]),
    
    .noc2_filter_val(uart_filter_noc2_valid),
    .noc2_filter_data(uart_filter_noc2_data),
    .filter_noc2_rdy(filter_uart_noc2_ready),
    
    .filter_noc3_val(filter_uart_noc3_valid),
    .filter_noc3_data(filter_uart_noc3_data),
    .noc3_filter_rdy(uart_filter_noc3_ready),
    
    .filter_xbar_val(uart_buf_noc2_valid),
    .filter_xbar_data(uart_buf_noc2_data),
    .xbar_filter_rdy(buf_uart_noc2_ready),
    
    .xbar_filter_val(buf_uart_noc3_valid),
    .xbar_filter_data(buf_uart_noc3_data),
    .filter_xbar_rdy(uart_buf_noc3_ready),
    .uart_boot_en(uart_boot_en)
);
io_xbar_top_wrap io_xbar_noc2 (
    .clk                (chipset_clk),
    .reset_in           (~chipset_rst_n),
    .myChipID                   (14'b10000000000000),    
    .myLocX                     (8'b0),  
    .myLocY                     (8'b0),  
    .dataIn_0(chip_buf_xbar_noc2_data),
    .validIn_0(chip_buf_xbar_noc2_valid),
    .yummyIn_0(chip_buf_xbar_noc2_yummy),
    .dataOut_0(xbar_buf_chip_noc2_data),
    .validOut_0(xbar_buf_chip_noc2_valid),
    .yummyOut_0(xbar_buf_chip_noc2_yummy),
    .dataIn_1(mem_buf_xbar_noc2_data),
    .validIn_1(mem_buf_xbar_noc2_valid),
    .yummyIn_1(mem_buf_xbar_noc2_yummy),
    .dataOut_1(xbar_buf_mem_noc2_data),
    .validOut_1(xbar_buf_mem_noc2_valid),
    .yummyOut_1(xbar_buf_mem_noc2_yummy),
    .dataIn_2(iob_buf_xbar_noc2_data),
    .validIn_2(iob_buf_xbar_noc2_valid),
    .yummyIn_2(iob_buf_xbar_noc2_yummy),
    .dataOut_2(xbar_buf_iob_noc2_data),
    .validOut_2(xbar_buf_iob_noc2_valid),
    .yummyOut_2(xbar_buf_iob_noc2_yummy),
    .dataIn_3(sd_buf_xbar_noc2_data),
    .validIn_3(sd_buf_xbar_noc2_valid),
    .yummyIn_3(sd_buf_xbar_noc2_yummy),
    .dataOut_3(xbar_buf_sd_noc2_data),
    .validOut_3(xbar_buf_sd_noc2_valid),
    .yummyOut_3(xbar_buf_sd_noc2_yummy),
    .dataIn_4(uart_buf_xbar_noc2_data),
    .validIn_4(uart_buf_xbar_noc2_valid),
    .yummyIn_4(uart_buf_xbar_noc2_yummy),
    .dataOut_4(xbar_buf_uart_noc2_data),
    .validOut_4(xbar_buf_uart_noc2_valid),
    .yummyOut_4(xbar_buf_uart_noc2_yummy),
    .dataIn_5(net_buf_xbar_noc2_data),
    .validIn_5(net_buf_xbar_noc2_valid),
    .yummyIn_5(net_buf_xbar_noc2_yummy),
    .dataOut_5(xbar_buf_net_noc2_data),
    .validOut_5(xbar_buf_net_noc2_valid),
    .yummyOut_5(xbar_buf_net_noc2_yummy)
);
io_xbar_top_wrap io_xbar_noc3 (
    .clk                (chipset_clk),
    .reset_in           (~chipset_rst_n),
    .myChipID                   (14'b10000000000000),    
    .myLocX                     (8'b0),  
    .myLocY                     (8'b0),  
    .dataIn_0(chip_buf_xbar_noc3_data),
    .validIn_0(chip_buf_xbar_noc3_valid),
    .yummyIn_0(chip_buf_xbar_noc3_yummy),
    .dataOut_0(xbar_buf_chip_noc3_data),
    .validOut_0(xbar_buf_chip_noc3_valid),
    .yummyOut_0(xbar_buf_chip_noc3_yummy),
    .dataIn_1(mem_buf_xbar_noc3_data),
    .validIn_1(mem_buf_xbar_noc3_valid),
    .yummyIn_1(mem_buf_xbar_noc3_yummy),
    .dataOut_1(xbar_buf_mem_noc3_data),
    .validOut_1(xbar_buf_mem_noc3_valid),
    .yummyOut_1(xbar_buf_mem_noc3_yummy),
    .dataIn_2(iob_buf_xbar_noc3_data),
    .validIn_2(iob_buf_xbar_noc3_valid),
    .yummyIn_2(iob_buf_xbar_noc3_yummy),
    .dataOut_2(xbar_buf_iob_noc3_data),
    .validOut_2(xbar_buf_iob_noc3_valid),
    .yummyOut_2(xbar_buf_iob_noc3_yummy),
    .dataIn_3(sd_buf_xbar_noc3_data),
    .validIn_3(sd_buf_xbar_noc3_valid),
    .yummyIn_3(sd_buf_xbar_noc3_yummy),
    .dataOut_3(xbar_buf_sd_noc3_data),
    .validOut_3(xbar_buf_sd_noc3_valid),
    .yummyOut_3(xbar_buf_sd_noc3_yummy),
    .dataIn_4(uart_buf_xbar_noc3_data),
    .validIn_4(uart_buf_xbar_noc3_valid),
    .yummyIn_4(uart_buf_xbar_noc3_yummy),
    .dataOut_4(xbar_buf_uart_noc3_data),
    .validOut_4(xbar_buf_uart_noc3_valid),
    .yummyOut_4(xbar_buf_uart_noc3_yummy),
    .dataIn_5(net_buf_xbar_noc3_data),
    .validIn_5(net_buf_xbar_noc3_valid),
    .yummyIn_5(net_buf_xbar_noc3_yummy),
    .dataOut_5(xbar_buf_net_noc3_data),
    .validOut_5(xbar_buf_net_noc3_valid),
    .yummyOut_5(xbar_buf_net_noc3_yummy)
    ,
    .thanksIn_5()
);
valrdy_to_credit noc2_chip_to_xbar (
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(chip_buf_noc2_data),
      .valid_in(chip_buf_noc2_valid),
      .ready_in(buf_chip_noc2_ready),
      .data_out(chip_buf_xbar_noc2_data),           
      .valid_out(chip_buf_xbar_noc2_valid),       
      .yummy_out(xbar_buf_chip_noc2_yummy)    
);
credit_to_valrdy noc2_xbar_to_chip(
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(xbar_buf_chip_noc2_data),
      .valid_in(xbar_buf_chip_noc2_valid),
      .yummy_in(chip_buf_xbar_noc2_yummy),
      .data_out(buf_chip_noc2_data),           
      .valid_out(buf_chip_noc2_valid),       
      .ready_out(chip_buf_noc2_ready)    
);
valrdy_to_credit noc3_chip_to_xbar (
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(chip_buf_noc3_data),
      .valid_in(chip_buf_noc3_valid),
      .ready_in(buf_chip_noc3_ready),
      .data_out(chip_buf_xbar_noc3_data),           
      .valid_out(chip_buf_xbar_noc3_valid),       
      .yummy_out(xbar_buf_chip_noc3_yummy)    
);
credit_to_valrdy noc3_xbar_to_chip(
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(xbar_buf_chip_noc3_data),
      .valid_in(xbar_buf_chip_noc3_valid),
      .yummy_in(chip_buf_xbar_noc3_yummy),
      .data_out(buf_chip_noc3_data),           
      .valid_out(buf_chip_noc3_valid),       
      .ready_out(chip_buf_noc3_ready)    
);
valrdy_to_credit noc2_mem_to_xbar (
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(mem_buf_noc2_data),
      .valid_in(mem_buf_noc2_valid),
      .ready_in(buf_mem_noc2_ready),
      .data_out(mem_buf_xbar_noc2_data),           
      .valid_out(mem_buf_xbar_noc2_valid),       
      .yummy_out(xbar_buf_mem_noc2_yummy)    
);
credit_to_valrdy noc2_xbar_to_mem(
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(xbar_buf_mem_noc2_data),
      .valid_in(xbar_buf_mem_noc2_valid),
      .yummy_in(mem_buf_xbar_noc2_yummy),
      .data_out(buf_mem_noc2_data),           
      .valid_out(buf_mem_noc2_valid),       
      .ready_out(mem_buf_noc2_ready)    
);
valrdy_to_credit noc3_mem_to_xbar (
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(mem_buf_noc3_data),
      .valid_in(mem_buf_noc3_valid),
      .ready_in(buf_mem_noc3_ready),
      .data_out(mem_buf_xbar_noc3_data),           
      .valid_out(mem_buf_xbar_noc3_valid),       
      .yummy_out(xbar_buf_mem_noc3_yummy)    
);
credit_to_valrdy noc3_xbar_to_mem(
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(xbar_buf_mem_noc3_data),
      .valid_in(xbar_buf_mem_noc3_valid),
      .yummy_in(mem_buf_xbar_noc3_yummy),
      .data_out(buf_mem_noc3_data),           
      .valid_out(buf_mem_noc3_valid),       
      .ready_out(mem_buf_noc3_ready)    
);
valrdy_to_credit noc2_iob_to_xbar (
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(iob_buf_noc2_data),
      .valid_in(iob_buf_noc2_valid),
      .ready_in(buf_iob_noc2_ready),
      .data_out(iob_buf_xbar_noc2_data),           
      .valid_out(iob_buf_xbar_noc2_valid),       
      .yummy_out(xbar_buf_iob_noc2_yummy)    
);
credit_to_valrdy noc2_xbar_to_iob(
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(xbar_buf_iob_noc2_data),
      .valid_in(xbar_buf_iob_noc2_valid),
      .yummy_in(iob_buf_xbar_noc2_yummy),
      .data_out(buf_iob_noc2_data),           
      .valid_out(buf_iob_noc2_valid),       
      .ready_out(iob_buf_noc2_ready)    
);
valrdy_to_credit noc3_iob_to_xbar (
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(iob_buf_noc3_data),
      .valid_in(iob_buf_noc3_valid),
      .ready_in(buf_iob_noc3_ready),
      .data_out(iob_buf_xbar_noc3_data),           
      .valid_out(iob_buf_xbar_noc3_valid),       
      .yummy_out(xbar_buf_iob_noc3_yummy)    
);
credit_to_valrdy noc3_xbar_to_iob(
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(xbar_buf_iob_noc3_data),
      .valid_in(xbar_buf_iob_noc3_valid),
      .yummy_in(iob_buf_xbar_noc3_yummy),
      .data_out(buf_iob_noc3_data),           
      .valid_out(buf_iob_noc3_valid),       
      .ready_out(iob_buf_noc3_ready)    
);
valrdy_to_credit noc2_sd_to_xbar (
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(sd_buf_noc2_data),
      .valid_in(sd_buf_noc2_valid),
      .ready_in(buf_sd_noc2_ready),
      .data_out(sd_buf_xbar_noc2_data),           
      .valid_out(sd_buf_xbar_noc2_valid),       
      .yummy_out(xbar_buf_sd_noc2_yummy)    
);
credit_to_valrdy noc2_xbar_to_sd(
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(xbar_buf_sd_noc2_data),
      .valid_in(xbar_buf_sd_noc2_valid),
      .yummy_in(sd_buf_xbar_noc2_yummy),
      .data_out(buf_sd_noc2_data),           
      .valid_out(buf_sd_noc2_valid),       
      .ready_out(sd_buf_noc2_ready)    
);
valrdy_to_credit noc3_sd_to_xbar (
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(sd_buf_noc3_data),
      .valid_in(sd_buf_noc3_valid),
      .ready_in(buf_sd_noc3_ready),
      .data_out(sd_buf_xbar_noc3_data),           
      .valid_out(sd_buf_xbar_noc3_valid),       
      .yummy_out(xbar_buf_sd_noc3_yummy)    
);
credit_to_valrdy noc3_xbar_to_sd(
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(xbar_buf_sd_noc3_data),
      .valid_in(xbar_buf_sd_noc3_valid),
      .yummy_in(sd_buf_xbar_noc3_yummy),
      .data_out(buf_sd_noc3_data),           
      .valid_out(buf_sd_noc3_valid),       
      .ready_out(sd_buf_noc3_ready)    
);
valrdy_to_credit noc2_uart_to_xbar (
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(uart_buf_noc2_data),
      .valid_in(uart_buf_noc2_valid),
      .ready_in(buf_uart_noc2_ready),
      .data_out(uart_buf_xbar_noc2_data),           
      .valid_out(uart_buf_xbar_noc2_valid),       
      .yummy_out(xbar_buf_uart_noc2_yummy)    
);
credit_to_valrdy noc2_xbar_to_uart(
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(xbar_buf_uart_noc2_data),
      .valid_in(xbar_buf_uart_noc2_valid),
      .yummy_in(uart_buf_xbar_noc2_yummy),
      .data_out(buf_uart_noc2_data),           
      .valid_out(buf_uart_noc2_valid),       
      .ready_out(uart_buf_noc2_ready)    
);
valrdy_to_credit noc3_uart_to_xbar (
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(uart_buf_noc3_data),
      .valid_in(uart_buf_noc3_valid),
      .ready_in(buf_uart_noc3_ready),
      .data_out(uart_buf_xbar_noc3_data),           
      .valid_out(uart_buf_xbar_noc3_valid),       
      .yummy_out(xbar_buf_uart_noc3_yummy)    
);
credit_to_valrdy noc3_xbar_to_uart(
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(xbar_buf_uart_noc3_data),
      .valid_in(xbar_buf_uart_noc3_valid),
      .yummy_in(uart_buf_xbar_noc3_yummy),
      .data_out(buf_uart_noc3_data),           
      .valid_out(buf_uart_noc3_valid),       
      .ready_out(uart_buf_noc3_ready)    
);
valrdy_to_credit noc2_net_to_xbar (
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(net_buf_noc2_data),
      .valid_in(net_buf_noc2_valid),
      .ready_in(buf_net_noc2_ready),
      .data_out(net_buf_xbar_noc2_data),           
      .valid_out(net_buf_xbar_noc2_valid),       
      .yummy_out(xbar_buf_net_noc2_yummy)    
);
credit_to_valrdy noc2_xbar_to_net(
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(xbar_buf_net_noc2_data),
      .valid_in(xbar_buf_net_noc2_valid),
      .yummy_in(net_buf_xbar_noc2_yummy),
      .data_out(buf_net_noc2_data),           
      .valid_out(buf_net_noc2_valid),       
      .ready_out(net_buf_noc2_ready)    
);
valrdy_to_credit noc3_net_to_xbar (
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(net_buf_noc3_data),
      .valid_in(net_buf_noc3_valid),
      .ready_in(buf_net_noc3_ready),
      .data_out(net_buf_xbar_noc3_data),           
      .valid_out(net_buf_xbar_noc3_valid),       
      .yummy_out(xbar_buf_net_noc3_yummy)    
);
credit_to_valrdy noc3_xbar_to_net(
      .clk(chipset_clk),
      .reset(~chipset_rst_n),
      .data_in(xbar_buf_net_noc3_data),
      .valid_in(xbar_buf_net_noc3_valid),
      .yummy_in(net_buf_xbar_noc3_yummy),
      .data_out(buf_net_noc3_data),           
      .valid_out(buf_net_noc3_valid),       
      .ready_out(net_buf_noc3_ready)    
);
    
        f1_mc_top mc_top(
            .sys_clk(chipset_clk),
            .sys_rst_n(chipset_rst_n),
            .mc_clk(mc_clk),
            .mc_flit_in_val(buf_mem_noc2_valid),
            .mc_flit_in_data(buf_mem_noc2_data),
            .mc_flit_in_rdy(mem_buf_noc2_ready),
            .mc_flit_out_val(mem_buf_noc3_valid),
            .mc_flit_out_data(mem_buf_noc3_data),
            .mc_flit_out_rdy(buf_mem_noc3_ready),
            .uart_boot_en(uart_boot_en),
            .init_calib_complete_out(init_calib_complete),
            .mc_ui_clk_sync_rst(mc_ui_clk_sync_rst),
            
            .m_axi_awid(m_axi_awid),
            .m_axi_awaddr(m_axi_awaddr),
            .m_axi_awlen(m_axi_awlen),
            .m_axi_awsize(m_axi_awsize),
            .m_axi_awburst(m_axi_awburst),
            .m_axi_awlock(m_axi_awlock),
            .m_axi_awcache(m_axi_awcache),
            .m_axi_awprot(m_axi_awprot),
            .m_axi_awqos(m_axi_awqos),
            .m_axi_awregion(m_axi_awregion),
            .m_axi_awuser(m_axi_awuser),
            .m_axi_awvalid(m_axi_awvalid),
            .m_axi_awready(m_axi_awready),
            
            .m_axi_wid(m_axi_wid),
            .m_axi_wdata(m_axi_wdata),
            .m_axi_wstrb(m_axi_wstrb),
            .m_axi_wlast(m_axi_wlast),
            .m_axi_wuser(m_axi_wuser),
            .m_axi_wvalid(m_axi_wvalid),
            .m_axi_wready(m_axi_wready),
            
            .m_axi_arid(m_axi_arid),
            .m_axi_araddr(m_axi_araddr),
            .m_axi_arlen(m_axi_arlen),
            .m_axi_arsize(m_axi_arsize),
            .m_axi_arburst(m_axi_arburst),
            .m_axi_arlock(m_axi_arlock),
            .m_axi_arcache(m_axi_arcache),
            .m_axi_arprot(m_axi_arprot),
            .m_axi_arqos(m_axi_arqos),
            .m_axi_arregion(m_axi_arregion),
            .m_axi_aruser(m_axi_aruser),
            .m_axi_arvalid(m_axi_arvalid),
            .m_axi_arready(m_axi_arready),
            
            .m_axi_rid(m_axi_rid),
            .m_axi_rdata(m_axi_rdata),
            .m_axi_rresp(m_axi_rresp),
            .m_axi_rlast(m_axi_rlast),
            .m_axi_ruser(m_axi_ruser),
            .m_axi_rvalid(m_axi_rvalid),
            .m_axi_rready(m_axi_rready),
            
            .m_axi_bid(m_axi_bid),
            .m_axi_bresp(m_axi_bresp),
            .m_axi_buser(m_axi_buser),
            .m_axi_bvalid(m_axi_bvalid),
            .m_axi_bready(m_axi_bready), 
            .ddr_ready(ddr_ready)
        );
    
        
        
        
        
         
        
        
        
     
 
 
wire net_interrupt;
wire uart_interrupt;
wire ciop_iob_rst_n;
assign ciop_iob_rst_n = io_ctrl_rst_n & test_start & ~piton_ready_n;
ciop_iob ciop_iob     (
    .chip_clk        ( chipset_clk           ),
    .fpga_clk        ( chipset_clk           ),
    .rst_n           ( ciop_iob_rst_n        ),
    .noc1_in_val     ( intf_chipset_val_noc1 ),
    .noc1_in_data    ( intf_chipset_data_noc1),
    .noc1_in_rdy     ( intf_chipset_rdy_noc1 ),
    .noc2_out_val    ( iob_filter_noc2_valid ),
    .noc2_out_data   ( iob_filter_noc2_data  ),
    .noc2_out_rdy    ( filter_iob_noc2_ready ),
    .noc3_in_val     ( filter_iob_noc3_valid ),
    .noc3_in_data    ( filter_iob_noc3_data  ),
    .noc3_in_rdy     ( iob_filter_noc3_ready ),
    .noc2_in_val     ( buf_iob_noc2_valid    ),
    .noc2_in_data    ( buf_iob_noc2_data     ),
    .noc2_in_rdy     ( iob_buf_noc2_ready    ),
    .noc3_out_val    ( iob_buf_noc3_valid    ),
    .noc3_out_data   ( iob_buf_noc3_data     ),
    .noc3_out_rdy    ( buf_iob_noc3_ready    ),
    .uart_interrupt ( uart_interrupt         ),
    .net_interrupt  ( net_interrupt          )
);
 
 
    assign uart_interrupt = 1'b0;
    assign test_start = 1'b1;
 
    
    
    
 
 
    wire [1:0] irq_sources, irq_le;
    
    
    
     
    assign irq_le      = ext_irq[1:0];
    assign irq_sources = ext_irq_trigger[1:0];
     
    
    wire ariane_boot_sel;
  assign ariane_boot_sel   = uart_boot_en;
  
  
  
    riscv_peripherals #(
        .DataWidth      ( 64 ),
        .NumHarts       ( 1),
        .NumSources     (               2 ),
        .SwapEndianess  (               1 ),
        .DmBase         ( 64'h0000000000000000 ),
        .RomBase        ( 64'h0000000000000000 ),
        .ClintBase      ( 64'h0000000000000000 ),
        .PlicBase       ( 64'h0000000000000000 )
    ) i_riscv_peripherals (
        .clk_i                           ( chipset_clk                   ),
        .rst_ni                          ( chipset_rst_n                 ),
        .testmode_i                      ( 1'b0                          ),
        .buf_ariane_debug_noc2_data_i    ( buf_ariane_debug_noc2_data    ),
        .buf_ariane_debug_noc2_valid_i   ( buf_ariane_debug_noc2_valid   ),
        .ariane_debug_buf_noc2_ready_o   ( ariane_debug_buf_noc2_ready   ),
        .ariane_debug_buf_noc3_data_o    ( ariane_debug_buf_noc3_data    ),
        .ariane_debug_buf_noc3_valid_o   ( ariane_debug_buf_noc3_valid   ),
        .buf_ariane_debug_noc3_ready_i   ( buf_ariane_debug_noc3_ready   ),
        .buf_ariane_bootrom_noc2_data_i  ( buf_ariane_bootrom_noc2_data  ),
        .buf_ariane_bootrom_noc2_valid_i ( buf_ariane_bootrom_noc2_valid ),
        .ariane_bootrom_buf_noc2_ready_o ( ariane_bootrom_buf_noc2_ready ),
        .ariane_bootrom_buf_noc3_data_o  ( ariane_bootrom_buf_noc3_data  ),
        .ariane_bootrom_buf_noc3_valid_o ( ariane_bootrom_buf_noc3_valid ),
        .buf_ariane_bootrom_noc3_ready_i ( buf_ariane_bootrom_noc3_ready ),
        .buf_ariane_clint_noc2_data_i    ( buf_ariane_clint_noc2_data    ),
        .buf_ariane_clint_noc2_valid_i   ( buf_ariane_clint_noc2_valid   ),
        .ariane_clint_buf_noc2_ready_o   ( ariane_clint_buf_noc2_ready   ),
        .ariane_clint_buf_noc3_data_o    ( ariane_clint_buf_noc3_data    ),
        .ariane_clint_buf_noc3_valid_o   ( ariane_clint_buf_noc3_valid   ),
        .buf_ariane_clint_noc3_ready_i   ( buf_ariane_clint_noc3_ready   ),
        .buf_ariane_plic_noc2_data_i     ( buf_ariane_plic_noc2_data     ),
        .buf_ariane_plic_noc2_valid_i    ( buf_ariane_plic_noc2_valid    ),
        .ariane_plic_buf_noc2_ready_o    ( ariane_plic_buf_noc2_ready    ),
        .ariane_plic_buf_noc3_data_o     ( ariane_plic_buf_noc3_data     ),
        .ariane_plic_buf_noc3_valid_o    ( ariane_plic_buf_noc3_valid    ),
        .buf_ariane_plic_noc3_ready_i    ( buf_ariane_plic_noc3_ready    ),
        
        .ariane_boot_sel_i               ( ariane_boot_sel               ),
        
        .ndmreset_o                      ( ndmreset_o                    ),
        .dmactive_o                      ( dmactive_o                    ),
        .debug_req_o                     ( debug_req_o                   ),
        .unavailable_i                   ( unavailable_i                 ),
        
        .tck_i                           ( tck_i                         ),
        .tms_i                           ( tms_i                         ),
        .trst_ni                         ( trst_ni                       ),
        .td_i                            ( td_i                          ),
        .td_o                            ( td_o                          ),
        .tdo_oe_o                        (                               ),
        
        .rtc_i                           ( rtc_i                         ),
        .timer_irq_o                     ( timer_irq_o                   ),
        .ipi_o                           ( ipi_o                         ),
        
        .irq_le_i                        ( irq_le                        ), 
        .irq_sources_i                   ( irq_sources                   ),
        .irq_o                           ( irq_o                         )
    );
endmodule
module packet_filter (
    input wire clk,
    input wire rst_n,
    
    input wire                          noc2_filter_val,
    input wire [64 - 1:0]  noc2_filter_data,
    output reg                         filter_noc2_rdy,
    
    output wire                         filter_noc3_val,
    output wire [64 - 1:0] filter_noc3_data,
    input wire                          noc3_filter_rdy,
    
    output reg                         filter_xbar_val,
    output reg [64 - 1:0] filter_xbar_data,
    input wire                          xbar_filter_rdy,
    
    input wire                          xbar_filter_val,
    input wire  [64 - 1:0] xbar_filter_data,
    output wire                         filter_xbar_rdy,
    
    input wire                          uart_boot_en,
    
    output wire                         invalid_access_o
);
    localparam IDLE = 3'b000;
    localparam ONLYHEADERFLIT = 3'b001;
    localparam ONEFLIT = 3'b010;
    localparam TWOFLITS = 3'b011;
    localparam SENDING = 3'b100;
    localparam DRAINTWO = 3'b101;
    localparam DRAINONE = 3'b110;
    reg [64-1:0] flit_buffer_0_reg;
    reg [64-1:0] flit_buffer_1_reg;
    reg [64-1:0] flit_buffer_0_next;
    reg [64-1:0] flit_buffer_1_next;
    reg [64-1:0] readdressed_flit0;
    reg [8-1:0] num_flits_reg; 
    reg [8-1:0] num_flits_next; 
    reg [8-1:0] flits_sent_reg; 
    reg [8-1:0] flits_sent_next; 
    reg [2:0] state_reg;
    reg [2:0] state_next;
    reg invalid_access, invalid_access_d, invalid_access_q;
    always @* begin
		    invalid_access_d = invalid_access_q;
        case (state_reg)
        IDLE: begin
            filter_xbar_val = 1'b0;
            filter_xbar_data = 64'b0;
            filter_noc2_rdy = 1'b1;
            flit_buffer_0_next = noc2_filter_val ? noc2_filter_data : 64'b0;
            flit_buffer_1_next = 64'b0;
            num_flits_next = noc2_filter_val ? noc2_filter_data[29:22] : 8'b0;
            flits_sent_next = 8'b0;
            
            if (noc2_filter_val & (noc2_filter_data[29:22] == 8'b0)) begin
                filter_xbar_val = 1'b1;
                filter_xbar_data = flit_buffer_0_reg;
                state_next = xbar_filter_rdy ? IDLE : ONLYHEADERFLIT;
            end
            else begin
                state_next = noc2_filter_val ? ONEFLIT : IDLE;
            end
        end
        ONLYHEADERFLIT: begin
            if (xbar_filter_rdy) begin
                
                filter_xbar_val = 1'b1;
                filter_xbar_data = flit_buffer_0_reg;
                filter_noc2_rdy = 1'b1;
                flit_buffer_0_next = noc2_filter_val ? noc2_filter_data : 64'b0;
                flit_buffer_1_next = 64'b0;
                num_flits_next = noc2_filter_val ? noc2_filter_data[29:22] : 8'b0;
                flits_sent_next = 8'b0;
                
                if (noc2_filter_val & (noc2_filter_data[29:22] == 8'b0)) begin
                    filter_xbar_val = 1'b1;
                    filter_xbar_data = flit_buffer_0_reg;
                    state_next = xbar_filter_rdy ? IDLE : ONLYHEADERFLIT;
                end
                else begin
                    state_next = noc2_filter_val ? ONEFLIT : IDLE;
                end
            end else begin
                
                filter_xbar_val = 1'b1;
                filter_xbar_data = flit_buffer_0_reg;
                filter_noc2_rdy = 1'b0;
                flit_buffer_0_next = flit_buffer_0_reg;
                flit_buffer_1_next = 64'b0;
                num_flits_next = num_flits_reg;
                flits_sent_next = 8'b0;
                state_next = ONLYHEADERFLIT;
            end
        end
        ONEFLIT: begin
            filter_xbar_val = 1'b0;
            filter_xbar_data = 64'b0;
            filter_noc2_rdy = 1'b1;
            flit_buffer_0_next = noc2_filter_val ? readdressed_flit0 : flit_buffer_0_reg;
            flit_buffer_1_next = noc2_filter_val ? noc2_filter_data : 64'b0;
            num_flits_next = num_flits_reg;
            flits_sent_next = 8'b0;
            state_next = noc2_filter_val ? TWOFLITS : ONEFLIT;
		        invalid_access_d = invalid_access_q | (noc2_filter_val & invalid_access);
		end
        TWOFLITS: begin
            if ((num_flits_reg == 8'd1)) begin
                if (xbar_filter_rdy) begin
                    filter_xbar_val = 1'b1;
                    filter_xbar_data = flit_buffer_0_reg;
                    filter_noc2_rdy = 1'b0;
                    flit_buffer_0_next = flit_buffer_1_reg;
                    flit_buffer_1_next = noc2_filter_data;
                    num_flits_next = num_flits_reg;
                    flits_sent_next = 8'b1;
                    state_next = DRAINONE;
                end
                else begin
                    filter_xbar_val = 1'b1;
                    filter_xbar_data = flit_buffer_0_reg;
                    filter_noc2_rdy = 1'b0;
                    flit_buffer_0_next = flit_buffer_0_reg;
                    flit_buffer_1_next = flit_buffer_1_reg;
                    num_flits_next = num_flits_reg;
                    flits_sent_next = 8'b0;
                    state_next = TWOFLITS;
                end
            end
            else if (xbar_filter_rdy & noc2_filter_val) begin
                filter_xbar_val = 1'b1;
                filter_xbar_data = flit_buffer_0_reg;
                filter_noc2_rdy = 1'b1;
                flit_buffer_0_next = flit_buffer_1_reg;
                flit_buffer_1_next = noc2_filter_data;
                num_flits_next = num_flits_reg;
                flits_sent_next = 8'b1;
                state_next = (num_flits_reg == 8'd2) ? DRAINTWO : SENDING;
            end
            else begin
                filter_xbar_val = 1'b0;
                filter_xbar_data = flit_buffer_0_reg;
                filter_noc2_rdy = 1'b0;
                flit_buffer_0_next = flit_buffer_0_reg;
                flit_buffer_1_next = flit_buffer_1_reg;
                num_flits_next = num_flits_reg;
                flits_sent_next = 8'b0;
                state_next = TWOFLITS;
            end
        end
        SENDING: begin
            if (xbar_filter_rdy & noc2_filter_val & (flits_sent_reg < (num_flits_reg + 1'b1))) begin
                filter_xbar_val = 1'b1;
                filter_xbar_data = flit_buffer_0_reg;
                filter_noc2_rdy = 1'b1;
                flit_buffer_0_next = flit_buffer_1_reg;
                flit_buffer_1_next = noc2_filter_data;
                num_flits_next = num_flits_reg;
                flits_sent_next = flits_sent_reg + 1'b1; 
                
                state_next = (flits_sent_reg == (num_flits_reg - 2'd2)) ? DRAINTWO : SENDING;
            end else begin
                filter_xbar_val = 1'b0;
                filter_xbar_data = flit_buffer_0_reg;
                filter_noc2_rdy = 1'b0;
                flit_buffer_0_next = flit_buffer_0_reg;
                flit_buffer_1_next = flit_buffer_1_reg;
                num_flits_next = num_flits_reg;
                flits_sent_next = flits_sent_reg;
                state_next = SENDING;
            end
        end
        DRAINTWO: begin
            if (xbar_filter_rdy) begin
                filter_xbar_val = 1'b1;
                filter_xbar_data = flit_buffer_0_reg;
                filter_noc2_rdy = 1'b0;
                flit_buffer_0_next = flit_buffer_1_reg;
                flit_buffer_1_next = 64'b0;
                num_flits_next = num_flits_reg;
                flits_sent_next = flits_sent_reg + 1'b1; 
                state_next = DRAINONE;
            end else begin
                filter_xbar_val = 1'b0;
                filter_xbar_data = flit_buffer_0_reg;
                filter_noc2_rdy = 1'b0;
                flit_buffer_0_next = flit_buffer_0_reg;
                flit_buffer_1_next = flit_buffer_1_reg;
                num_flits_next = num_flits_reg;
                flits_sent_next = flits_sent_reg;
                state_next = DRAINTWO;
            end
        end
        DRAINONE: begin
            if (xbar_filter_rdy) begin
                filter_xbar_val = 1'b1;
                filter_xbar_data = flit_buffer_0_reg;
                filter_noc2_rdy = 1'b0;
                flit_buffer_0_next = 64'b0;
                flit_buffer_1_next = 64'b0;
                num_flits_next = 8'b0;
                flits_sent_next = 8'b0; 
                state_next = IDLE;
            end else begin
                filter_xbar_val = 1'b0;
                filter_xbar_data = flit_buffer_0_reg;
                filter_noc2_rdy = 1'b0;
                flit_buffer_0_next = flit_buffer_0_reg;
                flit_buffer_1_next = flit_buffer_1_reg;
                num_flits_next = num_flits_reg;
                flits_sent_next = flits_sent_reg;
                state_next = DRAINONE;
            end
        end
        default: begin
            filter_xbar_val = 1'bX;
            filter_xbar_data = 64'bX;
            filter_noc2_rdy = 1'bX;
            flit_buffer_0_next = 64'bX;
            flit_buffer_1_next = 64'bX;
            num_flits_next = 8'bX;
            flits_sent_next = 8'bX;
            state_next = 3'bX;
        end
        endcase
    end
    always @* begin
        readdressed_flit0 = flit_buffer_0_reg;
        invalid_access  = 1'b0;
        if (flit_buffer_0_reg[21:14] == 8'd19 ||
            flit_buffer_0_reg[21:14] == 8'd20 ||
            flit_buffer_0_reg[21:14] == 8'd14 ||
            flit_buffer_0_reg[21:14] == 8'd15) begin
                if ((noc2_filter_data[((16 + 40 - 1)):(16)] >= 40'h9f00000000 && noc2_filter_data[((16 + 40 - 1)):(16)] < 40'h9f00000000 + 40'h10) & (~uart_boot_en))
                begin
                    readdressed_flit0[49:42] = 8'h2;
                end
                else if ((noc2_filter_data[((16 + 40 - 1)):(16)] >= 40'hf000000000 && noc2_filter_data[((16 + 40 - 1)):(16)] < 40'hf000000000 + 40'hff0300000) & (~uart_boot_en))
                begin
                    readdressed_flit0[49:42] = 8'h3;
                end
                else if ((noc2_filter_data[((16 + 40 - 1)):(16)] >= 40'hfff0c2c000 && noc2_filter_data[((16 + 40 - 1)):(16)] < 40'hfff0c2c000 + 40'hd4000))
                begin
                    readdressed_flit0[49:42] = 8'h4;
                end
                else if ((noc2_filter_data[((16 + 40 - 1)):(16)] >= 40'hfff0d00000 && noc2_filter_data[((16 + 40 - 1)):(16)] < 40'hfff0d00000 + 40'h100000) & (~uart_boot_en))
                begin
                    readdressed_flit0[49:42] = 8'h5;
                end
                else begin
 
                  
                  readdressed_flit0[49:42] = 8'h1;
 
                end
        end
    end
    assign invalid_access_o = invalid_access_q;
    always @(posedge clk) begin
        if (!rst_n) begin
            invalid_access_q  <= 1'b0;
            flit_buffer_0_reg <= 64'd0;
            flit_buffer_1_reg <= 64'd0;
            num_flits_reg     <= 8'd0;
            flits_sent_reg    <= 8'd0;
            state_reg         <= IDLE;
        end
        else
        begin
      			invalid_access_q  <= invalid_access_d;
			      flit_buffer_0_reg <= flit_buffer_0_next;
            flit_buffer_1_reg <= flit_buffer_1_next;
            num_flits_reg     <= num_flits_next;
            flits_sent_reg    <= flits_sent_next;
            state_reg         <= state_next;
        end
    end
    
    
    
    assign filter_xbar_rdy = noc3_filter_rdy;
    assign filter_noc3_val = xbar_filter_val;
    assign filter_noc3_data = xbar_filter_data;
endmodule
module storage_addr_trans #(parameter MEM_ADDR_WIDTH=64, VA_ADDR_WIDTH=40, STORAGE_ADDR_WIDTH=12)
(
    input       [VA_ADDR_WIDTH-1:0]         va_byte_addr,
    output      [STORAGE_ADDR_WIDTH-1:0]    storage_addr_out,
    output                                  hit_any_section
);
wire [63:0] storage_addr;
wire [63:0]                      bram_addr_0;
wire                          in_section_0;
assign storage_addr = ({STORAGE_ADDR_WIDTH{in_section_0}} & bram_addr_0[STORAGE_ADDR_WIDTH-1:0]);
assign storage_addr_out = {storage_addr, 3'b0};
assign hit_any_section = in_section_0 ;
endmodule
module storage_addr_trans_unified #(parameter MEM_ADDR_WIDTH=64, VA_ADDR_WIDTH=40, STORAGE_ADDR_WIDTH=12)
(
    input       [VA_ADDR_WIDTH-1:0]         va_byte_addr,
    output      [STORAGE_ADDR_WIDTH-1:0]    storage_addr_out,
    output                                  hit_any_section
);
wire [63:0] storage_addr;
wire [63:0]                      bram_addr_0;
wire                          in_section_0;
assign storage_addr = ({STORAGE_ADDR_WIDTH{in_section_0}} & bram_addr_0[STORAGE_ADDR_WIDTH-1:0]);
assign storage_addr_out = {storage_addr, 3'b0};
assign hit_any_section = in_section_0 ;
endmodule
module dynamic_node_top_wrap
(
    input clk,
    input reset_in,
       
    input [64-1:0] dataIn_N,   
    input [64-1:0] dataIn_E,
    input [64-1:0] dataIn_S,
    input [64-1:0] dataIn_W,
     input [64-1:0] dataIn_P,   
       
    input validIn_N,        
    input validIn_E,
    input validIn_S,
    input validIn_W,
    input validIn_P,        
       
    input yummyIn_N,        
    input yummyIn_E,
    input yummyIn_S,
    input yummyIn_W,
    input yummyIn_P,        
       
    input [8-1:0] myLocX,       
    input [8-1:0] myLocY,
    input [14-1:0] myChipID,
    output [64-1:0] dataOut_N, 
    output [64-1:0] dataOut_E,
    output [64-1:0] dataOut_S,
     output [64-1:0] dataOut_W,
     output [64-1:0] dataOut_P, 
    
    output validOut_N,      
    output validOut_E,
    output validOut_S,
    output validOut_W,
    output validOut_P,      
       
    output yummyOut_N,      
    output yummyOut_E,
    output yummyOut_S,
    output yummyOut_W,
    output yummyOut_P,      
    
    
    output thanksIn_P      
);
    dynamic_node_top dynamic_node_top
    (
        .clk(clk),
        .reset_in(reset_in),
        .dataIn_N(dataIn_N),
        .dataIn_E(dataIn_E),
        .dataIn_S(dataIn_S),
        .dataIn_W(dataIn_W),
        .dataIn_P(dataIn_P),
        .validIn_N(validIn_N),
        .validIn_E(validIn_E),
        .validIn_S(validIn_S),
        .validIn_W(validIn_W),
        .validIn_P(validIn_P),
        .yummyIn_N(yummyIn_N),
        .yummyIn_E(yummyIn_E),
        .yummyIn_S(yummyIn_S),
        .yummyIn_W(yummyIn_W),
        .yummyIn_P(yummyIn_P),
        .myLocX(myLocX),
        .myLocY(myLocY),
        .myChipID(myChipID),
        .ec_cfg(15'b0),
        .store_meter_partner_address_X(5'b0),
        .store_meter_partner_address_Y(5'b0),
        .dataOut_N(dataOut_N),
        .dataOut_E(dataOut_E),
        .dataOut_S(dataOut_S),
        .dataOut_W(dataOut_W),
        .dataOut_P(dataOut_P),
        .validOut_N(validOut_N),
        .validOut_E(validOut_E),
        .validOut_S(validOut_S),
        .validOut_W(validOut_W),
        .validOut_P(validOut_P),
        .yummyOut_N(yummyOut_N),
        .yummyOut_E(yummyOut_E),
        .yummyOut_W(yummyOut_W),
        .yummyOut_S(yummyOut_S),
        .yummyOut_P(yummyOut_P),
        .thanksIn_P(thanksIn_P),
        .external_interrupt(),
        .store_meter_ack_partner(),
        .store_meter_ack_non_partner(),
        .ec_out()
    ); 
endmodule
module dynamic_node_top(clk,
		    reset_in,
		    dataIn_N,
		    dataIn_E,
		    dataIn_S,
		    dataIn_W,
		    dataIn_P,
		    validIn_N,
		    validIn_E,
		    validIn_S,
		    validIn_W,
		    validIn_P,
		    yummyIn_N,
		    yummyIn_E,
		    yummyIn_S,
		    yummyIn_W,
		    yummyIn_P,
		    myLocX,
		    myLocY,
            myChipID,
		    store_meter_partner_address_X,
		    store_meter_partner_address_Y,
		    ec_cfg,
		    dataOut_N,
		    dataOut_E,
		    dataOut_S,
		    dataOut_W,
		    dataOut_P,
		    validOut_N,
		    validOut_E,
		    validOut_S,
		    validOut_W,
		    validOut_P,
		    yummyOut_N,
		    yummyOut_E,
		    yummyOut_S,
		    yummyOut_W,
		    yummyOut_P,
		    thanksIn_P,
		    external_interrupt,
		    store_meter_ack_partner,
		    store_meter_ack_non_partner,
		    ec_out);
input clk;
input reset_in;
   
input [64-1:0] dataIn_N;	
input [64-1:0] dataIn_E;
input [64-1:0] dataIn_S;
input [64-1:0] dataIn_W;
input [64-1:0] dataIn_P;	
   
input validIn_N;		
input validIn_E;
input validIn_S;
input validIn_W;
input validIn_P;		
   
input yummyIn_N;		
input yummyIn_E;
input yummyIn_S;
input yummyIn_W;
input yummyIn_P;		
   
input [8-1:0] myLocX;		
input [8-1:0] myLocY;
input [14-1:0] myChipID;
input [4:0] store_meter_partner_address_X;
input [4:0] store_meter_partner_address_Y;
input [14:0] ec_cfg;            
output [64-1:0] dataOut_N;	
output [64-1:0] dataOut_E;
output [64-1:0] dataOut_S;
output [64-1:0] dataOut_W;
output [64-1:0] dataOut_P;	
output validOut_N;		
output validOut_E;
output validOut_S;
output validOut_W;
output validOut_P;		
   
output yummyOut_N;		
output yummyOut_E;
output yummyOut_S;
output yummyOut_W;
output yummyOut_P;		
output thanksIn_P;		
output external_interrupt;	
				
output store_meter_ack_partner;      
                                     
output store_meter_ack_non_partner;  
                                     
output [4:0] ec_out;
wire   ec_wants_to_send_but_cannot_N,
       ec_wants_to_send_but_cannot_E,
       ec_wants_to_send_but_cannot_S,
       ec_wants_to_send_but_cannot_W,
       ec_wants_to_send_but_cannot_P;
   wire store_ack_received;
   wire store_ack_received_r;
   wire [9:0] store_ack_addr;
   wire [9:0] store_ack_addr_r;
wire north_input_tail;
wire east_input_tail;
wire south_input_tail;
wire west_input_tail;
wire proc_input_tail;
wire [64-1:0] north_input_data;
wire [64-1:0] east_input_data;
wire [64-1:0] south_input_data;
wire [64-1:0] west_input_data;
wire [64-1:0] proc_input_data;
wire north_input_valid;
wire east_input_valid;
wire south_input_valid;
wire west_input_valid;
wire proc_input_valid;
wire thanks_n_to_n;
wire thanks_n_to_e;
wire thanks_n_to_s;
wire thanks_n_to_w;
wire thanks_n_to_p;
wire thanks_e_to_n;
wire thanks_e_to_e;
wire thanks_e_to_s;
wire thanks_e_to_w;
wire thanks_e_to_p;
wire thanks_s_to_n;
wire thanks_s_to_e;
wire thanks_s_to_s;
wire thanks_s_to_w;
wire thanks_s_to_p;
wire thanks_w_to_n;
wire thanks_w_to_e;
wire thanks_w_to_s;
wire thanks_w_to_w;
wire thanks_w_to_p;
wire thanks_p_to_n;
wire thanks_p_to_e;
wire thanks_p_to_s;
wire thanks_p_to_w;
wire thanks_p_to_p;
wire route_req_n_to_n;
wire route_req_n_to_e;
wire route_req_n_to_s;
wire route_req_n_to_w;
wire route_req_n_to_p;
wire route_req_e_to_n;
wire route_req_e_to_e;
wire route_req_e_to_s;
wire route_req_e_to_w;
wire route_req_e_to_p;
wire route_req_s_to_n;
wire route_req_s_to_e;
wire route_req_s_to_s;
wire route_req_s_to_w;
wire route_req_s_to_p;
wire route_req_w_to_n;
wire route_req_w_to_e;
wire route_req_w_to_s;
wire route_req_w_to_w;
wire route_req_w_to_p;
wire route_req_p_to_n;
wire route_req_p_to_e;
wire route_req_p_to_s;
wire route_req_p_to_w;
wire route_req_p_to_p;
wire default_ready_n_to_s;
wire default_ready_e_to_w;
wire default_ready_s_to_n;
wire default_ready_s_to_p;
wire default_ready_w_to_e;
wire yummyOut_N_internal;
wire yummyOut_E_internal;
wire yummyOut_S_internal;
wire yummyOut_W_internal;
wire yummyOut_P_internal;
wire validOut_N_internal;
wire validOut_E_internal;
wire validOut_S_internal;
wire validOut_W_internal;
wire validOut_P_internal;
wire [64-1:0] dataOut_N_internal;
wire [64-1:0] dataOut_E_internal;
wire [64-1:0] dataOut_S_internal;
wire [64-1:0] dataOut_W_internal;
wire [64-1:0] dataOut_P_internal;
wire yummyOut_N_flip1_out;
wire yummyOut_E_flip1_out;
wire yummyOut_S_flip1_out;
wire yummyOut_W_flip1_out;
wire validOut_N_flip1_out;
wire validOut_E_flip1_out;
wire validOut_S_flip1_out;
wire validOut_W_flip1_out;
wire [64-1:0] dataOut_N_flip1_out;
wire [64-1:0] dataOut_E_flip1_out;
wire [64-1:0] dataOut_S_flip1_out;
wire [64-1:0] dataOut_W_flip1_out;
wire yummyIn_N_internal;
wire yummyIn_E_internal;
wire yummyIn_S_internal;
wire yummyIn_W_internal;
wire yummyIn_P_internal;
wire validIn_N_internal;
wire validIn_E_internal;
wire validIn_S_internal;
wire validIn_W_internal;
wire [64-1:0] dataIn_N_internal;
wire [64-1:0] dataIn_E_internal;
wire [64-1:0] dataIn_S_internal;
wire [64-1:0] dataIn_W_internal;
wire yummyIn_N_flip1_out;
wire yummyIn_E_flip1_out;
wire yummyIn_S_flip1_out;
wire yummyIn_W_flip1_out;
wire validIn_N_flip1_out;
wire validIn_E_flip1_out;
wire validIn_S_flip1_out;
wire validIn_W_flip1_out;
wire [64-1:0] dataIn_N_flip1_out;
wire [64-1:0] dataIn_E_flip1_out;
wire [64-1:0] dataIn_S_flip1_out;
wire [64-1:0] dataIn_W_flip1_out;
reg [8-1:0] myLocX_f;
reg [8-1:0] myLocY_f;
reg [14-1:0] myChipID_f;
wire   reset;
reg ec_thanks_n_to_n_reg, ec_thanks_n_to_e_reg, ec_thanks_n_to_s_reg, ec_thanks_n_to_w_reg, ec_thanks_n_to_p_reg;
reg ec_thanks_e_to_n_reg, ec_thanks_e_to_e_reg, ec_thanks_e_to_s_reg, ec_thanks_e_to_w_reg, ec_thanks_e_to_p_reg;
reg ec_thanks_s_to_n_reg, ec_thanks_s_to_e_reg, ec_thanks_s_to_s_reg, ec_thanks_s_to_w_reg, ec_thanks_s_to_p_reg;
reg ec_thanks_w_to_n_reg, ec_thanks_w_to_e_reg, ec_thanks_w_to_s_reg, ec_thanks_w_to_w_reg, ec_thanks_w_to_p_reg;
reg ec_thanks_p_to_n_reg, ec_thanks_p_to_e_reg, ec_thanks_p_to_s_reg, ec_thanks_p_to_w_reg, ec_thanks_p_to_p_reg;
reg ec_wants_to_send_but_cannot_N_reg, ec_wants_to_send_but_cannot_E_reg, ec_wants_to_send_but_cannot_S_reg, ec_wants_to_send_but_cannot_W_reg, ec_wants_to_send_but_cannot_P_reg;
reg ec_north_input_valid_reg, ec_east_input_valid_reg, ec_south_input_valid_reg, ec_west_input_valid_reg, ec_proc_input_valid_reg;
always @(posedge clk)
  begin
     ec_thanks_n_to_n_reg <= thanks_n_to_n; ec_thanks_n_to_e_reg <= thanks_n_to_e; ec_thanks_n_to_s_reg <= thanks_n_to_s; ec_thanks_n_to_w_reg <= thanks_n_to_w; ec_thanks_n_to_p_reg <= thanks_n_to_p;
     ec_thanks_e_to_n_reg <= thanks_e_to_n; ec_thanks_e_to_e_reg <= thanks_e_to_e; ec_thanks_e_to_s_reg <= thanks_e_to_s; ec_thanks_e_to_w_reg <= thanks_e_to_w; ec_thanks_e_to_p_reg <= thanks_e_to_p;
     ec_thanks_s_to_n_reg <= thanks_s_to_n; ec_thanks_s_to_e_reg <= thanks_s_to_e; ec_thanks_s_to_s_reg <= thanks_s_to_s; ec_thanks_s_to_w_reg <= thanks_s_to_w; ec_thanks_s_to_p_reg <= thanks_s_to_p;
     ec_thanks_w_to_n_reg <= thanks_w_to_n; ec_thanks_w_to_e_reg <= thanks_w_to_e; ec_thanks_w_to_s_reg <= thanks_w_to_s; ec_thanks_w_to_w_reg <= thanks_w_to_w; ec_thanks_w_to_p_reg <= thanks_w_to_p;
     ec_thanks_p_to_n_reg <= thanks_p_to_n; ec_thanks_p_to_e_reg <= thanks_p_to_e; ec_thanks_p_to_s_reg <= thanks_p_to_s; ec_thanks_p_to_w_reg <= thanks_p_to_w; ec_thanks_p_to_p_reg <= thanks_p_to_p;
     ec_wants_to_send_but_cannot_N_reg <= ec_wants_to_send_but_cannot_N;
     ec_wants_to_send_but_cannot_E_reg <= ec_wants_to_send_but_cannot_E;
     ec_wants_to_send_but_cannot_S_reg <= ec_wants_to_send_but_cannot_S;
     ec_wants_to_send_but_cannot_W_reg <= ec_wants_to_send_but_cannot_W;
     ec_wants_to_send_but_cannot_P_reg <= ec_wants_to_send_but_cannot_P;
     ec_north_input_valid_reg <= north_input_valid;
     ec_east_input_valid_reg  <= east_input_valid;
     ec_south_input_valid_reg <= south_input_valid;
     ec_west_input_valid_reg  <= west_input_valid;
     ec_proc_input_valid_reg  <= proc_input_valid;
  end
   wire ec_thanks_to_n = ec_thanks_n_to_n_reg | ec_thanks_e_to_n_reg | ec_thanks_s_to_n_reg | ec_thanks_w_to_n_reg | ec_thanks_p_to_n_reg;
   wire ec_thanks_to_e = ec_thanks_n_to_e_reg | ec_thanks_e_to_e_reg | ec_thanks_s_to_e_reg | ec_thanks_w_to_e_reg | ec_thanks_p_to_e_reg;
   wire ec_thanks_to_s = ec_thanks_n_to_s_reg | ec_thanks_e_to_s_reg | ec_thanks_s_to_s_reg | ec_thanks_w_to_s_reg | ec_thanks_p_to_s_reg;
   wire ec_thanks_to_w = ec_thanks_n_to_w_reg | ec_thanks_e_to_w_reg | ec_thanks_s_to_w_reg | ec_thanks_w_to_w_reg | ec_thanks_p_to_w_reg;
   wire ec_thanks_to_p = ec_thanks_n_to_p_reg | ec_thanks_e_to_p_reg | ec_thanks_s_to_p_reg | ec_thanks_w_to_p_reg | ec_thanks_p_to_p_reg;
one_of_eight #(1) ec_mux_north(.in0(ec_wants_to_send_but_cannot_N),
                        .in1(ec_thanks_p_to_n_reg),
                        .in2(ec_thanks_w_to_n_reg),
                        .in3(ec_thanks_s_to_n_reg),
                        .in4(ec_thanks_e_to_n_reg),
                        .in5(ec_thanks_n_to_n_reg),
                        .in6(ec_thanks_to_n),
                        .in7(ec_north_input_valid_reg & ~ec_thanks_to_n),
                        .sel(ec_cfg[14:12]),
                        .out(ec_out[4]));
one_of_eight #(1) ec_mux_east(.in0(ec_wants_to_send_but_cannot_E),
                       .in1(ec_thanks_p_to_e_reg),
                       .in2(ec_thanks_w_to_e_reg),
                       .in3(ec_thanks_s_to_e_reg),
                       .in4(ec_thanks_e_to_e_reg),
                       .in5(ec_thanks_n_to_e_reg),
                       .in6(ec_thanks_to_e),
                       .in7(ec_east_input_valid_reg & ~ec_thanks_to_e),
                       .sel(ec_cfg[11:9]),
                       .out(ec_out[3]));
one_of_eight #(1) ec_mux_south(.in0(ec_wants_to_send_but_cannot_S),
                        .in1(ec_thanks_p_to_s_reg),
                        .in2(ec_thanks_w_to_s_reg),
                        .in3(ec_thanks_s_to_s_reg),
                        .in4(ec_thanks_e_to_s_reg),
                        .in5(ec_thanks_n_to_s_reg),
                        .in6(ec_thanks_to_s),
                        .in7(ec_south_input_valid_reg & ~ec_thanks_to_s),
                        .sel(ec_cfg[8:6]),
                        .out(ec_out[2]));
one_of_eight #(1) ec_mux_west( .in0(ec_wants_to_send_but_cannot_W),
                        .in1(ec_thanks_p_to_w_reg),
                        .in2(ec_thanks_w_to_w_reg),
                        .in3(ec_thanks_s_to_w_reg),
                        .in4(ec_thanks_e_to_w_reg),
                        .in5(ec_thanks_n_to_w_reg),
                        .in6(ec_thanks_to_w),
                        .in7(ec_west_input_valid_reg & ~ec_thanks_to_w),
                        .sel(ec_cfg[5:3]),
                        .out(ec_out[1]));
one_of_eight #(1) ec_mux_proc( .in0(ec_wants_to_send_but_cannot_P),
                        .in1(ec_thanks_p_to_p_reg),
                        .in2(ec_thanks_w_to_p_reg),
                        .in3(ec_thanks_s_to_p_reg),
                        .in4(ec_thanks_e_to_p_reg),
                        .in5(ec_thanks_n_to_p_reg),
                        .in6(ec_thanks_to_p),
                        .in7(ec_proc_input_valid_reg & ~ec_thanks_to_p),
                        .sel(ec_cfg[2:0]),
                        .out(ec_out[0]));
net_dff #(1) REG_reset_fin(.d(reset_in), .q(reset), .clk(clk));
net_dff #(10) REG_store_ack_addr(   .d(store_ack_addr),     .q(store_ack_addr_r),     .clk(clk));
net_dff #(1) REG_store_ack_received(.d(store_ack_received), .q(store_ack_received_r), .clk(clk));
   wire is_partner_address_v_r;
   bus_compare_equal #(10) CMP_partner_address (.a(store_ack_addr_r),
                                        .b({ store_meter_partner_address_Y, store_meter_partner_address_X } ),
                                        .bus_equal(is_partner_address_v_r));
   assign store_meter_ack_partner     = is_partner_address_v_r & store_ack_received_r;
   assign store_meter_ack_non_partner = ~is_partner_address_v_r & store_ack_received_r;
always @ (posedge clk)
begin
        if(reset)
        begin
                myLocY_f <= 8'd0;
                myLocX_f <= 8'd0;
                myChipID_f <= 14'd0;
        end
        else
        begin
                myLocY_f <= myLocY;
                myLocX_f <= myLocX;
                myChipID_f <= myChipID;
        end
end
assign thanksIn_P = thanks_n_to_p | thanks_e_to_p | thanks_s_to_p | thanks_w_to_p | thanks_p_to_p;
assign validOut_P = validOut_P_internal;
assign dataOut_P = dataOut_P_internal;
assign yummyIn_P_internal = yummyIn_P;
assign yummyOut_P = yummyOut_P_internal;
   
flip_bus #(1, 14) yummyOut_N_flip1(yummyOut_N_internal, yummyOut_N_flip1_out);
flip_bus #(1, 14) yummyOut_E_flip1(yummyOut_E_internal, yummyOut_E_flip1_out);
flip_bus #(1, 14) yummyOut_S_flip1(yummyOut_S_internal, yummyOut_S_flip1_out);
flip_bus #(1, 14) yummyOut_W_flip1(yummyOut_W_internal, yummyOut_W_flip1_out);
flip_bus #(1, 21) yummyOut_N_flip2(yummyOut_N_flip1_out, yummyOut_N);
flip_bus #(1, 21) yummyOut_E_flip2(yummyOut_E_flip1_out, yummyOut_E);
flip_bus #(1, 21) yummyOut_S_flip2(yummyOut_S_flip1_out, yummyOut_S);
flip_bus #(1, 21) yummyOut_W_flip2(yummyOut_W_flip1_out, yummyOut_W);
flip_bus #(1, 14) validOut_N_flip1(validOut_N_internal, validOut_N_flip1_out);
flip_bus #(1, 14) validOut_E_flip1(validOut_E_internal, validOut_E_flip1_out);
flip_bus #(1, 14) validOut_S_flip1(validOut_S_internal, validOut_S_flip1_out);
flip_bus #(1, 14) validOut_W_flip1(validOut_W_internal, validOut_W_flip1_out);
flip_bus #(1, 21) validOut_N_flip2(validOut_N_flip1_out, validOut_N);
flip_bus #(1, 21) validOut_E_flip2(validOut_E_flip1_out, validOut_E);
flip_bus #(1, 21) validOut_S_flip2(validOut_S_flip1_out, validOut_S);
flip_bus #(1, 21) validOut_W_flip2(validOut_W_flip1_out, validOut_W);
flip_bus #(64, 14) dataOut_N_flip1(dataOut_N_internal, dataOut_N_flip1_out);
flip_bus #(64, 14) dataOut_E_flip1(dataOut_E_internal, dataOut_E_flip1_out);
flip_bus #(64, 14) dataOut_S_flip1(dataOut_S_internal, dataOut_S_flip1_out);
flip_bus #(64, 14) dataOut_W_flip1(dataOut_W_internal, dataOut_W_flip1_out);
flip_bus #(64, 21) dataOut_N_flip2(dataOut_N_flip1_out, dataOut_N);
flip_bus #(64, 21) dataOut_E_flip2(dataOut_E_flip1_out, dataOut_E);
flip_bus #(64, 21) dataOut_S_flip2(dataOut_S_flip1_out, dataOut_S);
flip_bus #(64, 21) dataOut_W_flip2(dataOut_W_flip1_out, dataOut_W);
flip_bus #(1, 14) yummyIn_N_flip1(yummyIn_N, yummyIn_N_flip1_out);
flip_bus #(1, 14) yummyIn_E_flip1(yummyIn_E, yummyIn_E_flip1_out);
flip_bus #(1, 14) yummyIn_S_flip1(yummyIn_S, yummyIn_S_flip1_out);
flip_bus #(1, 14) yummyIn_W_flip1(yummyIn_W, yummyIn_W_flip1_out);
flip_bus #(1, 10) yummyIn_N_flip2(yummyIn_N_flip1_out, yummyIn_N_internal);
flip_bus #(1, 10) yummyIn_E_flip2(yummyIn_E_flip1_out, yummyIn_E_internal);
flip_bus #(1, 10) yummyIn_S_flip2(yummyIn_S_flip1_out, yummyIn_S_internal);
flip_bus #(1, 10) yummyIn_W_flip2(yummyIn_W_flip1_out, yummyIn_W_internal);
flip_bus #(1, 14) validIn_N_flip1(validIn_N, validIn_N_flip1_out);
flip_bus #(1, 14) validIn_E_flip1(validIn_E, validIn_E_flip1_out);
flip_bus #(1, 14) validIn_S_flip1(validIn_S, validIn_S_flip1_out);
flip_bus #(1, 14) validIn_W_flip1(validIn_W, validIn_W_flip1_out);
flip_bus #(1, 10) validIn_N_flip2(validIn_N_flip1_out, validIn_N_internal);
flip_bus #(1, 10) validIn_E_flip2(validIn_E_flip1_out, validIn_E_internal);
flip_bus #(1, 10) validIn_S_flip2(validIn_S_flip1_out, validIn_S_internal);
flip_bus #(1, 10) validIn_W_flip2(validIn_W_flip1_out, validIn_W_internal);
flip_bus #(64, 14) dataIn_N_flip1(dataIn_N, dataIn_N_flip1_out);
flip_bus #(64, 14) dataIn_E_flip1(dataIn_E, dataIn_E_flip1_out);
flip_bus #(64, 14) dataIn_S_flip1(dataIn_S, dataIn_S_flip1_out);
flip_bus #(64, 14) dataIn_W_flip1(dataIn_W, dataIn_W_flip1_out);
flip_bus #(64, 10) dataIn_N_flip2(dataIn_N_flip1_out, dataIn_N_internal);
flip_bus #(64, 10) dataIn_E_flip2(dataIn_E_flip1_out, dataIn_E_internal);
flip_bus #(64, 10) dataIn_S_flip2(dataIn_S_flip1_out, dataIn_S_internal);
flip_bus #(64, 10) dataIn_W_flip2(dataIn_W_flip1_out, dataIn_W_internal);
dynamic_input_top_4 north_input(.route_req_n_out(route_req_n_to_n), .route_req_e_out(route_req_n_to_e), .route_req_s_out(route_req_n_to_s), .route_req_w_out(route_req_n_to_w), .route_req_p_out(route_req_n_to_p), .default_ready_n_out(), .default_ready_e_out(), .default_ready_s_out(default_ready_n_to_s), .default_ready_w_out(), .default_ready_p_out(), .tail_out(north_input_tail), .yummy_out(yummyOut_N_internal), .data_out(north_input_data), .valid_out(north_input_valid), .clk(clk), .reset(reset), .my_loc_x_in(myLocX_f), .my_loc_y_in(myLocY_f), .my_chip_id_in(myChipID_f), .valid_in(validIn_N_internal), .data_in(dataIn_N_internal), .thanks_n(thanks_n_to_n), .thanks_e(thanks_e_to_n), .thanks_s(thanks_s_to_n), .thanks_w(thanks_w_to_n), .thanks_p(thanks_p_to_n));
dynamic_input_top_4 east_input(.route_req_n_out(route_req_e_to_n), .route_req_e_out(route_req_e_to_e), .route_req_s_out(route_req_e_to_s), .route_req_w_out(route_req_e_to_w), .route_req_p_out(route_req_e_to_p), .default_ready_n_out(), .default_ready_e_out(), .default_ready_s_out(), .default_ready_w_out(default_ready_e_to_w), .default_ready_p_out(), .tail_out(east_input_tail), .yummy_out(yummyOut_E_internal), .data_out(east_input_data), .valid_out(east_input_valid), .clk(clk), .reset(reset), .my_loc_x_in(myLocX_f), .my_loc_y_in(myLocY_f), .my_chip_id_in(myChipID_f), .valid_in(validIn_E_internal), .data_in(dataIn_E_internal), .thanks_n(thanks_n_to_e), .thanks_e(thanks_e_to_e), .thanks_s(thanks_s_to_e), .thanks_w(thanks_w_to_e), .thanks_p(thanks_p_to_e));
dynamic_input_top_4 south_input(.route_req_n_out(route_req_s_to_n), .route_req_e_out(route_req_s_to_e), .route_req_s_out(route_req_s_to_s), .route_req_w_out(route_req_s_to_w), .route_req_p_out(route_req_s_to_p), .default_ready_n_out(default_ready_s_to_n), .default_ready_e_out(), .default_ready_s_out(), .default_ready_w_out(), .default_ready_p_out(default_ready_s_to_p), .tail_out(south_input_tail), .yummy_out(yummyOut_S_internal), .data_out(south_input_data), .valid_out(south_input_valid), .clk(clk), .reset(reset), .my_loc_x_in(myLocX_f), .my_loc_y_in(myLocY_f), .my_chip_id_in(myChipID_f), .valid_in(validIn_S_internal), .data_in(dataIn_S_internal), .thanks_n(thanks_n_to_s), .thanks_e(thanks_e_to_s), .thanks_s(thanks_s_to_s), .thanks_w(thanks_w_to_s), .thanks_p(thanks_p_to_s));
dynamic_input_top_4 west_input(.route_req_n_out(route_req_w_to_n), .route_req_e_out(route_req_w_to_e), .route_req_s_out(route_req_w_to_s), .route_req_w_out(route_req_w_to_w), .route_req_p_out(route_req_w_to_p), .default_ready_n_out(), .default_ready_e_out(default_ready_w_to_e), .default_ready_s_out(), .default_ready_w_out(), .default_ready_p_out(), .tail_out(west_input_tail), .yummy_out(yummyOut_W_internal), .data_out(west_input_data), .valid_out(west_input_valid), .clk(clk), .reset(reset), .my_loc_x_in(myLocX_f), .my_loc_y_in(myLocY_f), .my_chip_id_in(myChipID_f), .valid_in(validIn_W_internal), .data_in(dataIn_W_internal), .thanks_n(thanks_n_to_w), .thanks_e(thanks_e_to_w), .thanks_s(thanks_s_to_w), .thanks_w(thanks_w_to_w), .thanks_p(thanks_p_to_w));
dynamic_input_top_16 proc_input(.route_req_n_out(route_req_p_to_n), .route_req_e_out(route_req_p_to_e), .route_req_s_out(route_req_p_to_s), .route_req_w_out(route_req_p_to_w), .route_req_p_out(route_req_p_to_p), .default_ready_n_out(), .default_ready_e_out(), .default_ready_s_out(), .default_ready_w_out(), .default_ready_p_out(), .tail_out(proc_input_tail), .yummy_out(yummyOut_P_internal), .data_out(proc_input_data), .valid_out(proc_input_valid), .clk(clk), .reset(reset), .my_loc_x_in(myLocX_f), .my_loc_y_in(myLocY_f), .my_chip_id_in(myChipID_f), .valid_in(validIn_P), .data_in(dataIn_P), .thanks_n(thanks_n_to_p), .thanks_e(thanks_e_to_p), .thanks_s(thanks_s_to_p), .thanks_w(thanks_w_to_p), .thanks_p(thanks_p_to_p));
dynamic_output_top north_output(.data_out(dataOut_N_internal), .thanks_a_out(thanks_n_to_s), .thanks_b_out(thanks_n_to_w), .thanks_c_out(thanks_n_to_p), .thanks_d_out(thanks_n_to_e), .thanks_x_out(thanks_n_to_n), .valid_out(validOut_N_internal),  .popped_interrupt_mesg_out(), .popped_memory_ack_mesg_out(), .popped_memory_ack_mesg_out_sender(), .ec_wants_to_send_but_cannot(ec_wants_to_send_but_cannot_N), .clk(clk), .reset(reset), .route_req_a_in(route_req_s_to_n), .route_req_b_in(route_req_w_to_n), .route_req_c_in(route_req_p_to_n), .route_req_d_in(route_req_e_to_n), .route_req_x_in(route_req_n_to_n), .tail_a_in(south_input_tail), .tail_b_in(west_input_tail), .tail_c_in(proc_input_tail), .tail_d_in(east_input_tail), .tail_x_in(north_input_tail), .data_a_in(south_input_data), .data_b_in(west_input_data), .data_c_in(proc_input_data), .data_d_in(east_input_data), .data_x_in(north_input_data), .valid_a_in(south_input_valid), .valid_b_in(west_input_valid), .valid_c_in(proc_input_valid), .valid_d_in(east_input_valid), .valid_x_in(north_input_valid), .default_ready_in(default_ready_s_to_n), .yummy_in(yummyIn_N_internal));
dynamic_output_top east_output(.data_out(dataOut_E_internal), .thanks_a_out(thanks_e_to_w), .thanks_b_out(thanks_e_to_p), .thanks_c_out(thanks_e_to_n), .thanks_d_out(thanks_e_to_s), .thanks_x_out(thanks_e_to_e), .valid_out(validOut_E_internal),   .popped_interrupt_mesg_out(), .popped_memory_ack_mesg_out(), .popped_memory_ack_mesg_out_sender(),  .ec_wants_to_send_but_cannot(ec_wants_to_send_but_cannot_E), .clk(clk), .reset(reset), .route_req_a_in(route_req_w_to_e), .route_req_b_in(route_req_p_to_e), .route_req_c_in(route_req_n_to_e), .route_req_d_in(route_req_s_to_e), .route_req_x_in(route_req_e_to_e), .tail_a_in(west_input_tail), .tail_b_in(proc_input_tail), .tail_c_in(north_input_tail), .tail_d_in(south_input_tail), .tail_x_in(east_input_tail), .data_a_in(west_input_data), .data_b_in(proc_input_data), .data_c_in(north_input_data), .data_d_in(south_input_data), .data_x_in(east_input_data), .valid_a_in(west_input_valid), .valid_b_in(proc_input_valid), .valid_c_in(north_input_valid), .valid_d_in(south_input_valid), .valid_x_in(east_input_valid), .default_ready_in(default_ready_w_to_e), .yummy_in(yummyIn_E_internal));
dynamic_output_top south_output(.data_out(dataOut_S_internal), .thanks_a_out(thanks_s_to_n), .thanks_b_out(thanks_s_to_e), .thanks_c_out(thanks_s_to_w), .thanks_d_out(thanks_s_to_p), .thanks_x_out(thanks_s_to_s), .valid_out(validOut_S_internal),   .popped_interrupt_mesg_out(), .popped_memory_ack_mesg_out(), .popped_memory_ack_mesg_out_sender(),  .ec_wants_to_send_but_cannot(ec_wants_to_send_but_cannot_S), .clk(clk), .reset(reset), .route_req_a_in(route_req_n_to_s), .route_req_b_in(route_req_e_to_s), .route_req_c_in(route_req_w_to_s), .route_req_d_in(route_req_p_to_s), .route_req_x_in(route_req_s_to_s), .tail_a_in(north_input_tail), .tail_b_in(east_input_tail), .tail_c_in(west_input_tail), .tail_d_in(proc_input_tail), .tail_x_in(south_input_tail), .data_a_in(north_input_data), .data_b_in(east_input_data), .data_c_in(west_input_data), .data_d_in(proc_input_data), .data_x_in(south_input_data), .valid_a_in(north_input_valid), .valid_b_in(east_input_valid), .valid_c_in(west_input_valid), .valid_d_in(proc_input_valid), .valid_x_in(south_input_valid), .default_ready_in(default_ready_n_to_s), .yummy_in(yummyIn_S_internal));
dynamic_output_top west_output(.data_out(dataOut_W_internal), .thanks_a_out(thanks_w_to_e), .thanks_b_out(thanks_w_to_s), .thanks_c_out(thanks_w_to_p), .thanks_d_out(thanks_w_to_n), .thanks_x_out(thanks_w_to_w), .valid_out(validOut_W_internal),   .popped_interrupt_mesg_out(), .popped_memory_ack_mesg_out(), .popped_memory_ack_mesg_out_sender(),  .ec_wants_to_send_but_cannot(ec_wants_to_send_but_cannot_W), .clk(clk), .reset(reset), .route_req_a_in(route_req_e_to_w), .route_req_b_in(route_req_s_to_w), .route_req_c_in(route_req_p_to_w), .route_req_d_in(route_req_n_to_w), .route_req_x_in(route_req_w_to_w), .tail_a_in(east_input_tail), .tail_b_in(south_input_tail), .tail_c_in(proc_input_tail), .tail_d_in(north_input_tail), .tail_x_in(west_input_tail), .data_a_in(east_input_data), .data_b_in(south_input_data), .data_c_in(proc_input_data), .data_d_in(north_input_data), .data_x_in(west_input_data), .valid_a_in(east_input_valid), .valid_b_in(south_input_valid), .valid_c_in(proc_input_valid), .valid_d_in(north_input_valid), .valid_x_in(west_input_valid), .default_ready_in(default_ready_e_to_w), .yummy_in(yummyIn_W_internal));
dynamic_output_top #(1'b0) proc_output(.data_out(dataOut_P_internal), .thanks_a_out(thanks_p_to_s), .thanks_b_out(thanks_p_to_w), .thanks_c_out(thanks_p_to_n), .thanks_d_out(thanks_p_to_e), .thanks_x_out(thanks_p_to_p), .valid_out(validOut_P_internal),  .popped_interrupt_mesg_out(external_interrupt), .popped_memory_ack_mesg_out(store_ack_received), .popped_memory_ack_mesg_out_sender(store_ack_addr),  .ec_wants_to_send_but_cannot(ec_wants_to_send_but_cannot_P), .clk(clk), .reset(reset), .route_req_a_in(route_req_s_to_p), .route_req_b_in(route_req_w_to_p), .route_req_c_in(route_req_n_to_p), .route_req_d_in(route_req_e_to_p), .route_req_x_in(route_req_p_to_p), .tail_a_in(south_input_tail), .tail_b_in(west_input_tail), .tail_c_in(north_input_tail), .tail_d_in(east_input_tail), .tail_x_in(proc_input_tail), .data_a_in(south_input_data), .data_b_in(west_input_data), .data_c_in(north_input_data), .data_d_in(east_input_data), .data_x_in(proc_input_data), .valid_a_in(south_input_valid), .valid_b_in(west_input_valid), .valid_c_in(north_input_valid), .valid_d_in(east_input_valid), .valid_x_in(proc_input_valid), .default_ready_in(default_ready_s_to_p), .yummy_in(yummyIn_P_internal));
endmodule 
module dynamic_node_top_wrap_para
(
    input clk,
    input reset_in,
    
    input [64-1:0] dataIn_0,
    input [64-1:0] dataIn_1,
    input validIn_0,
    input validIn_1,
    input yummyIn_0,
    input yummyIn_1,
       
    input [8-1:0] myLocX,       
    input [8-1:0] myLocY,
    input [14-1:0] myChipID,
    
    output [64-1:0] dataOut_0,
    output [64-1:0] dataOut_1,
    output validOut_0,
    output validOut_1,
    output yummyOut_0,
    output yummyOut_1,
    
    
    output thanksIn_1      
);
    dynamic_node_top_para dynamic_node_top
    (
        .clk(clk),
        .reset_in(reset_in),
        
        .dataIn_0(dataIn_0),
        .dataIn_1(dataIn_1),
        .validIn_0(validIn_0),
        .validIn_1(validIn_1),
        .yummyIn_0(yummyIn_0),
        .yummyIn_1(yummyIn_1),
        .myLocX(myLocX),
        .myLocY(myLocY),
        .myChipID(myChipID),
        .ec_cfg(6'b0),
        .store_meter_partner_address_X(5'b0),
        .store_meter_partner_address_Y(5'b0),
        
        .dataOut_0(dataOut_0),
        .dataOut_1(dataOut_1),
        .validOut_0(validOut_0),
        .validOut_1(validOut_1),
        .yummyOut_0(yummyOut_0),
        .yummyOut_1(yummyOut_1),
        .thanksIn_1(thanksIn_1),
        .external_interrupt(),
        .store_meter_ack_partner(),
        .store_meter_ack_non_partner(),
        .ec_out()
    ); 
endmodule
module dynamic_node_top_para(clk,
		    reset_in,
        dataIn_0, dataIn_1, 
        validIn_0, validIn_1, 
        yummyIn_0,yummyIn_1,
		    myLocX,
		    myLocY,
            myChipID,
		    store_meter_partner_address_X,
		    store_meter_partner_address_Y,
		    ec_cfg,
        dataOut_0, dataOut_1, 
        validOut_0, validOut_1, 
        yummyOut_0,yummyOut_1,
		    thanksIn_1,
		    external_interrupt,
		    store_meter_ack_partner,
		    store_meter_ack_non_partner,
		    ec_out);
input clk;
input reset_in;
input [64-1:0] dataIn_0;
input [64-1:0] dataIn_1;
input validIn_0;
input validIn_1;
input yummyIn_0;
input yummyIn_1;
   
input [8-1:0] myLocX;		
input [8-1:0] myLocY;
input [14-1:0] myChipID;
input [4:0] store_meter_partner_address_X;
input [4:0] store_meter_partner_address_Y;
input [5:0] ec_cfg;            
output [64-1:0] dataOut_0;
output [64-1:0] dataOut_1;
output validOut_0;
output validOut_1;
output yummyOut_0;
output yummyOut_1;
output thanksIn_1;		
output external_interrupt;	
				
output store_meter_ack_partner;      
                                     
output store_meter_ack_non_partner;  
                                     
output [1:0] ec_out;
wire   ec_wants_to_send_but_cannot_0;
wire   ec_wants_to_send_but_cannot_1;
   wire store_ack_received;
   wire store_ack_received_r;
   wire [9:0] store_ack_addr;
   wire [9:0] store_ack_addr_r;
wire node_0_input_tail;
wire node_1_input_tail;
wire [64-1:0] node_0_input_data;
wire [64-1:0] node_1_input_data;
wire node_0_input_valid;
wire node_1_input_valid;
wire thanks_0_to_0;
wire thanks_0_to_1;
wire thanks_1_to_0;
wire thanks_1_to_1;
wire route_req_0_to_0;
wire route_req_0_to_1;
wire route_req_1_to_0;
wire route_req_1_to_1;
wire default_ready_0_to_0;
wire default_ready_0_to_1;
wire yummyOut_0_internal;
wire yummyOut_1_internal;
wire validOut_0_internal;
wire validOut_1_internal;
wire [64-1:0] dataOut_0_internal;
wire [64-1:0] dataOut_1_internal;
wire yummyOut_0_flip1_out;
wire validOut_0_flip1_out;
wire [64-1:0] dataOut_0_flip1_out;
wire yummyIn_0_internal;
wire yummyIn_1_internal;
wire validIn_0_internal;
wire [64-1:0] dataIn_0_internal;
wire yummyIn_0_flip1_out;
wire validIn_0_flip1_out;
wire [64-1:0] dataIn_0_flip1_out;
reg [8-1:0] myLocX_f;
reg [8-1:0] myLocY_f;
reg [14-1:0] myChipID_f;
wire   reset;
reg ec_thanks_0_to_0_reg, ec_thanks_0_to_1_reg;
reg ec_thanks_1_to_0_reg, ec_thanks_1_to_1_reg;
reg ec_wants_to_send_but_cannot_0_reg, ec_wants_to_send_but_cannot_1_reg;
reg ec_0_input_valid_reg, ec_1_input_valid_reg;
always @(posedge clk)
  begin
    
    ec_thanks_0_to_0_reg <= thanks_0_to_0; ec_thanks_0_to_1_reg <= thanks_0_to_1;
    ec_thanks_1_to_0_reg <= thanks_1_to_0; ec_thanks_1_to_1_reg <= thanks_1_to_1;
    ec_wants_to_send_but_cannot_0_reg <= ec_wants_to_send_but_cannot_0;
    ec_wants_to_send_but_cannot_1_reg <= ec_wants_to_send_but_cannot_1;
    ec_0_input_valid_reg <= node_0_input_valid;
    ec_1_input_valid_reg <= node_1_input_valid;
    
  end
wire ec_thanks_to_0= ec_thanks_0_to_0_reg | ec_thanks_1_to_0_reg ;
wire ec_thanks_to_1= ec_thanks_0_to_1_reg | ec_thanks_1_to_1_reg ;
one_of_n_plus_3 #(1) ec_mux_0(.in0(ec_wants_to_send_but_cannot_0),
                        .in1(ec_thanks_1_to_0_reg),
                        .in2(ec_thanks_0_to_0_reg),
                        .in3(ec_thanks_to_0),
                        .in4(ec_0_input_valid_reg & ~ec_thanks_to_0),
                        .sel(ec_cfg[5:3]),
                        .out(ec_out[1]));
one_of_n_plus_3 #(1) ec_mux_1(.in0(ec_wants_to_send_but_cannot_1),
                        .in1(ec_thanks_1_to_1_reg),
                        .in2(ec_thanks_0_to_1_reg),
                        .in3(ec_thanks_to_1),
                        .in4(ec_1_input_valid_reg & ~ec_thanks_to_1),
                        .sel(ec_cfg[2:0]),
                        .out(ec_out[0]));
net_dff #(1) REG_reset_fin(.d(reset_in), .q(reset), .clk(clk));
net_dff #(10) REG_store_ack_addr(   .d(store_ack_addr),     .q(store_ack_addr_r),     .clk(clk));
net_dff #(1) REG_store_ack_received(.d(store_ack_received), .q(store_ack_received_r), .clk(clk));
   wire is_partner_address_v_r;
   bus_compare_equal #(10) CMP_partner_address (.a(store_ack_addr_r),
                                        .b({ store_meter_partner_address_Y, store_meter_partner_address_X } ),
                                        .bus_equal(is_partner_address_v_r));
   assign store_meter_ack_partner     = is_partner_address_v_r & store_ack_received_r;
   assign store_meter_ack_non_partner = ~is_partner_address_v_r & store_ack_received_r;
always @ (posedge clk)
begin
        if(reset)
        begin
                myLocY_f <= 8'd0;
                myLocX_f <= 8'd0;
                myChipID_f <= 14'd0;
        end
        else
        begin
                myLocY_f <= myLocY;
                myLocX_f <= myLocX;
                myChipID_f <= myChipID;
        end
end
assign thanksIn_1 = thanks_0_to_1 | thanks_1_to_1 ;
assign validOut_1 = validOut_1_internal;
assign dataOut_1 = dataOut_1_internal;
assign yummyIn_1_internal = yummyIn_1;
assign yummyOut_1 = yummyOut_1_internal;
flip_bus #(1, 14) yummyOut_0_flip1(yummyOut_0_internal, yummyOut_0_flip1_out);
flip_bus #(1, 21) yummyOut_0_flip2(yummyOut_0_flip1_out, yummyOut_0);
flip_bus #(1, 14) validOut_0_flip1(validOut_0_internal, validOut_0_flip1_out);
flip_bus #(1, 21) validOut_0_flip2(validOut_0_flip1_out, validOut_0);
flip_bus #(64, 14) dataOut_0_flip1(dataOut_0_internal, dataOut_0_flip1_out);
flip_bus #(64, 21) dataOut_0_flip2(dataOut_0_flip1_out, dataOut_0);
flip_bus #(1, 14) yummyIn_0_flip1(yummyIn_0, yummyIn_0_flip1_out);
flip_bus #(1, 10) yummyIn_0_flip2(yummyIn_0_flip1_out, yummyIn_0_internal);
flip_bus #(1, 14) validIn_0_flip1(validIn_0, validIn_0_flip1_out);
flip_bus #(1, 10) validIn_0_flip2(validIn_0_flip1_out, validIn_0_internal);
flip_bus #(64, 14) dataIn_0_flip1(dataIn_0, dataIn_0_flip1_out);
flip_bus #(64, 10) dataIn_0_flip2(dataIn_0_flip1_out, dataIn_0_internal);
dynamic_input_top_4_para node_0_input(.route_req_0_out(route_req_0_to_0), .route_req_1_out(route_req_0_to_1), .default_ready_0_out(default_ready_0_to_0), .default_ready_1_out(default_ready_0_to_1), .tail_out(node_0_input_tail), .yummy_out(yummyOut_0_internal), .data_out(node_0_input_data), .valid_out(node_0_input_valid), .clk(clk), .reset(reset), .my_loc_x_in(myLocX_f), .my_loc_y_in(myLocY_f), .my_chip_id_in(myChipID_f), .valid_in(validIn_0_internal), .data_in(dataIn_0_internal), .thanks_0(thanks_0_to_0), .thanks_1(thanks_1_to_0));
dynamic_input_top_4_para node_1_input(.route_req_0_out(route_req_1_to_0), .route_req_1_out(route_req_1_to_1), .default_ready_0_out(), .default_ready_1_out(), .tail_out(node_1_input_tail), .yummy_out(yummyOut_1_internal), .data_out(node_1_input_data), .valid_out(node_1_input_valid), .clk(clk), .reset(reset), .my_loc_x_in(myLocX_f), .my_loc_y_in(myLocY_f), .my_chip_id_in(myChipID_f), .valid_in(validIn_1), .data_in(dataIn_1), .thanks_0(thanks_0_to_1), .thanks_1(thanks_1_to_1));
dynamic_output_top_para node_0_output(.data_out(dataOut_0_internal), .thanks_0_out(thanks_0_to_1), .thanks_1_out(thanks_0_to_0), .valid_out(validOut_0_internal), .popped_interrupt_mesg_out(), .popped_memory_ack_mesg_out(), .popped_memory_ack_mesg_out_sender(), .ec_wants_to_send_but_cannot(ec_wants_to_send_but_cannot_0), .clk(clk), .reset(reset), .route_req_0_in(route_req_1_to_0), .route_req_1_in(route_req_0_to_0), .tail_0_in(node_1_input_tail), .tail_1_in(node_0_input_tail), .data_0_in(node_1_input_data), .data_1_in(node_0_input_data), .valid_0_in(node_1_input_valid), .valid_1_in(node_0_input_valid), .default_ready_in(default_ready_0_to_0),.yummy_in(yummyIn_0_internal));
dynamic_output_top_para #(1'b0) node_1_output(.data_out(dataOut_1_internal), .thanks_0_out(thanks_1_to_0), .thanks_1_out(thanks_1_to_1), .valid_out(validOut_1_internal), .popped_interrupt_mesg_out(external_interrupt), .popped_memory_ack_mesg_out(store_ack_received), .popped_memory_ack_mesg_out_sender(store_ack_addr), .ec_wants_to_send_but_cannot(ec_wants_to_send_but_cannot_1), .clk(clk), .reset(reset), .route_req_0_in(route_req_0_to_1), .route_req_1_in(route_req_1_to_1), .tail_0_in(node_0_input_tail), .tail_1_in(node_1_input_tail), .data_0_in(node_0_input_data), .data_1_in(node_1_input_data), .valid_0_in(node_0_input_valid), .valid_1_in(node_1_input_valid), .default_ready_in(default_ready_0_to_1),.yummy_in(yummyIn_1_internal));
endmodule 
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
 
     
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	 
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
 
	
 
 
 
 
 
 
	
	
	
	
module l15 (
    input                                   clk,
    input                                   rst_n,
    
    input [4:0]                             transducer_l15_rqtype,
    input [4-1:0]           transducer_l15_amo_op,
    input                                   transducer_l15_nc,
    input [2:0]                             transducer_l15_size,
    input [0:0]              transducer_l15_threadid,
    input                                   transducer_l15_prefetch,
    input                                   transducer_l15_invalidate_cacheline,
    input                                   transducer_l15_blockstore,
    input                                   transducer_l15_blockinitstore,
    input [1:0]                             transducer_l15_l1rplway,
    input                                   transducer_l15_val,
    input [39:0]                            transducer_l15_address,
    input [63:0]                            transducer_l15_data,
    input [63:0]                            transducer_l15_data_next_entry,
    input [33-1:0]              transducer_l15_csm_data,
    output                                  l15_transducer_ack,
    output                                  l15_transducer_header_ack,
    output                                  l15_transducer_val,
    output [3:0]                            l15_transducer_returntype,
    output                                  l15_transducer_l2miss,
    output [1:0]                            l15_transducer_error,
    output                                  l15_transducer_noncacheable,
    output                                  l15_transducer_atomic,
    output [0:0]             l15_transducer_threadid,
    output                                  l15_transducer_prefetch,
    output                                  l15_transducer_f4b,
    output [63:0]                           l15_transducer_data_0,
    output [63:0]                           l15_transducer_data_1,
    output [63:0]                           l15_transducer_data_2,
    output [63:0]                           l15_transducer_data_3,
    output                                  l15_transducer_inval_icache_all_way,
    output                                  l15_transducer_inval_dcache_all_way,
    output [15:4]                           l15_transducer_inval_address_15_4,
    output                                  l15_transducer_cross_invalidate,
    output [1:0]                            l15_transducer_cross_invalidate_way,
    output                                  l15_transducer_inval_dcache_inval,
    output                                  l15_transducer_inval_icache_inval,
    output [1:0]                            l15_transducer_inval_way,
    output                                  l15_transducer_blockinitstore,
    input                                   transducer_l15_req_ack,
    input                                   noc1_out_rdy,
    input                                   noc2_in_val,
    input [64-1:0]             noc2_in_data,
    input                                   noc3_out_rdy,
    input                                   dmbr_l15_stall,
    input [14-1:0]           chipid,
    input [8-1:0]                coreid_x,
    input [8-1:0]                coreid_y,
    
    input [63:0]                            config_l15_read_res_data_s3,
    input                                   config_csm_en,
    input [31:0]                            config_system_tile_count,
    input [2-1:0]    config_home_alloc_method, 
    input [22-1:0]    config_hmt_base,
    output                                  noc1_out_val,
    output [64-1:0]            noc1_out_data,
    output                                  noc2_in_rdy,
    output                                  noc3_out_val,
    output [64-1:0]            noc3_out_data,
    output                                  l15_dmbr_l1missIn,
    output [4-1:0]            l15_dmbr_l1missTag,
    output                                  l15_dmbr_l2responseIn,
    output                                  l15_dmbr_l2missIn,
    output [4-1:0]            l15_dmbr_l2missTag,
    
    output                                  l15_config_req_val_s2,
    output                                  l15_config_req_rw_s2,
    output [63:0]                           l15_config_write_req_data_s2,
    output [15:8]       l15_config_req_address_s2,
    
    output [4-1:0]    srams_rtap_data,
    input  [4-1:0]             rtap_srams_bist_command,
    input  [4-1:0]    rtap_srams_bist_data
);
wire [4-1:0] dtag_rtap_data;
wire [4-1:0] dcache_rtap_data;
wire [4-1:0] hmt_rtap_data;
assign srams_rtap_data = dtag_rtap_data
                            | dcache_rtap_data
                            | hmt_rtap_data;
wire [40-1:0] l15_csm_req_address_s2;
wire l15_csm_req_val_s2;
wire l15_csm_stall_s3;
wire [3-1:0] l15_csm_req_ticket_s2;
wire  l15_csm_req_type_s2;
wire [127:0] l15_csm_req_data_s2;
wire  [33-1:0] l15_csm_req_pcx_data_s2;
wire csm_l15_res_val_s3;
wire [63:0] csm_l15_res_data_s3;
wire [3-1:0] l15_csm_read_ticket;
wire [3-1:0] l15_csm_clear_ticket;
wire l15_csm_clear_ticket_val;
wire [(14+8+8)-1:0] csm_l15_read_res_data;
wire csm_l15_read_res_val;
wire noc1encoder_csm_req_ack;
wire csm_noc1encoder_req_val;
wire [5-1:0] csm_noc1encoder_req_type;
wire [3-1:0] csm_noc1encoder_req_mshrid;
wire [40-1:0] csm_noc1encoder_req_address;
wire csm_noc1encoder_req_non_cacheable;
wire  [3-1:0] csm_noc1encoder_req_size;
l15_csm l15_csm(
    .clk(clk),
    .rst_n(rst_n),
    
    
    .l15_csm_read_ticket(l15_csm_read_ticket),
    .l15_csm_clear_ticket(l15_csm_clear_ticket),
    .l15_csm_clear_ticket_val(l15_csm_clear_ticket_val),
    .csm_l15_read_res_data(csm_l15_read_res_data),
    .csm_l15_read_res_val(csm_l15_read_res_val),
    
    
    .l15_hmt_base_reg(config_hmt_base),
    .csm_en(config_csm_en),
    .system_tile_count(config_system_tile_count[6-1:0]),
    .home_alloc_method(config_home_alloc_method),
    
    
    .l15_csm_req_address_s2(l15_csm_req_address_s2),
    .l15_csm_req_val_s2(l15_csm_req_val_s2),
    .l15_csm_stall_s3(l15_csm_stall_s3),
    .l15_csm_req_ticket_s2(l15_csm_req_ticket_s2),
    
    .l15_csm_req_type_s2(l15_csm_req_type_s2),
    .l15_csm_req_data_s2(l15_csm_req_data_s2),
    .l15_csm_req_pcx_data_s2(l15_csm_req_pcx_data_s2),
    .csm_l15_res_val_s3(csm_l15_res_val_s3),
    .csm_l15_res_data_s3(csm_l15_res_data_s3),
    
    
    .noc1encoder_csm_req_ack(noc1encoder_csm_req_ack),
    .csm_noc1encoder_req_val(csm_noc1encoder_req_val),
    .csm_noc1encoder_req_type(csm_noc1encoder_req_type),
    .csm_noc1encoder_req_mshrid(csm_noc1encoder_req_mshrid),
    .csm_noc1encoder_req_address(csm_noc1encoder_req_address),
    .csm_noc1encoder_req_non_cacheable(csm_noc1encoder_req_non_cacheable),
    .csm_noc1encoder_req_size(csm_noc1encoder_req_size)
);
wire [511:0] noc2_data;
wire noc2_data_val;
wire noc2_data_ack;
simplenocbuffer simplenocbuffer(
    .clk(clk),
    .rst_n(rst_n),
    .noc_in_val(noc2_in_val),
    .noc_in_data(noc2_in_data),
    .msg_ack(noc2_data_ack),
    .noc_in_rdy(noc2_in_rdy),
    .msg(noc2_data),
    .msg_val(noc2_data_val)
);
wire l15_noc2decoder_ack;
wire l15_noc2decoder_header_ack;
wire noc2decoder_l15_val;
wire [2-1:0] noc2decoder_l15_mshrid;
wire noc2decoder_l15_l2miss;
wire noc2decoder_l15_icache_type;
wire noc2decoder_l15_f4b;
wire [8-1:0] noc2decoder_l15_reqtype;
wire [2-1:0] noc2decoder_l15_ack_state;
wire [63:0] noc2decoder_l15_data_0;
wire [63:0] noc2decoder_l15_data_1;
wire [63:0] noc2decoder_l15_data_2;
wire [63:0] noc2decoder_l15_data_3;
wire [39:0] noc2decoder_l15_address;
wire [3:0] noc2decoder_l15_fwd_subcacheline_vector;
wire [(14+8+8)-1:0] noc2decoder_l15_src_homeid;
wire [3-1:0] noc2decoder_l15_csm_mshrid;
wire [0:0] noc2decoder_l15_threadid;
wire noc2decoder_l15_hmc_fill;
noc2decoder noc2decoder(
    .clk(clk),
    .rst_n(rst_n),
    .noc2_data(noc2_data),
    .noc2_data_val(noc2_data_val),
    .l15_noc2decoder_ack(l15_noc2decoder_ack),
    .l15_noc2decoder_header_ack(l15_noc2decoder_header_ack),
    .noc2_data_ack(noc2_data_ack),
    .noc2decoder_l15_val(noc2decoder_l15_val),
    .noc2decoder_l15_mshrid(noc2decoder_l15_mshrid),
    .noc2decoder_l15_l2miss(noc2decoder_l15_l2miss),
    .noc2decoder_l15_icache_type(noc2decoder_l15_icache_type),
    .noc2decoder_l15_f4b(noc2decoder_l15_f4b),
    .noc2decoder_l15_reqtype(noc2decoder_l15_reqtype),
    .noc2decoder_l15_ack_state(noc2decoder_l15_ack_state),
    .noc2decoder_l15_data_0(noc2decoder_l15_data_0),
    .noc2decoder_l15_data_1(noc2decoder_l15_data_1),
    .noc2decoder_l15_data_2(noc2decoder_l15_data_2),
    .noc2decoder_l15_data_3(noc2decoder_l15_data_3),
    .noc2decoder_l15_address(noc2decoder_l15_address),
    .noc2decoder_l15_fwd_subcacheline_vector(noc2decoder_l15_fwd_subcacheline_vector),
    .noc2decoder_l15_src_homeid(noc2decoder_l15_src_homeid),
    .noc2decoder_l15_csm_mshrid(noc2decoder_l15_csm_mshrid),
    .noc2decoder_l15_threadid(noc2decoder_l15_threadid),
    .noc2decoder_l15_hmc_fill(noc2decoder_l15_hmc_fill),
    .l15_dmbr_l2missIn(l15_dmbr_l2missIn),
    .l15_dmbr_l2missTag(l15_dmbr_l2missTag),
    .l15_dmbr_l2responseIn(l15_dmbr_l2responseIn)
);
wire noc1encoder_l15_req_ack;
wire noc1encoder_l15_req_sent;
wire l15_noc1buffer_req_val;
wire [2-1:0] noc1encoder_l15_req_data_sent;
wire [5-1:0] l15_noc1buffer_req_type;
wire [0:0] l15_noc1buffer_req_threadid;
wire [2-1:0] l15_noc1buffer_req_mshrid;
wire [39:0] l15_noc1buffer_req_address;
wire l15_noc1buffer_req_non_cacheable;
wire [2:0] l15_noc1buffer_req_size;
wire l15_noc1buffer_req_prefetch;
wire [63:0] l15_noc1buffer_req_data_0;
wire [63:0] l15_noc1buffer_req_data_1;
wire [33-1:0] l15_noc1buffer_req_csm_data;
wire [3-1:0] l15_noc1buffer_req_csm_ticket;
wire [(14+8+8)-1:0] l15_noc1buffer_req_homeid;
wire l15_noc1buffer_req_homeid_val;
wire [10-1:0] noc1buffer_noc1encoder_req_csm_sdid;
wire [6-1:0] noc1buffer_noc1encoder_req_csm_lsid;
wire [5-1:0] noc1buffer_noc1encoder_req_type;
wire [0:0] noc1buffer_noc1encoder_req_threadid;
wire [2-1:0] noc1buffer_noc1encoder_req_mshrid;
wire [39:0] noc1buffer_noc1encoder_req_address;
wire noc1buffer_noc1encoder_req_non_cacheable;
wire [2:0] noc1buffer_noc1encoder_req_size;
wire noc1buffer_noc1encoder_req_prefetch;
wire [63:0] noc1buffer_noc1encoder_req_data_0;
wire [63:0] noc1buffer_noc1encoder_req_data_1;
wire [(14+8+8)-1:0] noc1buffer_noc1encoder_req_homeid;
wire noc1encoder_noc1buffer_req_ack;
wire noc1buffer_noc1encoder_req_val;
wire noc3encoder_l15_req_ack;
wire noc3encoder_noc3buffer_req_ack;
wire l15_noc3encoder_req_val;
wire noc3buffer_noc3encoder_req_val;
wire [3-1:0] l15_noc3encoder_req_type;
wire [63:0] l15_noc3encoder_req_data_0;
wire [63:0] l15_noc3encoder_req_data_1;
wire [2-1:0] l15_noc3encoder_req_mshrid;
wire [1:0] l15_noc3encoder_req_sequenceid;
wire [0:0] l15_noc3encoder_req_threadid;
wire [39:0] l15_noc3encoder_req_address;
wire l15_noc3encoder_req_with_data;
wire l15_noc3encoder_req_was_inval;
wire [3:0] l15_noc3encoder_req_fwdack_vector;
wire [(14+8+8)-1:0] l15_noc3encoder_req_homeid;
wire [3-1:0] noc3buffer_noc3encoder_req_type;
wire [63:0] noc3buffer_noc3encoder_req_data_0;
wire [63:0] noc3buffer_noc3encoder_req_data_1;
wire [2-1:0] noc3buffer_noc3encoder_req_mshrid;
wire [1:0] noc3buffer_noc3encoder_req_sequenceid;
wire [0:0] noc3buffer_noc3encoder_req_threadid;
wire [39:0] noc3buffer_noc3encoder_req_address;
wire noc3buffer_noc3encoder_req_with_data;
wire noc3buffer_noc3encoder_req_was_inval;
wire [3:0] noc3buffer_noc3encoder_req_fwdack_vector;
wire [(14+8+8)-1:0] noc3buffer_noc3encoder_req_homeid;
wire l15_dtag_val_s1;
wire l15_dtag_rw_s1;
wire [((9-2))-1:0] l15_dtag_index_s1;
wire [33*4-1:0] l15_dtag_write_data_s1;
wire [33*4-1:0] l15_dtag_write_mask_s1;
wire [33*4-1:0] dtag_l15_dout_s2;
sram_l15_tag dtag(
    .MEMCLK(clk),
    .RESET_N(rst_n),
    .CE(l15_dtag_val_s1),
    .A(l15_dtag_index_s1),
    .DIN(l15_dtag_write_data_s1),
    .BW(l15_dtag_write_mask_s1),
    .RDWEN(l15_dtag_rw_s1),
    .DOUT(dtag_l15_dout_s2),
    .BIST_COMMAND(rtap_srams_bist_command),
    .BIST_DIN(rtap_srams_bist_data),
    .BIST_DOUT(dtag_rtap_data),
    .SRAMID(8'd6)
);
wire l15_dcache_val_s2;
wire l15_dcache_rw_s2;
wire [(((9-2))+2)-1:0] l15_dcache_index_s2;
wire [127:0] l15_dcache_write_data_s2;
wire [127:0] l15_dcache_write_mask_s2;
wire [127:0] dcache_l15_dout_s3;
wire [14 + 8 + 8-1:0] l15_hmt_write_data_s2;
wire [14 + 8 + 8-1:0] l15_hmt_write_mask_s2;
wire [14 + 8 + 8-1:0] hmt_l15_dout_s3;
sram_l15_data dcache(
    .MEMCLK(clk),
    .RESET_N(rst_n),
    .CE(l15_dcache_val_s2),
    .A(l15_dcache_index_s2),
    .DIN({l15_dcache_write_data_s2}),
    .BW({l15_dcache_write_mask_s2}),
    .RDWEN(l15_dcache_rw_s2),
    .DOUT({dcache_l15_dout_s3}),
    .BIST_COMMAND(rtap_srams_bist_command),
    .BIST_DIN(rtap_srams_bist_data),
    .BIST_DOUT(dcache_rtap_data),
    .SRAMID(8'd7)
);
wire [31:0] l15_hmt_write_data_s2_extended = l15_hmt_write_data_s2;
wire [31:0] l15_hmt_write_mask_s2_extended = l15_hmt_write_mask_s2;
wire [31:0] hmt_l15_dout_s3_extended;
assign hmt_l15_dout_s3 = hmt_l15_dout_s3_extended[14 + 8 + 8-1:0];
sram_l15_hmt hmt(
    .MEMCLK(clk),
    .RESET_N(rst_n),
    .CE(l15_dcache_val_s2),
    .A(l15_dcache_index_s2),
    .DIN(l15_hmt_write_data_s2_extended),
    .BW(l15_hmt_write_mask_s2_extended),
    .RDWEN(l15_dcache_rw_s2),
    .DOUT(hmt_l15_dout_s3_extended),
    .BIST_COMMAND(rtap_srams_bist_command),
    .BIST_DIN(rtap_srams_bist_data),
    .BIST_DOUT(hmt_rtap_data),
    .SRAMID(8'd8)
);
wire pipe_mshr_writereq_val_s1;
wire [3-1:0] pipe_mshr_writereq_op_s1;
wire [39:0] pipe_mshr_writereq_address_s1;
wire [127:0] pipe_mshr_writereq_write_buffer_data_s1;
wire [15:0] pipe_mshr_writereq_write_buffer_byte_mask_s1;
wire [((((((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) + 1) + 1) + 1)-1:0] pipe_mshr_writereq_control_s1;
wire [2-1:0] pipe_mshr_writereq_mshrid_s1;
wire [0:0] pipe_mshr_writereq_threadid_s1;
wire [0:0] pipe_mshr_readreq_threadid_s1;
wire [2-1:0] pipe_mshr_readreq_mshrid_s1;
wire [((((((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) + 1) + 1) + 1)-1:0] mshr_pipe_readres_control_s1;
wire [(14+8+8)-1:0] mshr_pipe_readres_homeid_s1;
wire [(4*2)-1:0] mshr_pipe_vals_s1;
wire [(40*2)-1:0] mshr_pipe_ld_address;
wire [(40*2)-1:0] mshr_pipe_st_address;
wire [(2*2)-1:0] mshr_pipe_st_way_s1;
wire [(2*2)-1:0] mshr_pipe_st_state_s1;
wire pipe_mshr_write_buffer_rd_en_s2;
wire [0:0] pipe_mshr_threadid_s2;
wire [127:0]mshr_pipe_write_buffer_s2;
wire [15:0] mshr_pipe_write_buffer_byte_mask_s2;
wire pipe_mshr_val_s3;
wire [3-1:0] pipe_mshr_op_s3;
wire [2-1:0] pipe_mshr_mshrid_s3;
wire [0:0] pipe_mshr_threadid_s3;
wire [2-1:0] pipe_mshr_write_update_state_s3;
wire [1:0] pipe_mshr_write_update_way_s3;
wire noc1buffer_mshr_homeid_write_val_s4;
wire [2-1:0] noc1buffer_mshr_homeid_write_mshrid_s4;
wire [(14+8+8)-1:0] noc1buffer_mshr_homeid_write_data_s4;
wire [0:0] noc1buffer_mshr_homeid_write_threadid_s4;
l15_mshr mshr(
    .clk(clk),
    .rst_n(rst_n),
    .pipe_mshr_writereq_val_s1(pipe_mshr_writereq_val_s1),
    .pipe_mshr_writereq_op_s1(pipe_mshr_writereq_op_s1),
    .pipe_mshr_writereq_address_s1(pipe_mshr_writereq_address_s1),
    .pipe_mshr_writereq_write_buffer_data_s1(pipe_mshr_writereq_write_buffer_data_s1),
    .pipe_mshr_writereq_write_buffer_byte_mask_s1(pipe_mshr_writereq_write_buffer_byte_mask_s1),
    .pipe_mshr_writereq_control_s1(pipe_mshr_writereq_control_s1),
    .pipe_mshr_writereq_mshrid_s1(pipe_mshr_writereq_mshrid_s1),
    .pipe_mshr_writereq_threadid_s1(pipe_mshr_writereq_threadid_s1),
    .pipe_mshr_readreq_threadid_s1(pipe_mshr_readreq_threadid_s1),
    .pipe_mshr_readreq_mshrid_s1(pipe_mshr_readreq_mshrid_s1),
    .mshr_pipe_readres_control_s1(mshr_pipe_readres_control_s1),
    .mshr_pipe_readres_homeid_s1(mshr_pipe_readres_homeid_s1),
    .mshr_pipe_vals_s1(mshr_pipe_vals_s1),
    .mshr_pipe_ld_address(mshr_pipe_ld_address),
    .mshr_pipe_st_address(mshr_pipe_st_address),
    .mshr_pipe_st_way_s1(mshr_pipe_st_way_s1),
    .mshr_pipe_st_state_s1(mshr_pipe_st_state_s1),
    .pipe_mshr_write_buffer_rd_en_s2(pipe_mshr_write_buffer_rd_en_s2),
    .pipe_mshr_threadid_s2(pipe_mshr_threadid_s2),
    .mshr_pipe_write_buffer_s2(mshr_pipe_write_buffer_s2),
    .mshr_pipe_write_buffer_byte_mask_s2(mshr_pipe_write_buffer_byte_mask_s2),
    .pipe_mshr_val_s3(pipe_mshr_val_s3),
    .pipe_mshr_op_s3(pipe_mshr_op_s3),
    .pipe_mshr_mshrid_s3(pipe_mshr_mshrid_s3),
    .pipe_mshr_threadid_s3(pipe_mshr_threadid_s3),
    .pipe_mshr_write_update_state_s3(pipe_mshr_write_update_state_s3),
    .pipe_mshr_write_update_way_s3(pipe_mshr_write_update_way_s3),
    
    .noc1buffer_mshr_homeid_write_threadid_s4(noc1buffer_mshr_homeid_write_threadid_s4),
    .noc1buffer_mshr_homeid_write_val_s4(noc1buffer_mshr_homeid_write_val_s4),
    .noc1buffer_mshr_homeid_write_mshrid_s4(noc1buffer_mshr_homeid_write_mshrid_s4),
    .noc1buffer_mshr_homeid_write_data_s4(noc1buffer_mshr_homeid_write_data_s4)
);
wire l15_mesi_read_val_s1;
wire [((9-2))-1:0] l15_mesi_read_index_s1;
wire l15_mesi_write_val_s2;
wire [((9-2))-1:0] l15_mesi_write_index_s2;
wire [7:0] l15_mesi_write_mask_s2;
wire [7:0] l15_mesi_write_data_s2;
wire [7:0] mesi_l15_dout_s2;
rf_l15_mesi mesi(
    .clk(clk),
    .rst_n(rst_n),
    .read_valid(l15_mesi_read_val_s1),
    .read_index(l15_mesi_read_index_s1),
    .write_valid(l15_mesi_write_val_s2),
    .write_index(l15_mesi_write_index_s2),
    .write_mask(l15_mesi_write_mask_s2),
    .write_data(l15_mesi_write_data_s2),
    .read_data(mesi_l15_dout_s2)
);
wire l15_lrsc_flag_read_val_s1;
wire [((9-2))-1:0] l15_lrsc_flag_read_index_s1;
wire l15_lrsc_flag_write_val_s2;
wire [((9-2))-1:0] l15_lrsc_flag_write_index_s2;
wire [3:0] l15_lrsc_flag_write_mask_s2;
wire [3:0] l15_lrsc_flag_write_data_s2;
wire [3:0] lrsc_flag_l15_dout_s2;
rf_l15_lrsc_flag lrsc_flag(
    .clk(clk),
    .rst_n(rst_n),
    .read_valid(l15_lrsc_flag_read_val_s1),
    .read_index(l15_lrsc_flag_read_index_s1),
    .write_valid(l15_lrsc_flag_write_val_s2),
    .write_index(l15_lrsc_flag_write_index_s2),
    .write_mask(l15_lrsc_flag_write_mask_s2),
    .write_data(l15_lrsc_flag_write_data_s2),
    .read_data(lrsc_flag_l15_dout_s2)
);
wire l15_wmt_read_val_s2;
wire [6:0] l15_wmt_read_index_s2;
wire l15_wmt_write_val_s3;
wire [6:0] l15_wmt_write_index_s3;
wire [4*((2+0)+1)-1:0] l15_wmt_write_mask_s3;
wire [4*((2+0)+1)-1:0] l15_wmt_write_data_s3;
wire [4*((2+0)+1)-1:0] wmt_l15_data_s3;
rf_l15_wmt wmc(
    .clk(clk),
    .rst_n(rst_n),
    .read_valid(l15_wmt_read_val_s2),
    .read_index(l15_wmt_read_index_s2),
    .write_valid(l15_wmt_write_val_s3),
    .write_index(l15_wmt_write_index_s3),
    .write_mask(l15_wmt_write_mask_s3),
    .write_data(l15_wmt_write_data_s3),
    .read_data(wmt_l15_data_s3)
);
wire l15_lruarray_read_val_s1;
wire [((9-2))-1:0] l15_lruarray_read_index_s1;
wire l15_lruarray_write_val_s3;
wire [((9-2))-1:0] l15_lruarray_write_index_s3;
wire [5:0] l15_lruarray_write_mask_s3;
wire [5:0] l15_lruarray_write_data_s3;
wire [5:0] lruarray_l15_dout_s2;
rf_l15_lruarray lruarray(
    .clk(clk),
    .rst_n(rst_n),
    .read_valid(l15_lruarray_read_val_s1),
    .read_index(l15_lruarray_read_index_s1),
    .write_valid(l15_lruarray_write_val_s3),
    .write_index(l15_lruarray_write_index_s3),
    .write_mask(l15_lruarray_write_mask_s3),
    .write_data(l15_lruarray_write_data_s3),
    .read_data(lruarray_l15_dout_s2)
);
l15_pipeline pipeline(
    .clk(clk),
    .rst_n(rst_n),
    .dtag_l15_dout_s2(dtag_l15_dout_s2),
    .dcache_l15_dout_s3(dcache_l15_dout_s3),
    .mesi_l15_dout_s2(mesi_l15_dout_s2),
    .lrsc_flag_l15_dout_s2(lrsc_flag_l15_dout_s2),
    .lruarray_l15_dout_s2(lruarray_l15_dout_s2),
    .wmt_l15_data_s3(wmt_l15_data_s3),
    .pcxdecoder_l15_rqtype               (transducer_l15_rqtype),
    .pcxdecoder_l15_amo_op               (transducer_l15_amo_op),
    .pcxdecoder_l15_nc                   (transducer_l15_nc),
    .pcxdecoder_l15_size                 (transducer_l15_size),
    
    .pcxdecoder_l15_threadid             (transducer_l15_threadid),
    .pcxdecoder_l15_prefetch             (transducer_l15_prefetch),
    .pcxdecoder_l15_blockstore           (transducer_l15_blockstore),
    .pcxdecoder_l15_blockinitstore       (transducer_l15_blockinitstore),
    .pcxdecoder_l15_l1rplway             (transducer_l15_l1rplway),
    .pcxdecoder_l15_val                  (transducer_l15_val),
    .pcxdecoder_l15_invalidate_cacheline (transducer_l15_invalidate_cacheline),
    .pcxdecoder_l15_address              (transducer_l15_address),
    .pcxdecoder_l15_data                 (transducer_l15_data),
    .pcxdecoder_l15_data_next_entry      (transducer_l15_data_next_entry),
    .pcxdecoder_l15_csm_data             (transducer_l15_csm_data),
    .noc2decoder_l15_val(noc2decoder_l15_val),
    .noc2decoder_l15_mshrid(noc2decoder_l15_mshrid),
    .noc2decoder_l15_l2miss(noc2decoder_l15_l2miss),
    .noc2decoder_l15_icache_type(noc2decoder_l15_icache_type),
    .noc2decoder_l15_f4b(noc2decoder_l15_f4b),
    .noc2decoder_l15_reqtype(noc2decoder_l15_reqtype),
    .noc2decoder_l15_ack_state(noc2decoder_l15_ack_state),
    .noc2decoder_l15_data_0(noc2decoder_l15_data_0),
    .noc2decoder_l15_data_1(noc2decoder_l15_data_1),
    .noc2decoder_l15_data_2(noc2decoder_l15_data_2),
    .noc2decoder_l15_data_3(noc2decoder_l15_data_3),
    .noc2decoder_l15_address(noc2decoder_l15_address),
    .noc2decoder_l15_fwd_subcacheline_vector(noc2decoder_l15_fwd_subcacheline_vector),
    .noc2decoder_l15_src_homeid(noc2decoder_l15_src_homeid),
    .noc2decoder_l15_csm_mshrid(noc2decoder_l15_csm_mshrid),
    .noc2decoder_l15_threadid(noc2decoder_l15_threadid),
    .noc2decoder_l15_hmc_fill(noc2decoder_l15_hmc_fill),
    .cpxencoder_l15_req_ack(transducer_l15_req_ack),
    
    .noc1encoder_l15_req_sent(noc1encoder_l15_req_sent),
    .noc1encoder_l15_req_data_sent(noc1encoder_l15_req_data_sent),
    .noc3encoder_l15_req_ack(noc3encoder_l15_req_ack),
    
    
    
    
    
    .l15_dtag_val_s1(l15_dtag_val_s1),
    .l15_dtag_rw_s1(l15_dtag_rw_s1),
    .l15_dtag_index_s1(l15_dtag_index_s1),
    .l15_dtag_write_data_s1(l15_dtag_write_data_s1),
    .l15_dtag_write_mask_s1(l15_dtag_write_mask_s1),
    .l15_dcache_val_s2(l15_dcache_val_s2),
    .l15_dcache_rw_s2(l15_dcache_rw_s2),
    .l15_dcache_index_s2(l15_dcache_index_s2),
    .l15_dcache_write_data_s2(l15_dcache_write_data_s2),
    .l15_dcache_write_mask_s2(l15_dcache_write_mask_s2),
    .l15_mesi_read_val_s1(l15_mesi_read_val_s1),
    .l15_mesi_read_index_s1(l15_mesi_read_index_s1),
    .l15_mesi_write_val_s2(l15_mesi_write_val_s2),
    .l15_mesi_write_index_s2(l15_mesi_write_index_s2),
    .l15_mesi_write_mask_s2(l15_mesi_write_mask_s2),
    .l15_mesi_write_data_s2(l15_mesi_write_data_s2),
    .l15_lrsc_flag_read_val_s1(l15_lrsc_flag_read_val_s1),
    .l15_lrsc_flag_read_index_s1(l15_lrsc_flag_read_index_s1),
    .l15_lrsc_flag_write_val_s2(l15_lrsc_flag_write_val_s2),
    .l15_lrsc_flag_write_index_s2(l15_lrsc_flag_write_index_s2),
    .l15_lrsc_flag_write_mask_s2(l15_lrsc_flag_write_mask_s2),
    .l15_lrsc_flag_write_data_s2(l15_lrsc_flag_write_data_s2),
    .l15_wmt_read_val_s2(l15_wmt_read_val_s2),
    .l15_wmt_read_index_s2(l15_wmt_read_index_s2),
    .l15_wmt_write_val_s3(l15_wmt_write_val_s3),
    .l15_wmt_write_index_s3(l15_wmt_write_index_s3),
    .l15_wmt_write_mask_s3(l15_wmt_write_mask_s3),
    .l15_wmt_write_data_s3(l15_wmt_write_data_s3),
    .l15_lruarray_read_val_s1(l15_lruarray_read_val_s1),
    .l15_lruarray_read_index_s1(l15_lruarray_read_index_s1),
    .l15_lruarray_write_val_s3(l15_lruarray_write_val_s3),
    .l15_lruarray_write_index_s3(l15_lruarray_write_index_s3),
    .l15_lruarray_write_mask_s3(l15_lruarray_write_mask_s3),
    .l15_lruarray_write_data_s3(l15_lruarray_write_data_s3),
    .l15_cpxencoder_val                  (l15_transducer_val),
    .l15_cpxencoder_returntype           (l15_transducer_returntype),
    .l15_cpxencoder_l2miss               (l15_transducer_l2miss),
    .l15_cpxencoder_error                (l15_transducer_error),
    .l15_cpxencoder_noncacheable         (l15_transducer_noncacheable),
    .l15_cpxencoder_atomic               (l15_transducer_atomic),
    .l15_cpxencoder_threadid             (l15_transducer_threadid),
    .l15_cpxencoder_prefetch             (l15_transducer_prefetch),
    .l15_cpxencoder_f4b                  (l15_transducer_f4b),
    .l15_cpxencoder_data_0               (l15_transducer_data_0),
    .l15_cpxencoder_data_1               (l15_transducer_data_1),
    .l15_cpxencoder_data_2               (l15_transducer_data_2),
    .l15_cpxencoder_data_3               (l15_transducer_data_3),
    .l15_cpxencoder_inval_icache_all_way (l15_transducer_inval_icache_all_way),
    .l15_cpxencoder_inval_dcache_all_way (l15_transducer_inval_dcache_all_way),
    .l15_cpxencoder_inval_address_15_4   (l15_transducer_inval_address_15_4),
    .l15_cpxencoder_cross_invalidate     (l15_transducer_cross_invalidate),
    .l15_cpxencoder_cross_invalidate_way (l15_transducer_cross_invalidate_way),
    .l15_cpxencoder_inval_dcache_inval   (l15_transducer_inval_dcache_inval),
    .l15_cpxencoder_inval_icache_inval   (l15_transducer_inval_icache_inval),
    .l15_cpxencoder_inval_way            (l15_transducer_inval_way),
    .l15_cpxencoder_blockinitstore       (l15_transducer_blockinitstore),
    .l15_noc1buffer_req_val(l15_noc1buffer_req_val),
    .l15_noc1buffer_req_type(l15_noc1buffer_req_type),
    .l15_noc1buffer_req_threadid(l15_noc1buffer_req_threadid),
    .l15_noc1buffer_req_mshrid(l15_noc1buffer_req_mshrid),
    .l15_noc1buffer_req_address(l15_noc1buffer_req_address),
    .l15_noc1buffer_req_non_cacheable(l15_noc1buffer_req_non_cacheable),
    .l15_noc1buffer_req_size(l15_noc1buffer_req_size),
    .l15_noc1buffer_req_prefetch(l15_noc1buffer_req_prefetch),
    
    
    .l15_noc1buffer_req_data_0(l15_noc1buffer_req_data_0),
    .l15_noc1buffer_req_data_1(l15_noc1buffer_req_data_1),
    .l15_noc1buffer_req_csm_data(l15_noc1buffer_req_csm_data),
    .l15_noc3encoder_req_val(l15_noc3encoder_req_val),
    .l15_noc3encoder_req_type(l15_noc3encoder_req_type),
    .l15_noc3encoder_req_data_0(l15_noc3encoder_req_data_0),
    .l15_noc3encoder_req_data_1(l15_noc3encoder_req_data_1),
    .l15_noc3encoder_req_mshrid(l15_noc3encoder_req_mshrid),
    .l15_noc3encoder_req_sequenceid(l15_noc3encoder_req_sequenceid),
    .l15_noc3encoder_req_threadid(l15_noc3encoder_req_threadid),
    .l15_noc3encoder_req_address(l15_noc3encoder_req_address),
    .l15_noc3encoder_req_with_data(l15_noc3encoder_req_with_data),
    .l15_noc3encoder_req_was_inval(l15_noc3encoder_req_was_inval),
    .l15_noc3encoder_req_fwdack_vector(l15_noc3encoder_req_fwdack_vector),
    .l15_noc3encoder_req_homeid(l15_noc3encoder_req_homeid),
    .l15_pcxdecoder_ack(l15_transducer_ack),
    .l15_noc2decoder_ack(l15_noc2decoder_ack),
    .l15_pcxdecoder_header_ack(l15_transducer_header_ack),
    .l15_noc2decoder_header_ack(l15_noc2decoder_header_ack),
    
    
    .l15_csm_req_address_s2(l15_csm_req_address_s2),
    .l15_csm_req_val_s2(l15_csm_req_val_s2),
    .l15_csm_stall_s3(l15_csm_stall_s3),
    .l15_csm_req_ticket_s2(l15_csm_req_ticket_s2),
    
    .l15_csm_req_type_s2(l15_csm_req_type_s2),
    .l15_csm_req_data_s2(l15_csm_req_data_s2),
    .l15_csm_req_pcx_data_s2(l15_csm_req_pcx_data_s2),
    .csm_l15_res_val_s3(csm_l15_res_val_s3),
    .csm_l15_res_data_s3(csm_l15_res_data_s3),
    
    .l15_noc1buffer_req_csm_ticket(l15_noc1buffer_req_csm_ticket),
    .l15_noc1buffer_req_homeid(l15_noc1buffer_req_homeid),
    .l15_noc1buffer_req_homeid_val(l15_noc1buffer_req_homeid_val),
    
    
    
    
     
    .l15_hmt_write_data_s2(l15_hmt_write_data_s2),
    .l15_hmt_write_mask_s2(l15_hmt_write_mask_s2),
    .hmt_l15_dout_s3(hmt_l15_dout_s3),
     
    
    
    .l15_config_req_val_s2(l15_config_req_val_s2),
    .l15_config_req_rw_s2(l15_config_req_rw_s2),
    .l15_config_write_req_data_s2(l15_config_write_req_data_s2),
    .l15_config_req_address_s2(l15_config_req_address_s2),
    .config_l15_read_res_data_s3(config_l15_read_res_data_s3),
    
    
    .pipe_mshr_writereq_val_s1(pipe_mshr_writereq_val_s1),
    .pipe_mshr_writereq_op_s1(pipe_mshr_writereq_op_s1),
    .pipe_mshr_writereq_address_s1(pipe_mshr_writereq_address_s1),
    .pipe_mshr_writereq_write_buffer_data_s1(pipe_mshr_writereq_write_buffer_data_s1),
    .pipe_mshr_writereq_write_buffer_byte_mask_s1(pipe_mshr_writereq_write_buffer_byte_mask_s1),
    .pipe_mshr_writereq_control_s1(pipe_mshr_writereq_control_s1),
    .pipe_mshr_writereq_mshrid_s1(pipe_mshr_writereq_mshrid_s1),
    .pipe_mshr_writereq_threadid_s1(pipe_mshr_writereq_threadid_s1),
    .pipe_mshr_readreq_threadid_s1(pipe_mshr_readreq_threadid_s1),
    .pipe_mshr_readreq_mshrid_s1(pipe_mshr_readreq_mshrid_s1),
    .mshr_pipe_readres_control_s1(mshr_pipe_readres_control_s1),
    .mshr_pipe_readres_homeid_s1(mshr_pipe_readres_homeid_s1),
    .mshr_pipe_vals_s1(mshr_pipe_vals_s1),
    .mshr_pipe_ld_address(mshr_pipe_ld_address),
    .mshr_pipe_st_address(mshr_pipe_st_address),
    .mshr_pipe_st_way_s1(mshr_pipe_st_way_s1),
    .mshr_pipe_st_state_s1(mshr_pipe_st_state_s1),
    .pipe_mshr_write_buffer_rd_en_s2(pipe_mshr_write_buffer_rd_en_s2),
    .pipe_mshr_threadid_s2(pipe_mshr_threadid_s2),
    .mshr_pipe_write_buffer_s2(mshr_pipe_write_buffer_s2),
    .mshr_pipe_write_buffer_byte_mask_s2(mshr_pipe_write_buffer_byte_mask_s2),
    .pipe_mshr_val_s3(pipe_mshr_val_s3),
    .pipe_mshr_op_s3(pipe_mshr_op_s3),
    .pipe_mshr_mshrid_s3(pipe_mshr_mshrid_s3),
    .pipe_mshr_threadid_s3(pipe_mshr_threadid_s3),
    .pipe_mshr_write_update_state_s3(pipe_mshr_write_update_state_s3),
    .pipe_mshr_write_update_way_s3(pipe_mshr_write_update_way_s3)
);
noc1buffer noc1buffer(
    .clk(clk),
    .rst_n(rst_n),
    .l15_noc1buffer_req_data_0(l15_noc1buffer_req_data_0),
    .l15_noc1buffer_req_data_1(l15_noc1buffer_req_data_1),
    .l15_noc1buffer_req_val(l15_noc1buffer_req_val),
    .l15_noc1buffer_req_type(l15_noc1buffer_req_type),
    .l15_noc1buffer_req_threadid(l15_noc1buffer_req_threadid),
    .l15_noc1buffer_req_mshrid(l15_noc1buffer_req_mshrid),
    .l15_noc1buffer_req_address(l15_noc1buffer_req_address),
    .l15_noc1buffer_req_non_cacheable(l15_noc1buffer_req_non_cacheable),
    .l15_noc1buffer_req_size(l15_noc1buffer_req_size),
    .l15_noc1buffer_req_prefetch(l15_noc1buffer_req_prefetch),
    
    
    .l15_noc1buffer_req_csm_data(l15_noc1buffer_req_csm_data),
    
    .l15_noc1buffer_req_csm_ticket(l15_noc1buffer_req_csm_ticket),
    .l15_noc1buffer_req_homeid(l15_noc1buffer_req_homeid),
    .l15_noc1buffer_req_homeid_val(l15_noc1buffer_req_homeid_val),
    .noc1buffer_noc1encoder_req_csm_sdid(noc1buffer_noc1encoder_req_csm_sdid),
    .noc1buffer_noc1encoder_req_csm_lsid(noc1buffer_noc1encoder_req_csm_lsid),
    
    .noc1encoder_noc1buffer_req_ack(noc1encoder_noc1buffer_req_ack),
    
    .noc1buffer_noc1encoder_req_data_0(noc1buffer_noc1encoder_req_data_0),
    .noc1buffer_noc1encoder_req_data_1(noc1buffer_noc1encoder_req_data_1),
    .noc1buffer_noc1encoder_req_val(noc1buffer_noc1encoder_req_val),
    .noc1buffer_noc1encoder_req_type(noc1buffer_noc1encoder_req_type),
    .noc1buffer_noc1encoder_req_mshrid(noc1buffer_noc1encoder_req_mshrid),
    .noc1buffer_noc1encoder_req_threadid(noc1buffer_noc1encoder_req_threadid),
    .noc1buffer_noc1encoder_req_address(noc1buffer_noc1encoder_req_address),
    .noc1buffer_noc1encoder_req_non_cacheable(noc1buffer_noc1encoder_req_non_cacheable),
    .noc1buffer_noc1encoder_req_size(noc1buffer_noc1encoder_req_size),
    .noc1buffer_noc1encoder_req_prefetch(noc1buffer_noc1encoder_req_prefetch),
    
    
    
    
    
    
    
    
    
    .l15_csm_read_ticket(l15_csm_read_ticket),
    .l15_csm_clear_ticket(l15_csm_clear_ticket),
    .l15_csm_clear_ticket_val(l15_csm_clear_ticket_val),
    .csm_l15_read_res_data(csm_l15_read_res_data),
    .csm_l15_read_res_val(csm_l15_read_res_val),
    .noc1buffer_noc1encoder_req_homeid(noc1buffer_noc1encoder_req_homeid),
    
    
    .noc1buffer_l15_req_sent(noc1encoder_l15_req_sent),
    .noc1buffer_l15_req_data_sent(noc1encoder_l15_req_data_sent),
    
    
    .noc1buffer_mshr_homeid_write_threadid_s4(noc1buffer_mshr_homeid_write_threadid_s4),
    .noc1buffer_mshr_homeid_write_val_s4(noc1buffer_mshr_homeid_write_val_s4),
    .noc1buffer_mshr_homeid_write_mshrid_s4(noc1buffer_mshr_homeid_write_mshrid_s4),
    .noc1buffer_mshr_homeid_write_data_s4(noc1buffer_mshr_homeid_write_data_s4)
);
noc1encoder noc1encoder(
    .clk(clk),
    .rst_n(rst_n),
    .noc1buffer_noc1encoder_req_data_0(noc1buffer_noc1encoder_req_data_0),
    .noc1buffer_noc1encoder_req_data_1(noc1buffer_noc1encoder_req_data_1),
    .noc1buffer_noc1encoder_req_val(noc1buffer_noc1encoder_req_val),
    .noc1buffer_noc1encoder_req_type(noc1buffer_noc1encoder_req_type),
    .noc1buffer_noc1encoder_req_mshrid(noc1buffer_noc1encoder_req_mshrid),
    .noc1buffer_noc1encoder_req_threadid(noc1buffer_noc1encoder_req_threadid),
    .noc1buffer_noc1encoder_req_address(noc1buffer_noc1encoder_req_address),
    .noc1buffer_noc1encoder_req_non_cacheable(noc1buffer_noc1encoder_req_non_cacheable),
    .noc1buffer_noc1encoder_req_size(noc1buffer_noc1encoder_req_size),
    .noc1buffer_noc1encoder_req_prefetch(noc1buffer_noc1encoder_req_prefetch),
    
    
    .noc1buffer_noc1encoder_req_csm_sdid(noc1buffer_noc1encoder_req_csm_sdid),
    .noc1buffer_noc1encoder_req_csm_lsid(noc1buffer_noc1encoder_req_csm_lsid),
    .noc1buffer_noc1encoder_req_homeid(noc1buffer_noc1encoder_req_homeid),
    
    .dmbr_l15_stall(dmbr_l15_stall),
    .chipid(chipid),
    .coreid_x(coreid_x),
    .coreid_y(coreid_y),
    .noc1out_ready(noc1_out_rdy),
    
    .l15_dmbr_l1missIn(l15_dmbr_l1missIn),
    .l15_dmbr_l1missTag(l15_dmbr_l1missTag),
    .noc1encoder_noc1buffer_req_ack(noc1encoder_noc1buffer_req_ack),
    .noc1encoder_noc1out_val(noc1_out_val),
    .noc1encoder_noc1out_data(noc1_out_data),
    
    
    .noc1encoder_csm_req_ack(noc1encoder_csm_req_ack),
    .csm_noc1encoder_req_val(csm_noc1encoder_req_val),
    .csm_noc1encoder_req_type(csm_noc1encoder_req_type),
    .csm_noc1encoder_req_mshrid(csm_noc1encoder_req_mshrid),
    .csm_noc1encoder_req_address(csm_noc1encoder_req_address),
    .csm_noc1encoder_req_non_cacheable(csm_noc1encoder_req_non_cacheable),
    .csm_noc1encoder_req_size(csm_noc1encoder_req_size)
);
noc3buffer noc3buffer(
    .clk(clk),
    .rst_n(rst_n),
    .l15_noc3encoder_req_val(l15_noc3encoder_req_val),
    .l15_noc3encoder_req_type(l15_noc3encoder_req_type),
    .l15_noc3encoder_req_data_0(l15_noc3encoder_req_data_0),
    .l15_noc3encoder_req_data_1(l15_noc3encoder_req_data_1),
    .l15_noc3encoder_req_mshrid(l15_noc3encoder_req_mshrid),
    .l15_noc3encoder_req_sequenceid(l15_noc3encoder_req_sequenceid),
    .l15_noc3encoder_req_threadid(l15_noc3encoder_req_threadid),
    .l15_noc3encoder_req_address(l15_noc3encoder_req_address),
    .l15_noc3encoder_req_with_data(l15_noc3encoder_req_with_data),
    .l15_noc3encoder_req_was_inval(l15_noc3encoder_req_was_inval),
    .l15_noc3encoder_req_fwdack_vector(l15_noc3encoder_req_fwdack_vector),
    .l15_noc3encoder_req_homeid(l15_noc3encoder_req_homeid),
    .noc3buffer_l15_req_ack(noc3encoder_l15_req_ack),
    
    
    .noc3buffer_noc3encoder_req_val(noc3buffer_noc3encoder_req_val),
    .noc3buffer_noc3encoder_req_type(noc3buffer_noc3encoder_req_type),
    .noc3buffer_noc3encoder_req_data_0(noc3buffer_noc3encoder_req_data_0),
    .noc3buffer_noc3encoder_req_data_1(noc3buffer_noc3encoder_req_data_1),
    .noc3buffer_noc3encoder_req_mshrid(noc3buffer_noc3encoder_req_mshrid),
    .noc3buffer_noc3encoder_req_sequenceid(noc3buffer_noc3encoder_req_sequenceid),
    .noc3buffer_noc3encoder_req_threadid(noc3buffer_noc3encoder_req_threadid),
    .noc3buffer_noc3encoder_req_address(noc3buffer_noc3encoder_req_address),
    .noc3buffer_noc3encoder_req_with_data(noc3buffer_noc3encoder_req_with_data),
    .noc3buffer_noc3encoder_req_was_inval(noc3buffer_noc3encoder_req_was_inval),
    .noc3buffer_noc3encoder_req_fwdack_vector(noc3buffer_noc3encoder_req_fwdack_vector),
    .noc3buffer_noc3encoder_req_homeid(noc3buffer_noc3encoder_req_homeid),
    .noc3encoder_noc3buffer_req_ack(noc3encoder_noc3buffer_req_ack)
);
noc3encoder noc3encoder(
    .clk(clk),
    .rst_n(rst_n),
    .l15_noc3encoder_req_val(noc3buffer_noc3encoder_req_val),
    .l15_noc3encoder_req_type(noc3buffer_noc3encoder_req_type),
    .l15_noc3encoder_req_data_0(noc3buffer_noc3encoder_req_data_0),
    .l15_noc3encoder_req_data_1(noc3buffer_noc3encoder_req_data_1),
    .l15_noc3encoder_req_mshrid(noc3buffer_noc3encoder_req_mshrid),
    .l15_noc3encoder_req_sequenceid(noc3buffer_noc3encoder_req_sequenceid),
    .l15_noc3encoder_req_threadid(noc3buffer_noc3encoder_req_threadid),
    .l15_noc3encoder_req_address(noc3buffer_noc3encoder_req_address),
    .l15_noc3encoder_req_with_data(noc3buffer_noc3encoder_req_with_data),
    .l15_noc3encoder_req_was_inval(noc3buffer_noc3encoder_req_was_inval),
    .l15_noc3encoder_req_fwdack_vector(noc3buffer_noc3encoder_req_fwdack_vector),
    .l15_noc3encoder_req_homeid(noc3buffer_noc3encoder_req_homeid),
    .chipid(chipid),
    .coreid_x(coreid_x),
    .coreid_y(coreid_y),
    .noc3out_ready(noc3_out_rdy),
    .noc3encoder_l15_req_ack(noc3encoder_noc3buffer_req_ack),
    .noc3encoder_noc3out_val(noc3_out_val),
    .noc3encoder_noc3out_data(noc3_out_data)
);
endmodule
module l15_cpxencoder(
    input wire          clk,
    input wire          rst_n,
    input wire          l15_cpxencoder_val,
    input wire [3:0]    l15_cpxencoder_returntype,
    input wire          l15_cpxencoder_l2miss,
    input wire [1:0]    l15_cpxencoder_error,
    input wire          l15_cpxencoder_noncacheable,
    input wire          l15_cpxencoder_atomic,
    input wire [0:0]    l15_cpxencoder_threadid,
    input wire          l15_cpxencoder_prefetch,
    input wire          l15_cpxencoder_f4b,
    input wire [63:0]  l15_cpxencoder_data_0,
    input wire [63:0]  l15_cpxencoder_data_1,
    input wire [63:0]  l15_cpxencoder_data_2,
    input wire [63:0]  l15_cpxencoder_data_3,
    input wire          l15_cpxencoder_inval_icache_all_way,
    input wire          l15_cpxencoder_inval_dcache_all_way,
    input wire [15:4]   l15_cpxencoder_inval_address_15_4,
    input wire          l15_cpxencoder_cross_invalidate,
    input wire [1:0]    l15_cpxencoder_cross_invalidate_way,
    input wire          l15_cpxencoder_inval_dcache_inval,
    input wire          l15_cpxencoder_inval_icache_inval,
    input wire [1:0]    l15_cpxencoder_inval_way,
    input wire          l15_cpxencoder_blockinitstore,
    output reg uncore_spc_data_ready,
    output reg [145-1:0] uncore_spc_data,
    output reg cpxencoder_l15_req_ack
    );
reg [145-1:0] out;
wire [2:0] cpuid = 3'b000;
reg state;
reg next_state;
reg [1:0] inval_index_5_4;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        state <= 1'b0;
    end
    else
    begin
        state <= next_state;
    end
end
always @ *
begin
    uncore_spc_data[145-1:0] = out[145-1:0];
    uncore_spc_data_ready = l15_cpxencoder_val;
    cpxencoder_l15_req_ack = (l15_cpxencoder_val && (next_state == 1'b0));
end
always @ *
begin
    out[144] = l15_cpxencoder_val;
    out[143:140] = l15_cpxencoder_returntype;
    out[139:0] = 1'b0;
    next_state = 1'b0;
    inval_index_5_4 = l15_cpxencoder_inval_address_15_4[5:4];
    if (l15_cpxencoder_val)
    begin
    case(l15_cpxencoder_returntype)
        4'b0000:
        begin
            
            out[139] = l15_cpxencoder_l2miss;
            out[138:137] = l15_cpxencoder_error;
            out[136] = l15_cpxencoder_noncacheable;
            out[135:134] = l15_cpxencoder_threadid;
            out[133] = l15_cpxencoder_cross_invalidate;
            out[132:131] = l15_cpxencoder_cross_invalidate_way;
            
            out[129] = l15_cpxencoder_atomic;
            out[128] = l15_cpxencoder_prefetch;
            out[127:0] = {l15_cpxencoder_data_0, l15_cpxencoder_data_1};
        end
        4'b0001:
        begin
            case (state)
                1'b0:
                begin
                    out[139] = l15_cpxencoder_l2miss;
                    out[138:137] = l15_cpxencoder_error;
                    out[136] = l15_cpxencoder_noncacheable;
                    out[135:134] = l15_cpxencoder_threadid;
                    out[133] = l15_cpxencoder_cross_invalidate;
                    out[132:131] = l15_cpxencoder_cross_invalidate_way;
                    out[130] = l15_cpxencoder_f4b;
                    out[129] = 1'b0;
                    out[128] = 1'b0;
                    out[127:0] = {l15_cpxencoder_data_0, l15_cpxencoder_data_1};
                    next_state = 1'b1;
                end
                1'b1:
                begin
                    
                    out[138:137] = l15_cpxencoder_error;
                    out[136] = l15_cpxencoder_noncacheable;
                    out[135:134] = l15_cpxencoder_threadid;
                    out[133] = l15_cpxencoder_cross_invalidate;
                    out[132:131] = l15_cpxencoder_cross_invalidate_way;
                    out[130] = 1'b0;
                    out[129] = 1'b1;
                    out[128] = 1'b0;
                    out[127:0] = {l15_cpxencoder_data_2, l15_cpxencoder_data_3};
                    next_state = 1'b0;
                end
            endcase
        end
        4'b0011:
        begin
            
            out[136] = l15_cpxencoder_noncacheable;
            out[128] = 1'b0;
            
                out[127:126] = 2'b0;
                out[125] = l15_cpxencoder_blockinitstore;
                out[124:123] = {l15_cpxencoder_inval_icache_all_way,
                                l15_cpxencoder_inval_dcache_all_way};
                out[122:121] = l15_cpxencoder_inval_address_15_4[5:4];
                out[120:118] = cpuid[2:0];
                out[117:112] = l15_cpxencoder_inval_address_15_4[11:6];
                
                if (l15_cpxencoder_inval_dcache_inval == 1)
                begin
                    out[5:2] = l15_cpxencoder_inval_way;
                    out[0] = 1'b1;
                end
                
        end
        4'b0100:
        begin
            out[136] = l15_cpxencoder_noncacheable;
            out[135:134] = l15_cpxencoder_threadid;
            out[129] = l15_cpxencoder_atomic;
            
                out[127:126] = 2'b0;
                out[125] = l15_cpxencoder_blockinitstore;
                out[124:123] = {l15_cpxencoder_inval_icache_all_way,
                                l15_cpxencoder_inval_dcache_all_way};
                out[122:121] = l15_cpxencoder_inval_address_15_4[5:4];
                out[120:118] = cpuid[2:0];
                out[117:112] = l15_cpxencoder_inval_address_15_4[11:6];
                
                if (l15_cpxencoder_inval_dcache_inval == 1)
                begin
                    out[5:2] = l15_cpxencoder_inval_way;
                    out[0] = 1'b1;
                end
        end
        4'b0111:
        begin
            
            
            
            out[136] = l15_cpxencoder_noncacheable; 
            out[63:0] = l15_cpxencoder_data_0;
            
            out[135:134] = l15_cpxencoder_threadid;
        end
        4'b1110:
        begin
            case (state)
                1'b0:
                begin
                    
                    out[143:140] = 4'b0000;
                    out[139] = l15_cpxencoder_l2miss;
                    out[138:137] = l15_cpxencoder_error;
                    out[136] = l15_cpxencoder_noncacheable;
                    out[135:134] = l15_cpxencoder_threadid;
                    out[133] = l15_cpxencoder_cross_invalidate;
                    out[132:131] = l15_cpxencoder_cross_invalidate_way;
                    
                    out[129] = l15_cpxencoder_atomic;
                    out[128] = l15_cpxencoder_prefetch;
                    out[127:0] = {l15_cpxencoder_data_0, l15_cpxencoder_data_1};
                    next_state = 1'b1;
                end
                1'b1:
                begin
                    
                    out[143:140] = 4'b0100;
                    out[136] = l15_cpxencoder_noncacheable;
                    out[135:134] = l15_cpxencoder_threadid;
                    out[129] = l15_cpxencoder_atomic;
                    
                        out[127:126] = 2'b0;
                        out[125] = l15_cpxencoder_blockinitstore;
                        out[124:123] = {l15_cpxencoder_inval_icache_all_way,
                                        l15_cpxencoder_inval_dcache_all_way};
                        out[122:121] = l15_cpxencoder_inval_address_15_4[5:4];
                        out[120:118] = cpuid[2:0];
                        out[117:112] = l15_cpxencoder_inval_address_15_4[11:6];
                        
                    next_state = 1'b0;
                end
            endcase
        end
        4'b1100:
        begin
            out[138:137] = l15_cpxencoder_error;
            out[135] = 1'b0;
            out[134] = 1'b0;
        end
        default:
        begin
            out[144] = 1'b0;
        end
    endcase
    end
end
endmodule
module l15_picoencoder(
    input wire          clk,
    input wire          rst_n,
    
    input wire          l15_picoencoder_val,
    input wire [3:0]    l15_picoencoder_returntype,
    
    input wire [63:0]   l15_picoencoder_data_0,
    input wire [63:0]   l15_picoencoder_data_1,
    
    input wire [39:0]   picodecoder_l15_address,  
    
    output reg          pico_mem_ready,
    output wire [31:0]  pico_mem_rdata,
    
    output wire         picoencoder_l15_req_ack,
    output reg          pico_int
);
    
    reg [31:0] rdata_part;
    assign pico_mem_rdata = {rdata_part[7:0], rdata_part[15:8],
                             rdata_part[23:16], rdata_part[31:24]};
    assign picoencoder_l15_req_ack = l15_picoencoder_val;
     
    
    reg int_recv;
    always @ (posedge clk) begin
        if (!rst_n) begin
            pico_int <= 1'b0;
        end
        else if (int_recv) begin
            pico_int <= 1'b1;
        end
        else if (pico_int) begin
            pico_int <= 1'b0;
        end
    end
       
    always @ * begin
        if (l15_picoencoder_val) begin
            case(l15_picoencoder_returntype)
                4'b0000, 4'b1110: begin
                    
                    int_recv = 1'b0;
                    pico_mem_ready = 1'b1;
                    case(picodecoder_l15_address[3:2])
                        2'b00: begin
                            rdata_part = l15_picoencoder_data_0[63:32];
                        end
                        2'b01: begin
                            rdata_part = l15_picoencoder_data_0[31:0];
                        end
                        2'b10: begin
                            rdata_part = l15_picoencoder_data_1[63:32];
                        end
                        2'b11: begin
                            rdata_part = l15_picoencoder_data_1[31:0];
                        end
                        default: begin
                        end
                    endcase 
                end
                4'b0100: begin
                    int_recv = 1'b0;
                    pico_mem_ready = 1'b1;
                    rdata_part = 32'b0;
                end
                4'b0111: begin
                    if (l15_picoencoder_data_0[17:16] == 2'b01) begin
                        int_recv = 1'b1;
                    end
                    else begin
                        int_recv = 1'b0;
                    end
                    pico_mem_ready = 1'b0;
                    rdata_part = 32'b0;
                end
                default: begin
                    int_recv = 1'b0;
                    pico_mem_ready = 1'b0;
                    rdata_part = 32'b0;
                end
            endcase 
        end
        else begin
            int_recv = 1'b0;
            pico_mem_ready = 1'b0;
            rdata_part = 32'b0;
        end
    end
    
endmodule 
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
module l15_wrap (
    input                                   clk,
    input                                   rst_n,
    input [4:0]                             transducer_l15_rqtype,
    input [4-1:0]           transducer_l15_amo_op,
    input                                   transducer_l15_nc,
    input [2:0]                             transducer_l15_size,
    input [0:0]              transducer_l15_threadid,
    input                                   transducer_l15_prefetch,
    input                                   transducer_l15_invalidate_cacheline,
    input                                   transducer_l15_blockstore,
    input                                   transducer_l15_blockinitstore,
    input [1:0]                             transducer_l15_l1rplway,
    input                                   transducer_l15_val,
    input [39:0]                            transducer_l15_address,
    input [63:0]                            transducer_l15_data,
    input [63:0]                            transducer_l15_data_next_entry,
    input [33-1:0]              transducer_l15_csm_data,
    output                                  l15_transducer_ack,
    output                                  l15_transducer_header_ack,
    output                                  l15_transducer_val,
    output [3:0]                            l15_transducer_returntype,
    output                                  l15_transducer_l2miss,
    output [1:0]                            l15_transducer_error,
    output                                  l15_transducer_noncacheable,
    output                                  l15_transducer_atomic,
    output [0:0]             l15_transducer_threadid,
    output                                  l15_transducer_prefetch,
    output                                  l15_transducer_f4b,
    output [63:0]                           l15_transducer_data_0,
    output [63:0]                           l15_transducer_data_1,
    output [63:0]                           l15_transducer_data_2,
    output [63:0]                           l15_transducer_data_3,
    output                                  l15_transducer_inval_icache_all_way,
    output                                  l15_transducer_inval_dcache_all_way,
    output [15:4]                           l15_transducer_inval_address_15_4,
    output                                  l15_transducer_cross_invalidate,
    output [1:0]                            l15_transducer_cross_invalidate_way,
    output                                  l15_transducer_inval_dcache_inval,
    output                                  l15_transducer_inval_icache_inval,
    output [1:0]                            l15_transducer_inval_way,
    output                                  l15_transducer_blockinitstore,
    input                                   transducer_l15_req_ack,
    input                                   noc1_out_rdy,
    input                                   noc2_in_val,
    input [64-1:0]             noc2_in_data,
    input                                   noc3_out_rdy,
    input                                   dmbr_l15_stall,
    input [14-1:0]           chipid,
    input [8-1:0]                coreid_x,
    input [8-1:0]                coreid_y,
    
    input [63:0]                            config_l15_read_res_data_s3,
    input                                   config_csm_en,
    input [5:0]                             config_system_tile_count_5_0,
    input [2-1:0]    config_home_alloc_method, 
    input [22-1:0]    config_hmt_base,
    output                                  noc1_out_val,
    output [64-1:0]            noc1_out_data,
    output                                  noc2_in_rdy,
    output                                  noc3_out_val,
    output [64-1:0]            noc3_out_data,
    
    output                                  l15_dmbr_l1missIn,
    output [4-1:0]            l15_dmbr_l1missTag,
    output                                  l15_dmbr_l2responseIn,
    output                                  l15_dmbr_l2missIn,
    output [4-1:0]            l15_dmbr_l2missTag,
    
    output                                  l15_config_req_val_s2,
    output                                  l15_config_req_rw_s2,
    output [63:0]                           l15_config_write_req_data_s2,
    output [15:8]       l15_config_req_address_s2,
    
    output [4-1:0]    srams_rtap_data,
    input  [4-1:0]             rtap_srams_bist_command,
    input  [4-1:0]    rtap_srams_bist_data
);
    wire [31:0]   config_system_tile_count = {26'bx, config_system_tile_count_5_0};
   
    l15 l15 (
        .clk(clk),
        .rst_n(rst_n),
        .transducer_l15_rqtype              (transducer_l15_rqtype),
        .transducer_l15_amo_op              (transducer_l15_amo_op),
        .transducer_l15_nc                  (transducer_l15_nc),
        .transducer_l15_size                (transducer_l15_size),
        
        .transducer_l15_threadid            (transducer_l15_threadid),
        .transducer_l15_prefetch            (transducer_l15_prefetch),
        .transducer_l15_blockstore          (transducer_l15_blockstore),
        .transducer_l15_blockinitstore      (transducer_l15_blockinitstore),
        .transducer_l15_l1rplway            (transducer_l15_l1rplway),
        .transducer_l15_val                 (transducer_l15_val),
        .transducer_l15_invalidate_cacheline(transducer_l15_invalidate_cacheline),
        .transducer_l15_address             (transducer_l15_address),
        .transducer_l15_csm_data            (transducer_l15_csm_data),
        .transducer_l15_data                (transducer_l15_data),
        .transducer_l15_data_next_entry     (transducer_l15_data_next_entry),
        .l15_transducer_ack                 (l15_transducer_ack),
        .l15_transducer_header_ack          (l15_transducer_header_ack),
                               
        .l15_transducer_val                 (l15_transducer_val),
        .l15_transducer_returntype          (l15_transducer_returntype),
        .l15_transducer_l2miss              (l15_transducer_l2miss),
        .l15_transducer_error               (l15_transducer_error),
        .l15_transducer_noncacheable        (l15_transducer_noncacheable),
        .l15_transducer_atomic              (l15_transducer_atomic),
        .l15_transducer_threadid            (l15_transducer_threadid),
        .l15_transducer_prefetch            (l15_transducer_prefetch),
        .l15_transducer_f4b                 (l15_transducer_f4b),
        .l15_transducer_data_0              (l15_transducer_data_0),
        .l15_transducer_data_1              (l15_transducer_data_1),
        .l15_transducer_data_2              (l15_transducer_data_2),
        .l15_transducer_data_3              (l15_transducer_data_3),
        .l15_transducer_inval_icache_all_way(l15_transducer_inval_icache_all_way),
        .l15_transducer_inval_dcache_all_way(l15_transducer_inval_dcache_all_way),
        .l15_transducer_inval_address_15_4  (l15_transducer_inval_address_15_4),
        .l15_transducer_cross_invalidate    (l15_transducer_cross_invalidate),
        .l15_transducer_cross_invalidate_way(l15_transducer_cross_invalidate_way),
        .l15_transducer_inval_dcache_inval  (l15_transducer_inval_dcache_inval),
        .l15_transducer_inval_icache_inval  (l15_transducer_inval_icache_inval),
        .l15_transducer_inval_way           (l15_transducer_inval_way),
        .l15_transducer_blockinitstore      (l15_transducer_blockinitstore),
        .transducer_l15_req_ack             (transducer_l15_req_ack),
        .noc1_out_rdy(noc1_out_rdy),
        .noc2_in_val(noc2_in_val),
        .noc2_in_data(noc2_in_data),
        .noc3_out_rdy(noc3_out_rdy),
        .dmbr_l15_stall(dmbr_l15_stall),
        .chipid(chipid),
        .coreid_x(coreid_x),
        .coreid_y(coreid_y),
        .noc1_out_val(noc1_out_val),
        .noc1_out_data(noc1_out_data),
        .noc2_in_rdy(noc2_in_rdy),
        .noc3_out_val(noc3_out_val),
        .noc3_out_data(noc3_out_data),
        
        .l15_dmbr_l1missIn(l15_dmbr_l1missIn),
        .l15_dmbr_l1missTag(l15_dmbr_l1missTag),
        .l15_dmbr_l2missIn(l15_dmbr_l2missIn),
        .l15_dmbr_l2missTag(l15_dmbr_l2missTag),
        .l15_dmbr_l2responseIn(l15_dmbr_l2responseIn),
        
        .l15_config_req_val_s2(l15_config_req_val_s2),
        .l15_config_req_rw_s2(l15_config_req_rw_s2),
        .l15_config_write_req_data_s2(l15_config_write_req_data_s2),
        .l15_config_req_address_s2(l15_config_req_address_s2),
        .config_l15_read_res_data_s3(config_l15_read_res_data_s3),
        
        .config_csm_en(config_csm_en),
        .config_hmt_base(config_hmt_base),
        .config_system_tile_count(config_system_tile_count),
        .config_home_alloc_method(config_home_alloc_method),
        
        
        .srams_rtap_data (srams_rtap_data),
        .rtap_srams_bist_command (rtap_srams_bist_command),
        .rtap_srams_bist_data (rtap_srams_bist_data)
    );
endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
module noc1encoder(
   input wire clk,
   input wire rst_n,
   
   input wire [63:0] noc1buffer_noc1encoder_req_data_0,
   input wire [63:0] noc1buffer_noc1encoder_req_data_1,
   input wire noc1buffer_noc1encoder_req_val,
   input wire [5-1:0] noc1buffer_noc1encoder_req_type,
   input wire [2-1:0] noc1buffer_noc1encoder_req_mshrid,
   input wire [0:0] noc1buffer_noc1encoder_req_threadid,
   input wire [39:0] noc1buffer_noc1encoder_req_address,
   input wire noc1buffer_noc1encoder_req_non_cacheable,
   input wire [3-1:0] noc1buffer_noc1encoder_req_size,
   input wire noc1buffer_noc1encoder_req_prefetch,
   
   
   input wire [(14+8+8)-1:0] noc1buffer_noc1encoder_req_homeid,
   input wire [10-1:0] noc1buffer_noc1encoder_req_csm_sdid,
   input wire [6-1:0] noc1buffer_noc1encoder_req_csm_lsid,
   output reg noc1encoder_noc1buffer_req_ack,
   
   input wire [14-1:0] chipid,
   input wire [8-1:0] coreid_x,
   input wire [8-1:0] coreid_y,
   
   input wire noc1out_ready,
   output reg noc1encoder_noc1out_val,
   output reg [63:0] noc1encoder_noc1out_data,
   
   input wire dmbr_l15_stall,
   output reg                       l15_dmbr_l1missIn,
   output reg [4-1:0] l15_dmbr_l1missTag,
   
   input wire csm_noc1encoder_req_val,
   input wire [5-1:0] csm_noc1encoder_req_type,
   input wire [3-1:0] csm_noc1encoder_req_mshrid,
   input wire [40-1:0] csm_noc1encoder_req_address,
   input wire csm_noc1encoder_req_non_cacheable,
   input wire  [3-1:0] csm_noc1encoder_req_size,
   output reg noc1encoder_csm_req_ack
);
reg [63:0] flit;
reg [4-1:0] flit_state;
reg [4-1:0] flit_state_next;
reg sending;
reg dmbr_stall;
reg control_raw_data_flit1;
always @ (posedge clk)
begin
   if (!rst_n)
   begin
      flit_state <= 0;
   end
   else
   begin
      flit_state <= flit_state_next;
   end
end
always @ *
begin
   
   noc1encoder_noc1out_data = flit;
   
   dmbr_stall = dmbr_l15_stall && (flit_state == 0); 
   sending = (noc1buffer_noc1encoder_req_val || csm_noc1encoder_req_val) && !dmbr_stall;
   noc1encoder_noc1out_val = sending;
end
reg [1-1:0] last_req_source;
reg [1-1:0] req_source;
reg [5-1:0] req_type;
reg req_prefetch;
reg req_nc;
reg [63:0] req_data0;
reg [63:0] req_data1;
reg [39:0] req_address;
reg [8-1:0] req_mshrid;
reg [3-1:0] req_size;
reg [8-1:0] req_dest_l2_xpos;
reg [8-1:0] req_dest_l2_ypos;
reg [14-1:0] req_dest_chipid;
reg [6-1:0] req_csm_lsid;
reg [10-1:0] req_csm_sdid;
always @ (posedge clk)
begin
   if (!rst_n)
      last_req_source <= 0;
   else
      last_req_source <= req_source;
end
always @ *
begin
   req_source = 0;
   req_type = 0;
   req_prefetch = 0;
   req_nc = 0;
   
   
   req_data0 = 0;
   req_data1 = 0;
   req_address = 0;
   req_mshrid = 0;
   req_size = 0;
   req_dest_l2_xpos = 0;
   req_dest_l2_ypos = 0;
   req_dest_chipid = 0;
   req_csm_lsid = 0;
   req_csm_sdid = 0;
   if ((last_req_source == 1'b0 && (flit_state != 0)) ||
         csm_noc1encoder_req_val == 1'b0)
   begin
      
      
      
      req_source = 1'b0;
   end
   else
   begin
      
      req_source = 1'b1;
   end
   if (req_source == 1'b0)
   begin
      req_type = noc1buffer_noc1encoder_req_type;
      req_prefetch = noc1buffer_noc1encoder_req_prefetch;
      req_nc = noc1buffer_noc1encoder_req_non_cacheable;
      
      
      req_data0 = noc1buffer_noc1encoder_req_data_0;
      req_data1 = noc1buffer_noc1encoder_req_data_1;
      req_address = noc1buffer_noc1encoder_req_address;
      req_mshrid = {noc1buffer_noc1encoder_req_threadid,noc1buffer_noc1encoder_req_mshrid};
      req_size = noc1buffer_noc1encoder_req_size;
      req_dest_l2_xpos = noc1buffer_noc1encoder_req_homeid[8-1:0];
      req_dest_l2_ypos = noc1buffer_noc1encoder_req_homeid[8+8-1:8];
      req_dest_chipid = noc1buffer_noc1encoder_req_homeid[((14+8+8)-1):(8+8)];
      if (req_type != 5'd1)
      begin
        req_csm_lsid = noc1buffer_noc1encoder_req_csm_lsid;
        req_csm_sdid = noc1buffer_noc1encoder_req_csm_sdid;
      end
   end
   else
   begin
      req_type = csm_noc1encoder_req_type;
      req_nc = csm_noc1encoder_req_non_cacheable;
      req_address = csm_noc1encoder_req_address;
      req_size = csm_noc1encoder_req_size;
      req_mshrid = csm_noc1encoder_req_mshrid;
      
      req_dest_l2_xpos = coreid_x;
      req_dest_l2_ypos = coreid_y;
      req_dest_chipid = chipid;
      
      req_mshrid = req_mshrid | {1'b1, {8-1{1'b0}}};
   end
end
reg [40-1:0]              msg_address;
reg [8-1:0]                 msg_dest_l2_xpos;
reg [8-1:0]                 msg_dest_l2_ypos;
reg [8-1:0]                 msg_dest_l2_xpos_new;
reg [8-1:0]                 msg_dest_l2_ypos_new;
wire [8-1:0]                msg_dest_l2_xpos_compat;
wire [8-1:0]                msg_dest_l2_ypos_compat;
reg [14-1:0]            msg_dest_chipid;
reg [4-1:0]             msg_dest_fbits;
reg [8-1:0]                 msg_src_xpos;
reg [8-1:0]                 msg_src_ypos;
reg [14-1:0]            msg_src_chipid;
reg [4-1:0]             msg_src_fbits;
reg [8-1:0]            msg_length;
reg [8-1:0]              msg_type;
reg [8-1:0]            msg_mshrid;
reg [2-1:0]               msg_mesi;
reg [1-1:0]      msg_last_subline;
reg [5:0]                   msg_options_1;
reg [15:0]                  msg_options_2;
reg [29:0]                  msg_options_3;
reg [1-1:0]        msg_cache_type;
reg [4-1:0]    msg_subline_vector;
reg [3-1:0]         msg_data_size;
reg [5:0] t1_interrupt_cpuid;
always @ *
begin
   msg_length = 0;
   msg_type = 0;
   msg_mesi = 0;
   msg_last_subline = 0;
   msg_cache_type = 0;
   msg_subline_vector = 0; 
   control_raw_data_flit1 = 0;
   t1_interrupt_cpuid = 0;
   msg_address = req_address;
   msg_mshrid = req_mshrid;
   msg_data_size = req_size;
   
   msg_src_xpos = coreid_x;
   msg_src_ypos = coreid_y;
   msg_src_chipid = chipid;
   msg_src_fbits = 4'd0;
   msg_dest_fbits = 4'd0;
   
   msg_dest_l2_xpos = req_dest_l2_xpos;
   msg_dest_l2_ypos = req_dest_l2_ypos;
   msg_dest_chipid = req_dest_chipid;
   
   msg_dest_l2_xpos_new = 0;
   msg_dest_l2_ypos_new = 0;
   case (req_type)
      5'd1:
      begin
         msg_type = 8'd13;
         msg_length = 2; 
         msg_cache_type = 1'b0;
      end
      5'd2:
      begin
         
         
         if (req_prefetch)
            msg_type = 8'd1;
         else if (req_nc)
            msg_type = 8'd14;
         else
            msg_type = 8'd31;
         msg_length = 2; 
         msg_cache_type = 1'b0;
      end
      5'd3:
      begin
         
         if (req_nc)
            msg_type = 8'd14;
         else
            msg_type = 8'd31;
         msg_length = 2; 
         msg_cache_type = 1'b1;
      end
      5'd4:
      begin
         
         if (req_nc)
            msg_type = 8'd15;
         
            
         
            
         msg_cache_type = 1'b0;
         msg_length = 3; 
      end
      5'd5, 5'd6:
      begin
         
         
         msg_type = 8'd2;
         msg_cache_type = 1'b0;
         msg_length = 2; 
      end
      5'd7:
      begin
         msg_type = 8'd5;
         msg_cache_type = 1'b0;
         msg_length = 4; 
      end
      5'd8:
      begin
         msg_type = 8'd9;
         msg_cache_type = 1'b0;
         msg_length = 3; 
      end
      5'd9:
      begin
         msg_type = 8'd32;
         msg_length = 1; 
         control_raw_data_flit1 = 1'b1;
         t1_interrupt_cpuid = req_data0[14:9];
         msg_dest_l2_xpos_new = req_data0[8+17:18];
         msg_dest_l2_ypos_new = req_data0[8+8+17:8+18];
         msg_dest_l2_xpos = req_data0[63] ? msg_dest_l2_xpos_new : msg_dest_l2_xpos_compat; 
         msg_dest_l2_ypos = req_data0[63] ? msg_dest_l2_ypos_new : msg_dest_l2_ypos_compat; 
         msg_dest_chipid  = req_data0[63] ? req_data0[14+8+8+17:8+8+18] : 14'b0;
      end
      5'd18:
      begin
         msg_type = 8'd60;
         msg_length = 2; 
         msg_cache_type = 1'b0;
      end
      5'd10:
      begin
         msg_type = 8'd36;
         msg_cache_type = 1'b0;
         msg_length = 3; 
      end
      5'd11:
      begin
         msg_type = 8'd37;
         msg_cache_type = 1'b0;
         msg_length = 3; 
      end
      5'd12:
      begin
         msg_type = 8'd38;
         msg_cache_type = 1'b0;
         msg_length = 3; 
      end
      5'd13:
      begin
         msg_type = 8'd39;
         msg_cache_type = 1'b0;
         msg_length = 3; 
      end
      5'd14:
      begin
         msg_type = 8'd40;
         msg_cache_type = 1'b0;
         msg_length = 3; 
      end
      5'd15:
      begin
         msg_type = 8'd41;
         msg_cache_type = 1'b0;
         msg_length = 3; 
      end
      5'd16:
      begin
         msg_type = 8'd42;
         msg_cache_type = 1'b0;
         msg_length = 3; 
      end
      5'd17:
      begin
         msg_type = 8'd43;
         msg_cache_type = 1'b0;
         msg_length = 3; 
      end
   endcase
end
flat_id_to_xy cpuid_to_xy (
    .flat_id(t1_interrupt_cpuid),
    .x_coord(msg_dest_l2_xpos_compat),
    .y_coord(msg_dest_l2_ypos_compat)
    );
always @ *
begin
   msg_options_1 = 0;
   msg_options_2 = 0;
   msg_options_3 = 0;
   msg_options_2[10:8] = msg_data_size;
   msg_options_2[11] = msg_cache_type;
   msg_options_2[15:12] = msg_subline_vector;
   msg_options_3[29:20] = req_csm_sdid;
   msg_options_3[19:14] = req_csm_lsid;
end
always @ *
begin
   flit[64-1:0] = 0; 
   if (flit_state == 4'd0)
   begin
      flit[63:50] = msg_dest_chipid;
      flit[49:42] = msg_dest_l2_xpos;
      flit[41:34] = msg_dest_l2_ypos;
      flit[33:30] = msg_dest_fbits;
      flit[29:22] = msg_length;
      flit[21:14] = msg_type;
      flit[13:6] = msg_mshrid;
      flit[5:0] = msg_options_1;
   end
   else if (flit_state == 4'd1)
   begin
      if (control_raw_data_flit1)
      begin
         flit[64-1:0] = req_data0;
         
         flit[15:9] = 0;
      end
      else
      begin
         flit[((16 + 40 - 1)):(16)] = msg_address;
         flit[11] = msg_cache_type;
         flit[15:0] = msg_options_2;
      end
   end
   else if (flit_state == 4'd2)
   begin
      flit[63:50] = msg_src_chipid;
      flit[49:42] = msg_src_xpos;
      flit[41:34] = msg_src_ypos;
      flit[33:30] = msg_src_fbits;
      flit[29:0] = msg_options_3;
   end
   else if (flit_state == 4'd3)
   begin
      flit[64-1:0] = req_data0;
   end
   else if (flit_state == 4'd4)
   begin
      flit[64-1:0] = req_data1;
   end
end
always @ *
begin
   
   if (sending)
   begin
      if (noc1out_ready)
      begin
         if (flit_state != msg_length)
            flit_state_next = flit_state + 1;
         else
            flit_state_next = 4'd0;
      end
      else
         flit_state_next = flit_state;
   end
   else
      flit_state_next = 4'd0;
end
always @ *
begin
   
   noc1encoder_noc1buffer_req_ack = 0;
   if (noc1buffer_noc1encoder_req_val && (flit_state == msg_length) && noc1out_ready
   && (req_source == 1'b0))
      noc1encoder_noc1buffer_req_ack = 1'b1;
   else
      noc1encoder_noc1buffer_req_ack = 1'b0;
   
   noc1encoder_csm_req_ack = 0;
   if (csm_noc1encoder_req_val && (flit_state == msg_length) && noc1out_ready 
   && (req_source == 1'b1))
      noc1encoder_csm_req_ack = 1'b1;
   else
      noc1encoder_csm_req_ack = 1'b0;
end
always @ *
begin
   
   l15_dmbr_l1missIn = 0;
   l15_dmbr_l1missTag = 0;
   
   
   
   if (noc1encoder_noc1buffer_req_ack)
   begin
      if (req_type == 5'd2 ||
         req_type == 5'd3 ||
         req_type == 5'd5 ||
         req_type == 5'd6 ||
         req_type == 5'd7 ||
         req_type == 5'd8 ||
         req_type == 5'd10 ||
         req_type == 5'd11 ||
         req_type == 5'd12 ||
         req_type == 5'd13 ||
         req_type == 5'd14 ||
         req_type == 5'd15 ||
         req_type == 5'd16 ||
         req_type == 5'd17)
      begin
         l15_dmbr_l1missIn = 1'b1;
         l15_dmbr_l1missTag = msg_mshrid[4-1:0]; 
      end
   end
end
endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
module noc2decoder(
    input wire clk,
    input wire rst_n,
    input wire [511:0] noc2_data,
    input wire noc2_data_val,
    input wire l15_noc2decoder_ack,
    input wire l15_noc2decoder_header_ack,
    output reg noc2_data_ack,
    output reg                       l15_dmbr_l2responseIn,
    output reg                       l15_dmbr_l2missIn,
    output reg [4-1:0] l15_dmbr_l2missTag,
    output reg noc2decoder_l15_val,
    output reg [2-1:0] noc2decoder_l15_mshrid,
    output reg [0:0] noc2decoder_l15_threadid,
    output reg noc2decoder_l15_hmc_fill,
    output reg noc2decoder_l15_l2miss,
    output reg noc2decoder_l15_icache_type,
    output reg noc2decoder_l15_f4b,
    output reg [8-1:0] noc2decoder_l15_reqtype,
    output reg [2-1:0] noc2decoder_l15_ack_state,
    output reg [63:0] noc2decoder_l15_data_0,
    output reg [63:0] noc2decoder_l15_data_1,
    output reg [63:0] noc2decoder_l15_data_2,
    output reg [63:0] noc2decoder_l15_data_3,
    output reg [39:0] noc2decoder_l15_address,
    output reg [3:0] noc2decoder_l15_fwd_subcacheline_vector,
    output reg [3-1:0] noc2decoder_l15_csm_mshrid,
    output reg [(14+8+8)-1:0] noc2decoder_l15_src_homeid
    );
reg is_message_new;
reg is_message_new_next;
always @ (posedge clk)
begin
    if (!rst_n)
      is_message_new <= 1'b1;
    else
      is_message_new <= is_message_new_next;
end
reg [8-1:0] noc2_mshrid;
reg [8-1:0] msg_len;
always @ *
begin
    noc2_data_ack = l15_noc2decoder_ack;
    noc2decoder_l15_val = noc2_data_val && is_message_new;
    
    noc2decoder_l15_reqtype = noc2_data[21:14];
    msg_len = noc2_data[29:22];
    
    noc2_mshrid = noc2_data[13:6];
    noc2decoder_l15_mshrid = noc2_mshrid[2-1:0];
    noc2decoder_l15_csm_mshrid = noc2_mshrid[3-1:0];
    
    noc2decoder_l15_threadid = noc2_mshrid[2+1 -1 -: 1];
    noc2decoder_l15_hmc_fill = noc2_mshrid[8-1];
    noc2decoder_l15_l2miss = noc2_data[3];
    noc2decoder_l15_icache_type = noc2_data[75];
    noc2decoder_l15_f4b = 0;
    noc2decoder_l15_ack_state = noc2_data[5:4];
    noc2decoder_l15_fwd_subcacheline_vector = noc2_data[79:76];
    noc2decoder_l15_address = noc2_data[119:80];
    
    
    
    
    
    
    
    noc2decoder_l15_data_0 = noc2_data[2*64 - 1 -: 64];
    noc2decoder_l15_data_1 = (msg_len == 8'd1) ? noc2_data[2*64 - 1 -: 64] : noc2_data[3*64 - 1 -: 64];
    noc2decoder_l15_data_2 = (msg_len <= 8'd2) ? noc2_data[2*64 - 1 -: 64] : noc2_data[4*64 - 1 -: 64];
    noc2decoder_l15_data_3 = (msg_len == 8'd1) ? noc2_data[2*64 - 1 -: 64] :
                                    (msg_len == 8'd2) ? noc2_data[3*64 - 1 -: 64] : noc2_data[5*64 - 1 -: 64];
    noc2decoder_l15_src_homeid = 0;
    noc2decoder_l15_src_homeid[8+8-1:8] = noc2_data[169:162];
    noc2decoder_l15_src_homeid[8-1:0] = noc2_data[177:170];
    noc2decoder_l15_src_homeid[((14+8+8)-1):(8+8)] = noc2_data[191:178];
    
    
    
    is_message_new_next = l15_noc2decoder_ack ? 1'b1 :
                                 l15_noc2decoder_header_ack ? 1'b0 : is_message_new;
end
reg dmbr_response_val_next;
reg dmbr_l2_miss_next;
reg [4-1:0]dmbr_l2_miss_mshrid_next;
reg dmbr_response_val;
reg dmbr_l2_miss;
reg [4-1:0]dmbr_l2_miss_mshrid;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        dmbr_response_val = 0;
        dmbr_l2_miss = 0;
        dmbr_l2_miss_mshrid = 0;
    end
    else
    begin
        dmbr_response_val = dmbr_response_val_next;
        dmbr_l2_miss = dmbr_l2_miss_next;
        dmbr_l2_miss_mshrid = dmbr_l2_miss_mshrid_next;
    end
end
always @ *
begin
    
    dmbr_response_val_next = 0;
    dmbr_l2_miss_next = 0;
    dmbr_l2_miss_mshrid_next = 0;
    if (l15_noc2decoder_ack)
    begin
        if (noc2decoder_l15_reqtype == 8'd29)
        begin
            dmbr_response_val_next = 1'b1;
            dmbr_l2_miss_next = noc2decoder_l15_l2miss;
            dmbr_l2_miss_mshrid_next = {1'b0, noc2decoder_l15_threadid, noc2decoder_l15_mshrid};
        end
    end
    l15_dmbr_l2responseIn = dmbr_response_val;
    l15_dmbr_l2missIn = dmbr_l2_miss;
    l15_dmbr_l2missTag = dmbr_l2_miss_mshrid;
end
endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
 
module noc3buffer(
    input wire clk,
    input wire rst_n,
    input wire l15_noc3encoder_req_val,
    input wire [3-1:0] l15_noc3encoder_req_type,
    input wire [63:0] l15_noc3encoder_req_data_0,
    input wire [63:0] l15_noc3encoder_req_data_1,
    input wire [2-1:0] l15_noc3encoder_req_mshrid,
    input wire [0:0] l15_noc3encoder_req_threadid,
    input wire [1:0] l15_noc3encoder_req_sequenceid,
    input wire [39:0] l15_noc3encoder_req_address,
    input wire l15_noc3encoder_req_with_data,
    input wire l15_noc3encoder_req_was_inval,
    input wire [3:0] l15_noc3encoder_req_fwdack_vector,
    input wire [(14+8+8)-1:0] l15_noc3encoder_req_homeid,
    output reg noc3buffer_noc3encoder_req_val,
    output reg [3-1:0] noc3buffer_noc3encoder_req_type,
    output reg [63:0] noc3buffer_noc3encoder_req_data_0,
    output reg [63:0] noc3buffer_noc3encoder_req_data_1,
    output reg [2-1:0] noc3buffer_noc3encoder_req_mshrid,
    output reg [1:0] noc3buffer_noc3encoder_req_sequenceid,
    output reg [0:0] noc3buffer_noc3encoder_req_threadid,
    output reg [39:0] noc3buffer_noc3encoder_req_address,
    output reg noc3buffer_noc3encoder_req_with_data,
    output reg noc3buffer_noc3encoder_req_was_inval,
    output reg [3:0] noc3buffer_noc3encoder_req_fwdack_vector,
    output reg [(14+8+8)-1:0] noc3buffer_noc3encoder_req_homeid,
    input wire noc3encoder_noc3buffer_req_ack,
    output reg noc3buffer_l15_req_ack
   );
reg buffer_val;
reg buffer_val_next;
reg new_buffer;
reg [3-1:0] l15_noc3encoder_req_type_buf;
reg [63:0] l15_noc3encoder_req_data_0_buf;
reg [63:0] l15_noc3encoder_req_data_1_buf;
reg [2-1:0] l15_noc3encoder_req_mshrid_buf;
reg [1:0] l15_noc3encoder_req_threadid_buf;
reg [1:0] l15_noc3encoder_req_sequenceid_buf;
reg [39:0] l15_noc3encoder_req_address_buf;
reg l15_noc3encoder_req_with_data_buf;
reg l15_noc3encoder_req_was_inval_buf;
reg [3:0] l15_noc3encoder_req_fwdack_vector_buf;
reg [(14+8+8)-1:0] l15_noc3encoder_req_homeid_buf;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        buffer_val <= 1'b0;
    end
    else
    begin
        buffer_val <= buffer_val_next;
        if (new_buffer)
        begin
            l15_noc3encoder_req_type_buf <= l15_noc3encoder_req_type;
            l15_noc3encoder_req_data_0_buf <= l15_noc3encoder_req_data_0;
            l15_noc3encoder_req_data_1_buf <= l15_noc3encoder_req_data_1;
            l15_noc3encoder_req_mshrid_buf <= l15_noc3encoder_req_mshrid;
            l15_noc3encoder_req_threadid_buf <= l15_noc3encoder_req_threadid;
            l15_noc3encoder_req_sequenceid_buf <= l15_noc3encoder_req_sequenceid;
            l15_noc3encoder_req_address_buf <= l15_noc3encoder_req_address;
            l15_noc3encoder_req_with_data_buf <= l15_noc3encoder_req_with_data;
            l15_noc3encoder_req_was_inval_buf <= l15_noc3encoder_req_was_inval;
            l15_noc3encoder_req_fwdack_vector_buf <= l15_noc3encoder_req_fwdack_vector;
            l15_noc3encoder_req_homeid_buf <= l15_noc3encoder_req_homeid;
        end
    end
end
always @ *
begin
    noc3buffer_noc3encoder_req_val = buffer_val;
    noc3buffer_noc3encoder_req_type = l15_noc3encoder_req_type_buf;
    noc3buffer_noc3encoder_req_data_0 = l15_noc3encoder_req_data_0_buf;
    noc3buffer_noc3encoder_req_data_1 = l15_noc3encoder_req_data_1_buf;
    noc3buffer_noc3encoder_req_mshrid = l15_noc3encoder_req_mshrid_buf;
    noc3buffer_noc3encoder_req_threadid = l15_noc3encoder_req_threadid_buf;
    noc3buffer_noc3encoder_req_sequenceid = l15_noc3encoder_req_sequenceid_buf;
    noc3buffer_noc3encoder_req_address = l15_noc3encoder_req_address_buf;
    noc3buffer_noc3encoder_req_with_data = l15_noc3encoder_req_with_data_buf;
    noc3buffer_noc3encoder_req_was_inval = l15_noc3encoder_req_was_inval_buf;
    noc3buffer_noc3encoder_req_fwdack_vector = l15_noc3encoder_req_fwdack_vector_buf;
    noc3buffer_noc3encoder_req_homeid = l15_noc3encoder_req_homeid_buf;
end
always @ *
begin
    noc3buffer_l15_req_ack = 1'b0;
    if (l15_noc3encoder_req_val && (!buffer_val || noc3encoder_noc3buffer_req_ack))
        noc3buffer_l15_req_ack = 1'b1;
    new_buffer = noc3buffer_l15_req_ack;
    buffer_val_next = 1'b0;
    if (noc3buffer_l15_req_ack)
        buffer_val_next = 1'b1;
    else if (noc3encoder_noc3buffer_req_ack)
        buffer_val_next = 1'b0;
    else
        buffer_val_next = buffer_val;
end
endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
 
module noc3encoder(
    input wire clk,
    input wire rst_n,
    input wire l15_noc3encoder_req_val,
    input wire [3-1:0] l15_noc3encoder_req_type,
    input wire [63:0] l15_noc3encoder_req_data_0,
    input wire [63:0] l15_noc3encoder_req_data_1,
    input wire [2-1:0] l15_noc3encoder_req_mshrid,
    input wire [0:0] l15_noc3encoder_req_threadid,
    input wire [1:0] l15_noc3encoder_req_sequenceid,
    input wire [39:0] l15_noc3encoder_req_address,
    input wire l15_noc3encoder_req_with_data,
    
    input wire l15_noc3encoder_req_was_inval,
    input wire [3:0] l15_noc3encoder_req_fwdack_vector,
    input wire [(14+8+8)-1:0] l15_noc3encoder_req_homeid,
    input wire [14-1:0] chipid,
    input wire [8-1:0] coreid_x,
    input wire [8-1:0] coreid_y,
    input wire noc3out_ready,
    output reg noc3encoder_l15_req_ack,
    output reg noc3encoder_noc3out_val,
    output reg [63:0] noc3encoder_noc3out_data
   );
reg [63:0] flit;
reg [4-1:0] flit_state;
reg [4-1:0] flit_state_next;
reg [40-1:0] address;
reg [8-1:0] dest_l2_xpos;
reg [8-1:0] dest_l2_ypos;
reg [14-1:0] dest_chipid;
reg [4-1:0] dest_fbits;
reg [8-1:0] src_l2_xpos;
reg [8-1:0] src_l2_ypos;
reg [14-1:0] src_chipid;
reg [4-1:0] src_fbits;
reg [8-1:0] msg_length;
reg [8-1:0] msg_type;
reg [8-1:0] msg_mshrid;
reg [2-1:0] msg_mesi;
reg [1-1:0] msg_last_subline;
reg [5:0] msg_options_1;
reg [15:0] msg_options_2;
reg [29:0] msg_options_3;
reg [5:0] msg_options_4;
reg [1-1:0] msg_cache_type;
reg [4-1:0] msg_subline_vector;
reg [3-1:0] msg_data_size;
reg sending;
reg is_request;
reg is_response;
reg [1:0] last_subcacheline_id;
reg [63:0] l15_noc3encoder_req_data_0_f;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        l15_noc3encoder_req_data_0_f <= 0;
        
    end
    else
    begin
        if (l15_noc3encoder_req_val && is_request && flit_state_next == 4'd3)
            l15_noc3encoder_req_data_0_f <= l15_noc3encoder_req_data_0;
        else if (l15_noc3encoder_req_val && is_request && flit_state_next == 4'd4)
            l15_noc3encoder_req_data_0_f <= l15_noc3encoder_req_data_1;
        else if (l15_noc3encoder_req_val && is_response && flit_state_next == 4'd1)
            l15_noc3encoder_req_data_0_f <= l15_noc3encoder_req_data_0;
        else if (l15_noc3encoder_req_val && is_response && flit_state_next == 4'd2)
            l15_noc3encoder_req_data_0_f <= l15_noc3encoder_req_data_1;
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        flit_state <= 0;
    end
    else
    begin
        flit_state <= flit_state_next;
    end
end
always @ *
begin
    is_request = (l15_noc3encoder_req_type == 3'd1);
    is_response = !is_request;
    last_subcacheline_id =  (l15_noc3encoder_req_fwdack_vector[3] == 1'b1) ? 2'b11 :
                            (l15_noc3encoder_req_fwdack_vector[2] == 1'b1) ? 2'b10 :
                            (l15_noc3encoder_req_fwdack_vector[1] == 1'b1) ? 2'b01 :
                                                                             2'b00 ;
    msg_last_subline = last_subcacheline_id == l15_noc3encoder_req_sequenceid;
    address = l15_noc3encoder_req_address;
    dest_l2_xpos = l15_noc3encoder_req_homeid[8-1:0];
    dest_l2_ypos = l15_noc3encoder_req_homeid[8+8-1:8];
    dest_chipid = l15_noc3encoder_req_homeid[((14+8+8)-1):(8+8)];
    dest_fbits = 4'd0;
    src_l2_xpos = coreid_x;
    src_l2_ypos = coreid_y;
    src_chipid = chipid;
    src_fbits = 4'd0;
    msg_length = 0;
    msg_type = 0;
    msg_mshrid = {l15_noc3encoder_req_threadid, l15_noc3encoder_req_mshrid};
    msg_mesi = 0;
    
    
    msg_cache_type = 0;
    msg_subline_vector = 0; 
    msg_data_size = 0;
    sending = l15_noc3encoder_req_val;
    noc3encoder_noc3out_val = sending;
    case (l15_noc3encoder_req_type)
        3'd1:
        begin
            
            msg_type = 8'd12;
            msg_length = 4; 
            
        end
        3'd3:
        begin
            msg_type = 8'd21;
            if (l15_noc3encoder_req_with_data)
            begin
                msg_length = 2;
                msg_data_size = 3'b110;
            end
            else
                msg_length = 0;
        end
        3'd2:
        begin
            
            if (l15_noc3encoder_req_was_inval)
               msg_type = 8'd23;
            else
               msg_type = 8'd22;
           
            if (l15_noc3encoder_req_with_data)
            begin
                msg_length = 2;
                msg_data_size = 3'b110;
            end
            else
                msg_length = 0;
        end
        3'd4:
        begin
            
            msg_type = 8'd23;
            msg_length = 0;
        end
    endcase
    msg_options_1 = 0;
    msg_options_2 = 0;
    msg_options_3 = 0;
    msg_options_4 = 0;
    
    msg_options_2[10:8] = msg_data_size;
    msg_options_2[11] = msg_cache_type;
    msg_options_2[15:12] = msg_subline_vector;
    msg_options_4[0] = msg_last_subline || (l15_noc3encoder_req_type == 3'd4);
    msg_options_4[2:1] = l15_noc3encoder_req_sequenceid;
    
    
    
    flit[64-1:0] = 0; 
    if (is_request)
    begin
        if (flit_state == 4'd0)
        begin
            flit[63:50] = dest_chipid;
            flit[49:42] = dest_l2_xpos;
            flit[41:34] = dest_l2_ypos;
            flit[33:30] = dest_fbits;
            flit[29:22] = msg_length;
            flit[21:14] = msg_type;
            flit[13:6] = msg_mshrid;
            flit[5:0] = msg_options_1;
        end
        else if (flit_state == 4'd1)
        begin
            flit[((16 + 40 - 1)):(16)] = address;
            flit[15:0] = msg_options_2;
        end
        else if (flit_state == 4'd2)
        begin
            flit[63:50] = src_chipid;
            flit[49:42] = src_l2_xpos;
            flit[41:34] = src_l2_ypos;
            flit[33:30] = src_fbits;
            flit[29:0] = msg_options_3;
        end
        else if (flit_state == 4'd3)
        begin
            flit[64-1:0] = l15_noc3encoder_req_data_0_f;
        end
        else if (flit_state == 4'd4)
        begin
            flit[64-1:0] = l15_noc3encoder_req_data_0_f;
        end
    end
    else if (is_response)
    begin
        if (flit_state == 4'd0)
        begin
            flit[63:50] = dest_chipid;
            flit[49:42] = dest_l2_xpos;
            flit[41:34] = dest_l2_ypos;
            flit[33:30] = dest_fbits;
            flit[29:22] = msg_length;
            flit[21:14] = msg_type;
            flit[13:6] = msg_mshrid;
            flit[5:0] = msg_options_4;
        end
        else if (flit_state == 4'd1)
        begin
            flit[64-1:0] = l15_noc3encoder_req_data_0_f;
        end
        else if (flit_state == 4'd2)
        begin
            flit[64-1:0] = l15_noc3encoder_req_data_0_f;
        end
    end
    noc3encoder_noc3out_data = flit;
    
    flit_state_next = flit_state;
    if (sending)
    begin
        if (is_request || is_response)
            if (noc3out_ready)
            begin
                if (flit_state != msg_length)
                    flit_state_next = flit_state + 1;
                else
                    flit_state_next = 4'd0;
            end
            else
                flit_state_next = flit_state;
    end
    else
        flit_state_next = 4'd0;
    
    if (l15_noc3encoder_req_val && flit_state == msg_length && noc3out_ready)
        noc3encoder_l15_req_ack = 1'b1;
    else
        noc3encoder_l15_req_ack = 1'b0;
end
endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
module pcx_buffer(
   input wire clk,
   input wire rst_n,
   
   input wire [4:0] spc_uncore_req,
   input wire spc_uncore_atomic_req,
   input wire [124-1:0] spc_uncore_data,
   input wire [33-1:0] spc_uncore_csm_data,
   
   input wire pcxdecoder_pcxbuf_ack,
   
   output reg [4:0] uncore_spc_grant,
   
   output reg [124-1:0] pcxbuf_pcxdecoder_data,
   output reg [124-1:0] pcxbuf_pcxdecoder_data_buf1,
   output reg [33-1:0] pcxbuf_pcxdecoder_csm_data,
   output reg pcxbuf_pcxdecoder_valid
   
   );
reg [124-1:0]   buffer[0:1];
reg [124-1:0]   buffer_next[0:1];
reg                    buffer_atomic[0:1];
reg                    buffer_atomic_next[0:1];
reg                    buffer_atomic_next_next;
reg [124-1:0]   buffer_csm_data[0:1];
reg [124-1:0]   buffer_csm_data_next[0:1];
reg atomic_req_second_packet_coming;
reg atomic_req_second_packet_coming_next;
reg atomic_ack_second;
reg atomic_ack_second_next;
reg buffer_val [0:1];
reg buffer_val_next [0:1];
reg read_pos;
reg write_pos;
reg read_pos_next;
reg write_pos_next;
reg write_req;
reg write_req_next;
reg read_ack;
reg is_buffer_full;
reg is_buffer_full_1back;
reg is_req_squashed;
reg [4:0] uncore_spc_grant_next;
always @ (posedge clk)
if (~rst_n)
begin
   
   
   buffer[0] <= 1'b0;
   buffer[1] <= 1'b0;
   read_pos <= 1'b0;
   write_pos <= 1'b0;
   write_req <= 1'b0;
   buffer_val[0] <= 1'b0;
   buffer_val[1] <= 1'b0;
   buffer_atomic[0] <= 1'b0;
   buffer_atomic[1] <= 1'b0;
   buffer_atomic_next_next <= 1'b0;
   atomic_req_second_packet_coming <= 1'b0;
   atomic_ack_second <= 1'b0;
   
   
   is_buffer_full_1back <= 1'b0;
   uncore_spc_grant <= 0;
end
else
begin
   
   
      
      
      buffer[0] <= buffer_next[0];
      buffer[1] <= buffer_next[1];
      buffer_csm_data[0] <= buffer_csm_data_next[0];
      buffer_csm_data[1] <= buffer_csm_data_next[1];
      read_pos <= read_pos_next;
      write_pos <= write_pos_next;
      write_req <= write_req_next;
      buffer_val[0] <= buffer_val_next[0];
      buffer_val[1] <= buffer_val_next[1];
      buffer_atomic[0] <= buffer_atomic_next[0];
      buffer_atomic[1] <= buffer_atomic_next[1];
      buffer_atomic_next_next <= spc_uncore_atomic_req && !is_req_squashed;
      atomic_req_second_packet_coming <= atomic_req_second_packet_coming_next;
      atomic_ack_second <= atomic_ack_second_next;
      
      
      is_buffer_full_1back <= is_buffer_full;
      uncore_spc_grant <= uncore_spc_grant_next;
   
end
always @ *
begin
   
   
   
   read_ack = pcxdecoder_pcxbuf_ack;
   buffer_val_next[0] = buffer_val[0];
   buffer_val_next[1] = buffer_val[1];
   buffer_next[0] = buffer[0];
   buffer_next[1] = buffer[1];
   buffer_atomic_next[0] = buffer_atomic[0];
   buffer_atomic_next[1] = buffer_atomic[1];
   buffer_csm_data_next[0] = buffer_csm_data[0];
   buffer_csm_data_next[1] = buffer_csm_data[1];
   read_pos_next = read_pos;
   write_pos_next = write_pos;
   atomic_ack_second_next = 0;
   if (write_req)
   begin
      
      buffer_next[write_pos] = spc_uncore_data;
      buffer_csm_data_next[write_pos] = spc_uncore_csm_data;
      buffer_atomic_next[write_pos] = buffer_atomic_next_next;
      buffer_val_next[write_pos] = 1'b1;
      write_pos_next = write_pos ^ 1'b1;
   end
   if (read_ack)
   begin
      if (buffer_atomic[read_pos] == 1'b1)
      begin
         read_pos_next = read_pos;
         atomic_ack_second_next = 1'b1;
         buffer_val_next[0] = 1'b0;
         buffer_val_next[1] = 1'b0;
      end
      else
      begin
         read_pos_next = read_pos^1'b1;
         buffer_val_next[read_pos] = 1'b0;
      end
   end
   
   
   is_buffer_full = (write_pos_next == read_pos) && (buffer_val[read_pos] == 1'b1) && (uncore_spc_grant[0] != 1'b1);
   
   is_req_squashed = is_buffer_full && spc_uncore_req[0];
   
   atomic_req_second_packet_coming_next = spc_uncore_atomic_req && !is_req_squashed;
   pcxbuf_pcxdecoder_data = buffer[read_pos];
   pcxbuf_pcxdecoder_data_buf1 = buffer[read_pos^1'b1];
   pcxbuf_pcxdecoder_valid = buffer_val[read_pos];
   pcxbuf_pcxdecoder_csm_data = buffer_csm_data[read_pos];
   write_req_next = (spc_uncore_req[0] && !is_req_squashed) || atomic_req_second_packet_coming;
end
always @ *
begin
   
   
      
   
   
   
   uncore_spc_grant_next = {4'b0, pcxdecoder_pcxbuf_ack|atomic_ack_second};
end
endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
module pcx_decoder(
   input wire clk,
   input wire rst_n,
   input wire [124-1:0]   pcxbuf_pcxdecoder_data,
   input wire [124-1:0]   pcxbuf_pcxdecoder_data_buf1,
   input wire [33-1:0]   pcxbuf_pcxdecoder_csm_data,
   input wire                    pcxbuf_pcxdecoder_valid,
   input wire                    l15_pcxdecoder_ack,
   input wire                    l15_pcxdecoder_header_ack,
   output reg        pcxdecoder_pcxbuf_ack,
   output reg [4:0]  pcxdecoder_l15_rqtype,
   output reg [4-1:0]  pcxdecoder_l15_amo_op,
   output reg        pcxdecoder_l15_nc,
   output reg [2:0]  pcxdecoder_l15_size,
   output reg [0:0]  pcxdecoder_l15_threadid,
   output reg        pcxdecoder_l15_prefetch,
   output reg        pcxdecoder_l15_invalidate_cacheline,
   output reg        pcxdecoder_l15_blockstore,
   output reg        pcxdecoder_l15_blockinitstore,
   output reg [1:0]  pcxdecoder_l15_l1rplway,
   output reg        pcxdecoder_l15_val,
   output reg [39:0] pcxdecoder_l15_address,
   output reg [63:0] pcxdecoder_l15_data,
   output reg [63:0] pcxdecoder_l15_data_next_entry,
   output reg [33-1:0] pcxdecoder_l15_csm_data
   );
wire [124-1:0] message = pcxbuf_pcxdecoder_data;
reg is_message_new;
reg is_message_new_next;
always @ (posedge clk)
begin
   if (!rst_n)
      is_message_new <= 1'b1;
   else
      is_message_new <= is_message_new_next;
end
reg [2:0] pcxdecoder_l15_size_pcx_standard;
reg [2:0] pcxdecoder_l15_size_pmesh_standard;
always @ *
begin
   pcxdecoder_l15_val = pcxbuf_pcxdecoder_valid && message[123] && is_message_new;
   
   pcxdecoder_pcxbuf_ack = l15_pcxdecoder_ack || (pcxbuf_pcxdecoder_valid && !message[123]);
   pcxdecoder_l15_csm_data = pcxbuf_pcxdecoder_csm_data;
   pcxdecoder_l15_rqtype = message[122:118];
   pcxdecoder_l15_amo_op = 4'b0000;
   pcxdecoder_l15_nc = message[117];
   pcxdecoder_l15_threadid = message[113:112];
   pcxdecoder_l15_prefetch = message[110];
   pcxdecoder_l15_blockstore = message[110];
   pcxdecoder_l15_invalidate_cacheline = message[111];
   pcxdecoder_l15_blockinitstore = message[109];
   pcxdecoder_l15_l1rplway = message[108:107];
   pcxdecoder_l15_size_pcx_standard = message[106:104];
   pcxdecoder_l15_address = message[103:64]; 
   pcxdecoder_l15_data = message[63:0];
   pcxdecoder_l15_data_next_entry = pcxbuf_pcxdecoder_data_buf1[63:0];
   
   
   
   is_message_new_next = l15_pcxdecoder_ack ? 1'b1 :
                         l15_pcxdecoder_header_ack ? 1'b0 : is_message_new;
   if (message[122:118] == 5'b00010)
   begin
      pcxdecoder_l15_rqtype = 5'b00110;
      pcxdecoder_l15_amo_op = 4'b1100;
   end
   else if (message[122:118] == 5'b00011)
   begin
      pcxdecoder_l15_rqtype = 5'b00110;
      pcxdecoder_l15_amo_op = 4'b1101;
   end
   else if (message[122:118] == 5'b00110)
   begin
      pcxdecoder_l15_rqtype = 5'b00110;
      pcxdecoder_l15_amo_op = 4'b0011;
   end
end
always @(*) begin
   case (pcxdecoder_l15_size_pcx_standard)
      3'b000:
         pcxdecoder_l15_size_pmesh_standard = 3'b001;
      3'b001:
         pcxdecoder_l15_size_pmesh_standard = 3'b010;
      3'b010:
         pcxdecoder_l15_size_pmesh_standard = 3'b011;
      3'b011:
         pcxdecoder_l15_size_pmesh_standard = 3'b100;
      3'b111:
         pcxdecoder_l15_size_pmesh_standard = 3'b101;
   endcase
    pcxdecoder_l15_size = pcxdecoder_l15_size_pmesh_standard;
end
endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
 
module pico_decoder(
    input wire         clk,
    input wire         rst_n,
    
    input wire         pico_mem_valid,
    input wire [31:0]  pico_mem_addr,
    input wire [ 3:0]  pico_mem_wstrb,
    
    input wire [31:0]  pico_mem_wdata,
    input wire [4-1:0] pico_mem_amo_op,
    input wire         l15_picodecoder_ack,
    input wire         l15_picodecoder_header_ack,
    
    
    output reg  [4:0]  picodecoder_l15_rqtype,
    output      [4-1:0] picodecoder_l15_amo_op,
    output reg  [2:0]  picodecoder_l15_size,
    output wire        picodecoder_l15_val,
    output wire [39:0] picodecoder_l15_address,
    output wire [63:0] picodecoder_l15_data,
    output wire        picodecoder_l15_nc,
    
    
    
    output wire [0:0]  picodecoder_l15_threadid,
    output wire        picodecoder_l15_prefetch,
    output wire        picodecoder_l15_invalidate_cacheline,
    output wire        picodecoder_l15_blockstore,
    output wire        picodecoder_l15_blockinitstore,
    output wire [1:0]  picodecoder_l15_l1rplway,
    output wire [63:0] picodecoder_l15_data_next_entry,
    output wire [32:0] picodecoder_l15_csm_data
);
    localparam ACK_IDLE = 1'b0;
    localparam ACK_WAIT = 1'b1;
    assign picodecoder_l15_amo_op = pico_mem_amo_op;
    reg current_val;
    reg prev_val;
    
    wire new_request = current_val & ~prev_val;
    always @ (posedge clk)
    begin
        if (!rst_n) begin
           current_val <= 0;
           prev_val <= 0;
        end
        else begin
           current_val <= pico_mem_valid;
           prev_val <= current_val;
        end
    end 
    
    reg ack_reg;
    reg ack_next;
    always @ (posedge clk) begin
        if (!rst_n) begin
            ack_reg <= 0;
        end
        else begin
            ack_reg <= ack_next;
        end
    end
    always @ (*) begin
        
        if (l15_picodecoder_ack) begin
            ack_next = ACK_IDLE;
        end
        else if (new_request) begin
            ack_next = ACK_WAIT;
        end
        else begin
            ack_next = ack_reg;
        end
    end
    
    
    
    
	assign picodecoder_l15_val = (ack_reg == ACK_WAIT) ? pico_mem_valid 
                                 : (ack_reg == ACK_IDLE) ? new_request
                                 : pico_mem_valid;
    reg [31:0] pico_wdata_flipped;
    
	assign picodecoder_l15_threadid = 1'b0;
	assign picodecoder_l15_prefetch = 1'b0;
	assign picodecoder_l15_csm_data = 33'b0;
	assign picodecoder_l15_data_next_entry = 64'b0;
	assign picodecoder_l15_blockstore = 1'b0;
	assign picodecoder_l15_blockinitstore = 1'b0;
	
	assign picodecoder_l15_l1rplway = 2'b0;
	
	assign picodecoder_l15_invalidate_cacheline = 1'b0;
    
	assign picodecoder_l15_address = {{8{pico_mem_addr[31]}}, pico_mem_addr};
   	assign picodecoder_l15_nc = pico_mem_addr[31] | (picodecoder_l15_rqtype == 5'b00110);
    assign picodecoder_l15_data = {pico_wdata_flipped, pico_wdata_flipped};
	
	always @ *
	begin
        if (pico_mem_valid) begin
	        
            if (pico_mem_wstrb) begin
	            picodecoder_l15_rqtype = 5'b00001;
                
                pico_wdata_flipped = {pico_mem_wdata[7:0], pico_mem_wdata[15:8],
                                      pico_mem_wdata[23:16], pico_mem_wdata[31:24]};
                
                
                if (pico_mem_amo_op != 4'b0000) begin
                    picodecoder_l15_rqtype = 5'b00110;
                end
                case(pico_mem_wstrb)
		            4'b1111: begin
		                picodecoder_l15_size = 3'b011;
		            end
		            4'b1100, 4'b0011: begin
		                picodecoder_l15_size = 3'b010;
		            end
		            4'b1000, 4'b0100, 4'b0010, 4'b0001: begin
		                picodecoder_l15_size = 3'b001;
		            end
		            
		            default: begin
		                picodecoder_l15_size = 0;
		            end
	            endcase
	        end
	        
	        else begin
	            pico_wdata_flipped = 32'b0;
                picodecoder_l15_rqtype = 5'b00000;
	            picodecoder_l15_size = 3'b011;
	        end 
        end
        else begin
            pico_wdata_flipped = 32'b0;
            picodecoder_l15_rqtype = 5'b0;
            picodecoder_l15_size = 3'b0;
        end
    end
endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
module simplenocbuffer(
   input wire clk,
   input wire rst_n,
   input wire noc_in_val,
   input wire [64-1:0] noc_in_data,
   input wire msg_ack,
   output reg noc_in_rdy,
   output reg [511:0] msg,
   output reg msg_val
   );
reg [2:0] index;
reg [2:0] index_next;
reg [8-1:0] msg_len;
reg [2-1:0] state;
reg [2-1:0] state_next;
reg [64-1:0] buffer [0:7];
reg [64-1:0] buffer_next [0:7];
always @ (posedge clk)
begin
   if (~rst_n)
   begin
      buffer[0] <= 1'b0;
      buffer[1] <= 1'b0;
      buffer[2] <= 1'b0;
      buffer[3] <= 1'b0;
      buffer[4] <= 1'b0;
      buffer[5] <= 1'b0;
      buffer[6] <= 1'b0;
      buffer[7] <= 1'b0;
      index <= 0;
      state <= 0;
   end
   else
   begin
      buffer[0] <= buffer_next[0];
      buffer[1] <= buffer_next[1];
      buffer[2] <= buffer_next[2];
      buffer[3] <= buffer_next[3];
      buffer[4] <= buffer_next[4];
      buffer[5] <= buffer_next[5];
      buffer[6] <= buffer_next[6];
      buffer[7] <= buffer_next[7];
      index <= index_next;
      state <= state_next;
   end
end
always @ *
begin
   msg[(0+1)*64 - 1 -: 64] = buffer[0];
   msg[(1+1)*64 - 1 -: 64] = buffer[1];
   msg[(2+1)*64 - 1 -: 64] = buffer[2];
   msg[(3+1)*64 - 1 -: 64] = buffer[3];
   msg[(4+1)*64 - 1 -: 64] = buffer[4];
   msg[(5+1)*64 - 1 -: 64] = buffer[5];
   msg[(6+1)*64 - 1 -: 64] = buffer[6];
   msg[(7+1)*64 - 1 -: 64] = buffer[7];
end
always @ *
begin
   index_next = index;
   state_next = 0;
   msg_val = 0;
   msg_len = 0;
   buffer_next[0] = buffer[0];
   buffer_next[1] = buffer[1];
   buffer_next[2] = buffer[2];
   buffer_next[3] = buffer[3];
   buffer_next[4] = buffer[4];
   buffer_next[5] = buffer[5];
   buffer_next[6] = buffer[6];
   buffer_next[7] = buffer[7];
   noc_in_rdy = 1'b0;
   if (state == 2'd0)
   begin
      noc_in_rdy = 1'b1;
      msg_len = noc_in_data[29:22];
      if (noc_in_val)
      begin
         buffer_next[0] = noc_in_data;
         if (msg_len == 0)
         begin
            state_next = 2'd2;
         end
         else
         begin
            state_next = 2'd1;
            index_next = index + 1;
         end
      end
   end
   else if (state == 2'd1)
   begin
      noc_in_rdy = 1'b1;
      msg_len = buffer[0][29:22];
      if (noc_in_val)
      begin
         buffer_next[index] = noc_in_data;
         if (index == msg_len)
         begin
            state_next = 2'd2;
         end
         else
         begin
            state_next = 2'd1;
            index_next = index + 1;
         end
      end
      else state_next = state;
   end
   else if (state == 2'd2)
   begin
      noc_in_rdy = 1'b0;
      msg_val = 1'b1;
      if (msg_ack)
      begin
         state_next = 2'd0;
         index_next = 0;
      end
      else
         state_next = 2'd2;
   end
end
endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
module l15_csm(
   input wire clk,
   input wire rst_n,
   input wire csm_en,
   
   input wire [6-1:0] system_tile_count,
   input wire [2-1:0] home_alloc_method, 
   input wire [22-1:0] l15_hmt_base_reg,
   
   input wire [3-1:0] l15_csm_read_ticket,
   input wire [3-1:0] l15_csm_clear_ticket,
   input wire l15_csm_clear_ticket_val,
   output wire [(14+8+8)-1:0] csm_l15_read_res_data,
   output wire csm_l15_read_res_val,
   
   input wire [40-1:0] l15_csm_req_address_s2,
   input wire l15_csm_req_val_s2,
   input wire l15_csm_stall_s3,
   input wire [3-1:0] l15_csm_req_ticket_s2,
   input wire  l15_csm_req_type_s2,     
   input wire [128-1:0] l15_csm_req_data_s2,
   input wire [33-1:0] l15_csm_req_pcx_data_s2, 
   output reg csm_l15_res_val_s3,
   output reg [63:0] csm_l15_res_data_s3,
   
   input wire noc1encoder_csm_req_ack,
   output wire csm_noc1encoder_req_val,
   output wire [5-1:0] csm_noc1encoder_req_type,
   output wire [3-1:0] csm_noc1encoder_req_mshrid,
   output wire [40-1:0] csm_noc1encoder_req_address,
   output wire csm_noc1encoder_req_non_cacheable,
   output wire  [3-1:0] csm_noc1encoder_req_size
);
reg [(14+8+8)-1:0] ghid_ticketed_cache [8-1:0];
reg [16-1:0] ghid_ticketed_cache_addr [8-1:0];
reg [8-1:0] ghid_ticketed_cache_val;
reg [3-1:0] write_index_s2;
reg write_val_s2;
reg [3-1:0] read_index_s2;
reg read_val_s2;
reg [6-1:0] num_homes_s2;
wire [6-1:0] lhid_s2;
reg [(14+8+8)-1:0] ghid_s2;
reg ghid_val_s2;
reg diag_en_s2;
reg flush_en_s2;
reg rd_en_s2;
reg wr_en_s2;
reg [8-1:0] addr_type_s2;
reg [16-1:0] addr_in_s2;
reg [16-1:0] addr_in_s2_next;
reg [6-1:0] home_addr_bits_s2;
reg special_l2_addr_s2;
reg [6-1:0] l15_csm_clump_tile_count_s2;
reg [10-1:0] l15_csm_req_clump_id_s2;
reg [14-1:0] l15_csm_chipid_s2;
reg [8-1:0] l15_csm_x_s2;
reg [8-1:0] l15_csm_y_s2;
reg l15_csm_clump_sel_s2;
always @ *
begin
    l15_csm_clump_sel_s2 = l15_csm_req_pcx_data_s2[32];
end
always @ *
begin
    if (l15_csm_clump_sel_s2 == 1'b0)
    begin
        l15_csm_clump_tile_count_s2 = l15_csm_req_pcx_data_s2[21:16];
        l15_csm_req_clump_id_s2 =  l15_csm_req_pcx_data_s2[31:22];
    end
    else
    begin
        l15_csm_clump_tile_count_s2 = 0;
        l15_csm_req_clump_id_s2 =  0;
    end
end
always @ *
begin
    if (l15_csm_clump_sel_s2 == 1'b1)
    begin
        l15_csm_chipid_s2 = l15_csm_req_pcx_data_s2[29:16];
        l15_csm_x_s2 =  l15_csm_req_pcx_data_s2[7:0];
        l15_csm_y_s2 =  l15_csm_req_pcx_data_s2[15:8];
    end
    else
    begin
        l15_csm_chipid_s2 = 0;
        l15_csm_x_s2 =  0;
        l15_csm_y_s2 =  0;
    end
end
always @ *
begin
    addr_type_s2 = l15_csm_req_address_s2[39:32];
end
always @ *
begin
    
    special_l2_addr_s2 = (l15_csm_req_address_s2[39:36] == 4'b1010);
end
always @ *
begin
    if (special_l2_addr_s2)
    begin
        home_addr_bits_s2 = l15_csm_req_address_s2[6+23 : 24];
    end
    else
    begin
        case (home_alloc_method)
        2'd0:
        begin
            home_addr_bits_s2 = l15_csm_req_address_s2[6+5 : 6];
        end
        2'd1:
        begin
            home_addr_bits_s2 = l15_csm_req_address_s2[6+13 : 14];
        end
        2'd2:
        begin
            home_addr_bits_s2 = l15_csm_req_address_s2[6+23 : 24];
        end
        2'd3:
        begin
            home_addr_bits_s2 = (l15_csm_req_address_s2[6+5 : 6] ^ l15_csm_req_address_s2[6+13 : 14]);
        end
        endcase
    end
end
always @ *
begin
    diag_en_s2 = l15_csm_req_val_s2 && (addr_type_s2 == 8'hb2);
    flush_en_s2 = l15_csm_req_val_s2 && (addr_type_s2 == 8'hb5);
    rd_en_s2 = l15_csm_req_val_s2 && (l15_csm_req_type_s2 == 1'b0)
            && ~(~diag_en_s2 && ~flush_en_s2 && (l15_csm_clump_sel_s2 == 1'b1));
    wr_en_s2 = l15_csm_req_val_s2 && (l15_csm_req_type_s2 == 1'b1);
end
always @ *
begin
   if(diag_en_s2 || flush_en_s2)
   begin
      addr_in_s2 = l15_csm_req_address_s2[16+3:4];
   end
   else
   begin
      addr_in_s2 = {l15_csm_req_clump_id_s2, lhid_s2};
   end
end
always @ *
begin
   if (csm_en)
   begin
      num_homes_s2 = l15_csm_clump_tile_count_s2;
   end
   else
   begin
      num_homes_s2 = system_tile_count;
   end
end
l15_home_encoder    l15_home_encoder(
   
   
   .home_in        (home_addr_bits_s2),
   .num_homes      (num_homes_s2),
   .lhid_out       (lhid_s2)
);
always @ *
begin
   
   
   write_index_s2 = l15_csm_req_ticket_s2;
   write_val_s2 = l15_csm_req_val_s2 && wr_en_s2 && (~diag_en_s2) && (~flush_en_s2);
end
always @ *
begin
   read_index_s2 = l15_csm_req_ticket_s2;
   read_val_s2 = l15_csm_req_val_s2 && (l15_csm_req_type_s2 == 1'b0);
end
always @ *
begin  
    case(ghid_ticketed_cache_addr[write_index_s2][1:0])
    2'd0:
    begin
        ghid_s2 = l15_csm_req_data_s2;
        ghid_val_s2 = l15_csm_req_data_s2 >> ((128/4) - 1);
    end
    2'd1:
    begin
        ghid_s2 = l15_csm_req_data_s2 >> (128/4);
        ghid_val_s2 = l15_csm_req_data_s2 >> ((128/4) * 2 - 1);
    end
    2'd2:
    begin
        ghid_s2 = l15_csm_req_data_s2 >> ((128/4) * 2);
        ghid_val_s2 = l15_csm_req_data_s2 >> ((128/4) * 3 - 1);
    end
    2'd3:
    begin
        ghid_s2 = l15_csm_req_data_s2 >> ((128/4) * 3);
        ghid_val_s2 = l15_csm_req_data_s2 >> ((128/4) * 4 - 1);
    end
    endcase
end
always @ (posedge clk)
begin
   if (!rst_n)
   begin
      ghid_ticketed_cache_val[0] <= 0;
ghid_ticketed_cache[0] <= 0;
ghid_ticketed_cache_val[1] <= 0;
ghid_ticketed_cache[1] <= 0;
ghid_ticketed_cache_val[2] <= 0;
ghid_ticketed_cache[2] <= 0;
ghid_ticketed_cache_val[3] <= 0;
ghid_ticketed_cache[3] <= 0;
ghid_ticketed_cache_val[4] <= 0;
ghid_ticketed_cache[4] <= 0;
ghid_ticketed_cache_val[5] <= 0;
ghid_ticketed_cache[5] <= 0;
ghid_ticketed_cache_val[6] <= 0;
ghid_ticketed_cache[6] <= 0;
ghid_ticketed_cache_val[7] <= 0;
ghid_ticketed_cache[7] <= 0;
   end
   else
   begin
      if (write_val_s2)
      begin
         ghid_ticketed_cache[write_index_s2] <= ghid_s2;
         ghid_ticketed_cache_val[write_index_s2] <= ghid_val_s2;
         if (l15_csm_clear_ticket_val && (l15_csm_clear_ticket != write_index_s2))
         begin
            ghid_ticketed_cache_val[l15_csm_clear_ticket] <= 1'b0;
         end
      end
      else if (read_val_s2)
      begin
         ghid_ticketed_cache[read_index_s2] <= 0;
         ghid_ticketed_cache_val[read_index_s2] <=1'b0;
         if (l15_csm_clear_ticket_val && (l15_csm_clear_ticket != read_index_s2))
         begin
            ghid_ticketed_cache_val[l15_csm_clear_ticket] <= 1'b0;
         end
      end
      else if (l15_csm_clear_ticket_val)
      begin
          ghid_ticketed_cache_val[l15_csm_clear_ticket] <= 1'b0;
      end
   end
end
always @ *
begin
    if (write_val_s2)
    begin
        addr_in_s2_next = ghid_ticketed_cache_addr[write_index_s2];
    end
    else
    begin
        addr_in_s2_next = addr_in_s2;
    end
end
reg [40-1:0] l15_csm_req_address_s3;
reg [10-1:0] l15_csm_req_clump_id_s3;
reg l15_csm_req_val_s3;
reg [3-1:0] l15_csm_req_ticket_s3;
reg [16-1:0] addr_in_s3;
reg [128-1:0] data_in_s3;
reg [6-1:0] lhid_s3;
reg diag_en_s3;
reg flush_en_s3;
reg rd_en_s3;
reg wr_en_s3;
reg [14-1:0] l15_csm_chipid_s3;
reg [8-1:0] l15_csm_x_s3;
reg [8-1:0] l15_csm_y_s3;
reg l15_csm_clump_sel_s3;
always @ (posedge clk)
begin
   if (!rst_n)
   begin
      l15_csm_req_address_s3 <= 0;
      l15_csm_req_clump_id_s3 <= 0;
      l15_csm_req_val_s3 <= 0;
      l15_csm_req_ticket_s3 <= 0;
      addr_in_s3 <= 0;
      data_in_s3 <= 0;
      lhid_s3 <= 0;
      diag_en_s3 <= 0;
      flush_en_s3 <= 0;
      rd_en_s3 <= 0;
      wr_en_s3 <= 0;
      l15_csm_chipid_s3 <= 0;
      l15_csm_x_s3 <= 0;
      l15_csm_y_s3 <= 0;
      l15_csm_clump_sel_s3 <= 0;
   end
   else
   begin
      if (!l15_csm_stall_s3)
      begin
         l15_csm_req_address_s3 <= l15_csm_req_address_s2;
         l15_csm_req_clump_id_s3 <= l15_csm_req_clump_id_s2;
         l15_csm_req_val_s3 <= l15_csm_req_val_s2;
         l15_csm_req_ticket_s3 <= l15_csm_req_ticket_s2;
         addr_in_s3 <= addr_in_s2_next;
         data_in_s3 <= l15_csm_req_data_s2;
         lhid_s3 <= lhid_s2;
         diag_en_s3 <= diag_en_s2;
         flush_en_s3 <= flush_en_s2;
         rd_en_s3 <= rd_en_s2;
         wr_en_s3 <= wr_en_s2;
         l15_csm_chipid_s3 <= l15_csm_chipid_s2;
         l15_csm_x_s3 <= l15_csm_x_s2;
         l15_csm_y_s3 <= l15_csm_y_s2;
         l15_csm_clump_sel_s3 <= l15_csm_clump_sel_s2;
      end
   end
end
reg [2-1:0] addr_op_s3;
reg refill_req_val_s3;
wire hit_s3;
wire [30-1:0] data_out_s3;
wire [4-1:0] valid_out_s3;
wire [14-1:0] tag_out_s3;
wire [8-1:0] lhid_s3_x;
wire [8-1:0] lhid_s3_y;
always @ *
begin
    addr_op_s3 = l15_csm_req_address_s3[31:30];
end
l15_hmc l15_hmc(
   .clk            (clk),
   .rst_n          (rst_n),
   .rd_en          (rd_en_s3),
   .wr_en          (wr_en_s3),
   .rd_diag_en     (diag_en_s3),
   .wr_diag_en     (diag_en_s3),
   .flush_en       (flush_en_s3),
   .addr_op        (addr_op_s3),
   .rd_addr_in     (addr_in_s3),
   .wr_addr_in     (addr_in_s3),
   .data_in        (data_in_s3),
   .hit            (hit_s3),
   .data_out       (data_out_s3),
   .valid_out      (valid_out_s3),
   .tag_out        (tag_out_s3)
);
always @ *
begin
    refill_req_val_s3 = csm_en && rd_en_s3 && (~diag_en_s3) && (~flush_en_s3) && (~hit_s3);
end
always @ *
begin
    if (csm_en)
    begin
        csm_l15_res_val_s3 = rd_en_s3 && ~refill_req_val_s3;
    end
    else
    begin
        csm_l15_res_val_s3 = l15_csm_req_val_s3;
    end
end
always @ *
begin
    if (diag_en_s3)
    begin
        if (addr_op_s3 == 0)
        begin
            csm_l15_res_data_s3 = data_out_s3;
        end
        else if (addr_op_s3 == 1)
        begin
            csm_l15_res_data_s3 = valid_out_s3;
        end
        else if (addr_op_s3 == 2)
        begin
            csm_l15_res_data_s3 = tag_out_s3;
        end
        else
        begin
            csm_l15_res_data_s3 = 0;
        end
    end
    else
    begin
        if (csm_en)
        begin
            if (~diag_en_s3 && ~flush_en_s3 && (l15_csm_clump_sel_s3 == 1'b1))
            begin
                csm_l15_res_data_s3 = 0;
                csm_l15_res_data_s3[((14+8+8)-1):(8+8)] = l15_csm_chipid_s3;
                
                csm_l15_res_data_s3[8-1:0] = l15_csm_y_s3;
                csm_l15_res_data_s3[8+8-1:8] = l15_csm_x_s3;
            end
            else
            begin
                csm_l15_res_data_s3 = data_out_s3;
            end
        end
        else
        begin
            csm_l15_res_data_s3 = 0;
            csm_l15_res_data_s3[((14+8+8)-1):(8+8)] = 1'b0; 
            csm_l15_res_data_s3[8+8-1:8] = lhid_s3_y;
            csm_l15_res_data_s3[8-1:0] = lhid_s3_x;
        end
    end
end
flat_id_to_xy lhid_to_xy (
    .flat_id(lhid_s3[6-1:0]),
    .x_coord(lhid_s3_x),
    .y_coord(lhid_s3_y)
    );
always @ (posedge clk)
begin
   if (!rst_n)
   begin
      ghid_ticketed_cache_addr[0] <= 0;
ghid_ticketed_cache_addr[1] <= 0;
ghid_ticketed_cache_addr[2] <= 0;
ghid_ticketed_cache_addr[3] <= 0;
ghid_ticketed_cache_addr[4] <= 0;
ghid_ticketed_cache_addr[5] <= 0;
ghid_ticketed_cache_addr[6] <= 0;
ghid_ticketed_cache_addr[7] <= 0;
   end
   else
   begin
      if (refill_req_val_s3)
      begin
         ghid_ticketed_cache_addr[l15_csm_req_ticket_s3] <= addr_in_s3;
      end
   end
end
assign csm_l15_read_res_data = ghid_ticketed_cache[l15_csm_read_ticket];
assign csm_l15_read_res_val = ghid_ticketed_cache_val[l15_csm_read_ticket];
reg [40-1:0] refill_req_addr_buf [8-1:0];
reg [3-1:0] refill_req_ticket_buf [8-1:0];
reg [8-1:0] refill_req_val_buf;
reg [3-1:0] refill_req_buf_rd_ptr;
reg [3-1:0] refill_req_buf_rd_ptr_next;
reg [3-1:0] refill_req_buf_wr_ptr;
reg [3-1:0] refill_req_buf_wr_ptr_next;
reg [3:0] refill_req_buf_counter;
reg [3:0] refill_req_buf_counter_next;
always @ *
begin
    if (!rst_n)
    begin
        refill_req_buf_counter_next = 0;
    end
    else if (refill_req_val_s3 && noc1encoder_csm_req_ack)
    begin
        refill_req_buf_counter_next = refill_req_buf_counter;
    end
    else if (refill_req_val_s3)
    begin
        refill_req_buf_counter_next = refill_req_buf_counter + 1;
    end
    else if (noc1encoder_csm_req_ack)
    begin
        refill_req_buf_counter_next = refill_req_buf_counter - 1;
    end
    else
    begin
        refill_req_buf_counter_next = refill_req_buf_counter;
    end
end
always @ (posedge clk)
begin
    refill_req_buf_counter <= refill_req_buf_counter_next;
end
always @ *
begin
    if (!rst_n)
    begin
        refill_req_buf_rd_ptr_next = 0;
    end
    else if (noc1encoder_csm_req_ack)
    begin
        refill_req_buf_rd_ptr_next = refill_req_buf_rd_ptr + 1;
    end
    else
    begin
        refill_req_buf_rd_ptr_next = refill_req_buf_rd_ptr;
    end
end
always @ (posedge clk)
begin
    refill_req_buf_rd_ptr <= refill_req_buf_rd_ptr_next;
end
always @ *
begin
    if (!rst_n)
    begin
        refill_req_buf_wr_ptr_next = 0;
    end
    else if (refill_req_val_s3)
    begin
        refill_req_buf_wr_ptr_next = refill_req_buf_wr_ptr + 1;
    end
    else
    begin
        refill_req_buf_wr_ptr_next = refill_req_buf_wr_ptr;
    end
end
always @ (posedge clk)
begin
    refill_req_buf_wr_ptr <= refill_req_buf_wr_ptr_next;
end
always @ (posedge clk)
begin
   if (!rst_n)
   begin
      refill_req_addr_buf[0] <= 0;
refill_req_ticket_buf[0] <= 0;
refill_req_val_buf[0] <= 0;
refill_req_addr_buf[1] <= 0;
refill_req_ticket_buf[1] <= 0;
refill_req_val_buf[1] <= 0;
refill_req_addr_buf[2] <= 0;
refill_req_ticket_buf[2] <= 0;
refill_req_val_buf[2] <= 0;
refill_req_addr_buf[3] <= 0;
refill_req_ticket_buf[3] <= 0;
refill_req_val_buf[3] <= 0;
refill_req_addr_buf[4] <= 0;
refill_req_ticket_buf[4] <= 0;
refill_req_val_buf[4] <= 0;
refill_req_addr_buf[5] <= 0;
refill_req_ticket_buf[5] <= 0;
refill_req_val_buf[5] <= 0;
refill_req_addr_buf[6] <= 0;
refill_req_ticket_buf[6] <= 0;
refill_req_val_buf[6] <= 0;
refill_req_addr_buf[7] <= 0;
refill_req_ticket_buf[7] <= 0;
refill_req_val_buf[7] <= 0;
   end
   else
   begin
      if (refill_req_val_s3)
      begin
        refill_req_addr_buf[refill_req_buf_wr_ptr] <= {l15_hmt_base_reg, addr_in_s3[15:2], 4'd0};
        refill_req_ticket_buf[refill_req_buf_wr_ptr] <= l15_csm_req_ticket_s3;
        refill_req_val_buf[refill_req_buf_wr_ptr] <= refill_req_val_s3;
      end
   end
end
assign csm_noc1encoder_req_val = refill_req_val_buf[refill_req_buf_rd_ptr] && (refill_req_buf_counter > 0);
assign csm_noc1encoder_req_type = 5'd2;
assign csm_noc1encoder_req_mshrid = refill_req_ticket_buf[refill_req_buf_rd_ptr];
assign csm_noc1encoder_req_address = refill_req_addr_buf[refill_req_buf_rd_ptr];
assign csm_noc1encoder_req_non_cacheable = 1'b1;
assign csm_noc1encoder_req_size = 3'b101; 
endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
module l15_hmc(
    input wire clk,
    input wire rst_n,
    
    input wire rd_en,
    
    input wire wr_en,
    
    input wire rd_diag_en,
    
    input wire wr_diag_en,
    
    input wire flush_en,
    input wire [2-1:0] addr_op,
    
    input wire [16-1:0] rd_addr_in,
    input wire [16-1:0] wr_addr_in,
    
    input wire [128-1:0] data_in,
    output reg hit,
    
    output reg [30-1:0] data_out,
    output reg [4-1:0] valid_out,
    output reg [14-1:0] tag_out
);
reg [16-1:0] entry_used_f;
reg [16-1:0] entry_used_next;
reg [16-1:0] entry_used_and_mask;
reg [16-1:0] entry_used_or_mask;
reg [16-1:0] entry_locked_f;
reg [16-1:0] entry_locked_next;
reg [16-1:0] entry_locked_and_mask;
reg [16-1:0] entry_locked_or_mask;
reg [138-1:0] data_mem_f [16-1:0];
reg [14-1:0] smc_tag [16-1:0];
reg [4-1:0] smc_valid [16-1:0];
reg [120-1:0] smc_data [16-1:0];
reg [10-1:0] smc_sdid [16-1:0];
reg [14-1:0] rd_tag_in;
reg [14-1:0] wr_tag_in;
reg [4-1:0] rd_index_in;
reg [4-1:0] wr_index_in;
reg [2-1:0] rd_offset_in;
reg [2-1:0] wr_offset_in;
reg [10-1:0] wr_sdid_in;
reg [4-1:0] smc_valid_in;
reg [120-1:0] smc_data_in;
reg [4-1:0] hit_index;
reg [4-1:0] replace_index;
reg wr_hit;
reg [4-1:0] wr_hit_index;
reg [4-1:0] wr_index;
always @ *
begin
    smc_tag[0] = data_mem_f[0][137:124];
    smc_tag[1] = data_mem_f[1][137:124];
    smc_tag[2] = data_mem_f[2][137:124];
    smc_tag[3] = data_mem_f[3][137:124];
    smc_tag[4] = data_mem_f[4][137:124];
    smc_tag[5] = data_mem_f[5][137:124];
    smc_tag[6] = data_mem_f[6][137:124];
    smc_tag[7] = data_mem_f[7][137:124];
    smc_tag[8] = data_mem_f[8][137:124];
    smc_tag[9] = data_mem_f[9][137:124];
    smc_tag[10] = data_mem_f[10][137:124];
    smc_tag[11] = data_mem_f[11][137:124];
    smc_tag[12] = data_mem_f[12][137:124];
    smc_tag[13] = data_mem_f[13][137:124];
    smc_tag[14] = data_mem_f[14][137:124];
    smc_tag[15] = data_mem_f[15][137:124];
end
always @ *
begin
    smc_valid[0] = data_mem_f[0][123:120];
    smc_valid[1] = data_mem_f[1][123:120];
    smc_valid[2] = data_mem_f[2][123:120];
    smc_valid[3] = data_mem_f[3][123:120];
    smc_valid[4] = data_mem_f[4][123:120];
    smc_valid[5] = data_mem_f[5][123:120];
    smc_valid[6] = data_mem_f[6][123:120];
    smc_valid[7] = data_mem_f[7][123:120];
    smc_valid[8] = data_mem_f[8][123:120];
    smc_valid[9] = data_mem_f[9][123:120];
    smc_valid[10] = data_mem_f[10][123:120];
    smc_valid[11] = data_mem_f[11][123:120];
    smc_valid[12] = data_mem_f[12][123:120];
    smc_valid[13] = data_mem_f[13][123:120];
    smc_valid[14] = data_mem_f[14][123:120];
    smc_valid[15] = data_mem_f[15][123:120];
end
always @ *
begin
    smc_data[0] = data_mem_f[0][119:0];
    smc_data[1] = data_mem_f[1][119:0];
    smc_data[2] = data_mem_f[2][119:0];
    smc_data[3] = data_mem_f[3][119:0];
    smc_data[4] = data_mem_f[4][119:0];
    smc_data[5] = data_mem_f[5][119:0];
    smc_data[6] = data_mem_f[6][119:0];
    smc_data[7] = data_mem_f[7][119:0];
    smc_data[8] = data_mem_f[8][119:0];
    smc_data[9] = data_mem_f[9][119:0];
    smc_data[10] = data_mem_f[10][119:0];
    smc_data[11] = data_mem_f[11][119:0];
    smc_data[12] = data_mem_f[12][119:0];
    smc_data[13] = data_mem_f[13][119:0];
    smc_data[14] = data_mem_f[14][119:0];
    smc_data[15] = data_mem_f[15][119:0];
end
always @ *
begin
    smc_sdid[0] = data_mem_f[0][137:128];
    smc_sdid[1] = data_mem_f[1][137:128];
    smc_sdid[2] = data_mem_f[2][137:128];
    smc_sdid[3] = data_mem_f[3][137:128];
    smc_sdid[4] = data_mem_f[4][137:128];
    smc_sdid[5] = data_mem_f[5][137:128];
    smc_sdid[6] = data_mem_f[6][137:128];
    smc_sdid[7] = data_mem_f[7][137:128];
    smc_sdid[8] = data_mem_f[8][137:128];
    smc_sdid[9] = data_mem_f[9][137:128];
    smc_sdid[10] = data_mem_f[10][137:128];
    smc_sdid[11] = data_mem_f[11][137:128];
    smc_sdid[12] = data_mem_f[12][137:128];
    smc_sdid[13] = data_mem_f[13][137:128];
    smc_sdid[14] = data_mem_f[14][137:128];
    smc_sdid[15] = data_mem_f[15][137:128];
end
always @ *
begin
    rd_tag_in = rd_addr_in[15:2];
    rd_offset_in = rd_addr_in[1:0];
    rd_index_in = rd_addr_in[5:2];
end
always @ *
begin
    wr_tag_in = wr_addr_in[15:2];
    wr_offset_in = wr_addr_in[1:0];
    wr_index_in = wr_addr_in[5:2];
    wr_sdid_in = wr_addr_in[15:6];
end
always @ *
begin
    smc_valid_in = { data_in[127], data_in[95], data_in[63], data_in[31] };
    smc_data_in = { data_in[125:96], data_in[93:64], data_in[61:32], data_in[29:0] };
end
wire [4-1:0] tag_hit_index;
wire tag_hit;
reg [15:0] smc_tag_cmp;
always @ *
begin
    smc_tag_cmp[0] = (smc_tag[0] == rd_tag_in) && smc_valid[0][rd_offset_in];
    smc_tag_cmp[1] = (smc_tag[1] == rd_tag_in) && smc_valid[1][rd_offset_in];
    smc_tag_cmp[2] = (smc_tag[2] == rd_tag_in) && smc_valid[2][rd_offset_in];
    smc_tag_cmp[3] = (smc_tag[3] == rd_tag_in) && smc_valid[3][rd_offset_in];
    smc_tag_cmp[4] = (smc_tag[4] == rd_tag_in) && smc_valid[4][rd_offset_in];
    smc_tag_cmp[5] = (smc_tag[5] == rd_tag_in) && smc_valid[5][rd_offset_in];
    smc_tag_cmp[6] = (smc_tag[6] == rd_tag_in) && smc_valid[6][rd_offset_in];
    smc_tag_cmp[7] = (smc_tag[7] == rd_tag_in) && smc_valid[7][rd_offset_in];
    smc_tag_cmp[8] = (smc_tag[8] == rd_tag_in) && smc_valid[8][rd_offset_in];
    smc_tag_cmp[9] = (smc_tag[9] == rd_tag_in) && smc_valid[9][rd_offset_in];
    smc_tag_cmp[10] = (smc_tag[10] == rd_tag_in) && smc_valid[10][rd_offset_in];
    smc_tag_cmp[11] = (smc_tag[11] == rd_tag_in) && smc_valid[11][rd_offset_in];
    smc_tag_cmp[12] = (smc_tag[12] == rd_tag_in) && smc_valid[12][rd_offset_in];
    smc_tag_cmp[13] = (smc_tag[13] == rd_tag_in) && smc_valid[13][rd_offset_in];
    smc_tag_cmp[14] = (smc_tag[14] == rd_tag_in) && smc_valid[14][rd_offset_in];
    smc_tag_cmp[15] = (smc_tag[15] == rd_tag_in) && smc_valid[15][rd_offset_in];
end
l15_priority_encoder_4 priority_encoder_cmp_4bits( 
    .data_in        (smc_tag_cmp),
    .data_out       (tag_hit_index),
    .data_out_mask  (),
    .nonzero_out    (tag_hit)
);
always @ *
begin
    if (rd_en && rd_diag_en)
    begin
        hit = 1'b0;
        hit_index = rd_index_in;
    end
    else
    begin
        if(rd_en)
        begin
            hit = tag_hit;
            hit_index = tag_hit_index;
        end
        else
        begin
            hit = 1'b0;
            hit_index = 0;
        end
    end
end
wire [4-1:0] tag_wr_hit_index;
wire tag_wr_hit;
reg [15:0] smc_tag_wr_cmp;
always @ *
begin
    smc_tag_wr_cmp[0] = (smc_tag[0] == wr_tag_in) && (smc_valid[0] != 0);
    smc_tag_wr_cmp[1] = (smc_tag[1] == wr_tag_in) && (smc_valid[1] != 0);
    smc_tag_wr_cmp[2] = (smc_tag[2] == wr_tag_in) && (smc_valid[2] != 0);
    smc_tag_wr_cmp[3] = (smc_tag[3] == wr_tag_in) && (smc_valid[3] != 0);
    smc_tag_wr_cmp[4] = (smc_tag[4] == wr_tag_in) && (smc_valid[4] != 0);
    smc_tag_wr_cmp[5] = (smc_tag[5] == wr_tag_in) && (smc_valid[5] != 0);
    smc_tag_wr_cmp[6] = (smc_tag[6] == wr_tag_in) && (smc_valid[6] != 0);
    smc_tag_wr_cmp[7] = (smc_tag[7] == wr_tag_in) && (smc_valid[7] != 0);
    smc_tag_wr_cmp[8] = (smc_tag[8] == wr_tag_in) && (smc_valid[8] != 0);
    smc_tag_wr_cmp[9] = (smc_tag[9] == wr_tag_in) && (smc_valid[9] != 0);
    smc_tag_wr_cmp[10] = (smc_tag[10] == wr_tag_in) && (smc_valid[10] != 0);
    smc_tag_wr_cmp[11] = (smc_tag[11] == wr_tag_in) && (smc_valid[11] != 0);
    smc_tag_wr_cmp[12] = (smc_tag[12] == wr_tag_in) && (smc_valid[12] != 0);
    smc_tag_wr_cmp[13] = (smc_tag[13] == wr_tag_in) && (smc_valid[13] != 0);
    smc_tag_wr_cmp[14] = (smc_tag[14] == wr_tag_in) && (smc_valid[14] != 0);
    smc_tag_wr_cmp[15] = (smc_tag[15] == wr_tag_in) && (smc_valid[15] != 0);
end
l15_priority_encoder_4 priority_encoder_wr_cmp_4bits( 
    .data_in        (smc_tag_wr_cmp),
    .data_out       (tag_wr_hit_index),
    .data_out_mask  (),
    .nonzero_out    (tag_wr_hit)
);
always @ *
begin
    if(wr_en || (flush_en && (addr_op == 2'd1)))
    begin
        wr_hit = tag_wr_hit;
        wr_hit_index = tag_wr_hit_index;
    end
    else
    begin
        wr_hit = 1'b0;
        wr_hit_index = 0;
    end
end
always @ *
begin
    data_out = smc_data[hit_index]>>(rd_offset_in * 30);
    valid_out = smc_valid[hit_index];
    tag_out = smc_tag[hit_index];
end
always @ *
begin
    entry_locked_and_mask = {16{1'b1}};
    entry_locked_or_mask = {16{1'b0}};
    if (!rst_n)
    begin
        entry_locked_and_mask = {16{1'b0}};
    end
    else if (wr_en && ~wr_diag_en)
    begin
        if(smc_valid_in)
        begin
            entry_locked_or_mask[wr_index] = 1'b1;
        end
        else
        begin
            entry_locked_and_mask[wr_index] = 1'b0;
        end
        if (rd_en && ~rd_diag_en && hit && (wr_index != hit_index) && entry_locked_f[hit_index])
        begin
            entry_locked_and_mask[hit_index] = 1'b0;
        end
    end
    else if (rd_en && ~rd_diag_en && hit && entry_locked_f[hit_index])
    begin
        entry_locked_and_mask[hit_index] = 1'b0;
    end
end
always @ *
begin
    entry_locked_next = (entry_locked_f & entry_locked_and_mask) | entry_locked_or_mask;
end
always @ (posedge clk)
begin
    entry_locked_f <= entry_locked_next;
end
always @ *
begin
    entry_used_and_mask = {16{1'b1}};
    entry_used_or_mask = {16{1'b0}};
    if (!rst_n)
    begin
        entry_used_and_mask = {16{1'b0}};
    end
    else if (wr_en && ~wr_diag_en)
    begin
        if(smc_valid_in)
        begin
            entry_used_or_mask[wr_index] = 1'b1;
        end
        else
        begin
            entry_used_and_mask[wr_index] = 1'b0;
        end
        if (rd_en && ~rd_diag_en && hit && (wr_index != hit_index))
        begin
            entry_used_or_mask[hit_index] = 1'b1;
        end
    end
    else if (rd_en && ~rd_diag_en && hit)
    begin
        entry_used_or_mask[hit_index] = 1'b1;
    end
end
always @ *
begin
    entry_used_next = (entry_used_f & entry_used_and_mask) | entry_used_or_mask;
    if (entry_used_next == {16{1'b1}})
    begin
        entry_used_next = {16{1'b0}};
    end
end
always @ (posedge clk)
begin
    entry_used_f <= entry_used_next;
end
wire [4-1:0] entry_replace_index;
wire replace_hit;
reg [15:0] replace_cmp;
always @ *
begin
    replace_cmp[0] = (~entry_used_f[0] && ~entry_locked_f[0]);
    replace_cmp[1] = (~entry_used_f[1] && ~entry_locked_f[1]);
    replace_cmp[2] = (~entry_used_f[2] && ~entry_locked_f[2]);
    replace_cmp[3] = (~entry_used_f[3] && ~entry_locked_f[3]);
    replace_cmp[4] = (~entry_used_f[4] && ~entry_locked_f[4]);
    replace_cmp[5] = (~entry_used_f[5] && ~entry_locked_f[5]);
    replace_cmp[6] = (~entry_used_f[6] && ~entry_locked_f[6]);
    replace_cmp[7] = (~entry_used_f[7] && ~entry_locked_f[7]);
    replace_cmp[8] = (~entry_used_f[8] && ~entry_locked_f[8]);
    replace_cmp[9] = (~entry_used_f[9] && ~entry_locked_f[9]);
    replace_cmp[10] = (~entry_used_f[10] && ~entry_locked_f[10]);
    replace_cmp[11] = (~entry_used_f[11] && ~entry_locked_f[11]);
    replace_cmp[12] = (~entry_used_f[12] && ~entry_locked_f[12]);
    replace_cmp[13] = (~entry_used_f[13] && ~entry_locked_f[13]);
    replace_cmp[14] = (~entry_used_f[14] && ~entry_locked_f[14]);
    replace_cmp[15] = (~entry_used_f[15] && ~entry_locked_f[15]);
end
l15_priority_encoder_4 priority_encoder_replace_cmp_4bits( 
    .data_in        (replace_cmp),
    .data_out       (entry_replace_index),
    .data_out_mask  (),
    .nonzero_out    (replace_hit)
);
always @ *
begin
    if (replace_hit)
    begin
        replace_index = entry_replace_index;
    end
    else
    begin
        replace_index = {4{1'b0}};
    end
end
always @ *
begin
    if (wr_en && wr_diag_en)
    begin
        wr_index = wr_index_in;
    end
    else if ((flush_en || wr_en) && wr_hit)
    begin
        wr_index = wr_hit_index;
    end
    else
    begin
        wr_index = replace_index;
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        data_mem_f[0] <= {138{1'b0}};
        data_mem_f[1] <= {138{1'b0}};
        data_mem_f[2] <= {138{1'b0}};
        data_mem_f[3] <= {138{1'b0}};
        data_mem_f[4] <= {138{1'b0}};
        data_mem_f[5] <= {138{1'b0}};
        data_mem_f[6] <= {138{1'b0}};
        data_mem_f[7] <= {138{1'b0}};
        data_mem_f[8] <= {138{1'b0}};
        data_mem_f[9] <= {138{1'b0}};
        data_mem_f[10] <= {138{1'b0}};
        data_mem_f[11] <= {138{1'b0}};
        data_mem_f[12] <= {138{1'b0}};
        data_mem_f[13] <= {138{1'b0}};
        data_mem_f[14] <= {138{1'b0}};
        data_mem_f[15] <= {138{1'b0}};
    end
    else if (flush_en)
    begin
        case (addr_op)
        2'd0:
        begin
            data_mem_f[0][123:120] <= {4{1'b0}};
            data_mem_f[1][123:120] <= {4{1'b0}};
            data_mem_f[2][123:120] <= {4{1'b0}};
            data_mem_f[3][123:120] <= {4{1'b0}};
            data_mem_f[4][123:120] <= {4{1'b0}};
            data_mem_f[5][123:120] <= {4{1'b0}};
            data_mem_f[6][123:120] <= {4{1'b0}};
            data_mem_f[7][123:120] <= {4{1'b0}};
            data_mem_f[8][123:120] <= {4{1'b0}};
            data_mem_f[9][123:120] <= {4{1'b0}};
            data_mem_f[10][123:120] <= {4{1'b0}};
            data_mem_f[11][123:120] <= {4{1'b0}};
            data_mem_f[12][123:120] <= {4{1'b0}};
            data_mem_f[13][123:120] <= {4{1'b0}};
            data_mem_f[14][123:120] <= {4{1'b0}};
            data_mem_f[15][123:120] <= {4{1'b0}};
        end
        2'd1:
        begin
            if (wr_hit)
            begin
                data_mem_f[wr_index][120+wr_offset_in] <= 1'b0;
            end
        end
        2'd2:
        begin
            if ((smc_sdid[0] == wr_sdid_in) && (smc_valid[0] != 0))
                data_mem_f[0][123:120] <= {4{1'b0}};
            if ((smc_sdid[1] == wr_sdid_in) && (smc_valid[1] != 0))
                data_mem_f[1][123:120] <= {4{1'b0}};
            if ((smc_sdid[2] == wr_sdid_in) && (smc_valid[2] != 0))
                data_mem_f[2][123:120] <= {4{1'b0}};
            if ((smc_sdid[3] == wr_sdid_in) && (smc_valid[3] != 0))
                data_mem_f[3][123:120] <= {4{1'b0}};
            if ((smc_sdid[4] == wr_sdid_in) && (smc_valid[4] != 0))
                data_mem_f[4][123:120] <= {4{1'b0}};
            if ((smc_sdid[5] == wr_sdid_in) && (smc_valid[5] != 0))
                data_mem_f[5][123:120] <= {4{1'b0}};
            if ((smc_sdid[6] == wr_sdid_in) && (smc_valid[6] != 0))
                data_mem_f[6][123:120] <= {4{1'b0}};
            if ((smc_sdid[7] == wr_sdid_in) && (smc_valid[7] != 0))
                data_mem_f[7][123:120] <= {4{1'b0}};
            if ((smc_sdid[8] == wr_sdid_in) && (smc_valid[8] != 0))
                data_mem_f[8][123:120] <= {4{1'b0}};
            if ((smc_sdid[9] == wr_sdid_in) && (smc_valid[9] != 0))
                data_mem_f[9][123:120] <= {4{1'b0}};
            if ((smc_sdid[10] == wr_sdid_in) && (smc_valid[10] != 0))
                data_mem_f[10][123:120] <= {4{1'b0}};
            if ((smc_sdid[11] == wr_sdid_in) && (smc_valid[11] != 0))
                data_mem_f[11][123:120] <= {4{1'b0}};
            if ((smc_sdid[12] == wr_sdid_in) && (smc_valid[12] != 0))
                data_mem_f[12][123:120] <= {4{1'b0}};
            if ((smc_sdid[13] == wr_sdid_in) && (smc_valid[13] != 0))
                data_mem_f[13][123:120] <= {4{1'b0}};
            if ((smc_sdid[14] == wr_sdid_in) && (smc_valid[14] != 0))
                data_mem_f[14][123:120] <= {4{1'b0}};
            if ((smc_sdid[15] == wr_sdid_in) && (smc_valid[15] != 0))
                data_mem_f[15][123:120] <= {4{1'b0}};
        end
        default:
        begin
            data_mem_f[wr_index] <= data_mem_f[wr_index];
        end
        endcase
    end
    else if (wr_en)
    begin
        if (wr_diag_en)
        begin
            case (addr_op)
            2'd0:
            begin
                case (wr_offset_in)
                2'd0:
                begin
                    data_mem_f[wr_index][30-1:0] <=
                    data_in[30-1:0];
                end
                2'd1:
                begin
                    data_mem_f[wr_index][30*2-1:30] <=
                    data_in[30-1:0];
                end
                2'd2:
                begin
                    data_mem_f[wr_index][30*3-1:30*2] <=
                    data_in[30-1:0];
                end
                2'd3:
                begin
                    data_mem_f[wr_index][30*4-1:30*3] <=
                    data_in[30-1:0];
                end
                default:
                begin
                    data_mem_f[wr_index] <= data_mem_f[wr_index];
                end
                endcase
            end
            2'd1:
            begin
                data_mem_f[wr_index][123:120] <= data_in[4-1:0];
            end
            2'd2:
            begin
                data_mem_f[wr_index][137:124] <= data_in[14-1:0];
            end
            default:
            begin
                data_mem_f[wr_index] <= data_mem_f[wr_index];
            end
            endcase
        end
        else
        begin
            data_mem_f[wr_index] <= {wr_tag_in, smc_valid_in, smc_data_in};
        end
    end
end
endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
module l15_home_encoder(
    
    
    input wire [6-1:0] home_in,
    
    input wire [6-1:0] num_homes,
    output reg [6-1:0] lhid_out
);
reg [6-1:0] home_mask;
reg [6-1:0] home_low_mask;
reg [6-1:0] home_mod;
reg isPowerOf2;
always @ *
begin
    if (num_homes[5])
    begin
        home_low_mask = 6'b011111;
        isPowerOf2 = ~(|(num_homes[4:0]));
    end
    else if (num_homes[4])
    begin
        home_low_mask = 6'b001111;
        isPowerOf2 = ~(|(num_homes[3:0]));
    end
    else if (num_homes[3])
    begin
        home_low_mask = 6'b000111;
        isPowerOf2 = ~(|(num_homes[2:0]));
    end
    else if (num_homes[2])
    begin
        home_low_mask = 6'b000011;
        isPowerOf2 = ~(|(num_homes[1:0]));
    end
    else if (num_homes[1])
    begin
        home_low_mask = 6'b000001;
        isPowerOf2 = ~(|(num_homes[0:0]));
    end
    else if (num_homes[0])
    begin
        home_low_mask = 6'b000000;
        isPowerOf2 = 1'b1;
    end
    else
    begin
        home_low_mask = 6'b111111;
        isPowerOf2 = 1'b1;
    end
end
always @ *
begin
    if (isPowerOf2) 
    begin
        home_mask = home_low_mask;
    end
    else 
    begin
        home_mask = {home_low_mask[6-2:0], 1'b1};
    end
end
always @ *
begin
    home_mod = home_in & home_mask;
end
always @ *
begin
    if (home_mod < num_homes)
    begin
        lhid_out = home_mod;
    end
    else
    begin
        lhid_out = home_mod & home_low_mask;
    end
end
endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
module l15_mshr(
    input wire clk,
    input wire rst_n,
    
    input wire pipe_mshr_writereq_val_s1,
    input wire [3-1:0] pipe_mshr_writereq_op_s1,
    input wire [39:0] pipe_mshr_writereq_address_s1,
    input wire [127:0] pipe_mshr_writereq_write_buffer_data_s1,
    input wire [15:0] pipe_mshr_writereq_write_buffer_byte_mask_s1,
    input wire [((((((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) + 1) + 1) + 1)-1:0] pipe_mshr_writereq_control_s1,
    input wire [2-1:0] pipe_mshr_writereq_mshrid_s1,
    input wire [0:0] pipe_mshr_writereq_threadid_s1,
    input wire [0:0] pipe_mshr_readreq_threadid_s1,
    input wire [2-1:0] pipe_mshr_readreq_mshrid_s1,
    output reg [((((((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) + 1) + 1) + 1)-1:0]mshr_pipe_readres_control_s1,
    output reg [(14+8+8)-1:0] mshr_pipe_readres_homeid_s1,
    
    output reg [(4*2)-1:0] mshr_pipe_vals_s1,
    output reg [(40*2)-1:0] mshr_pipe_ld_address,
    output reg [(40*2)-1:0] mshr_pipe_st_address,
    output reg [(2*2)-1:0] mshr_pipe_st_way_s1,
    output reg [(2*2)-1:0] mshr_pipe_st_state_s1,
    
    input wire pipe_mshr_write_buffer_rd_en_s2,
    input wire [0:0] pipe_mshr_threadid_s2,
    output reg [127:0]mshr_pipe_write_buffer_s2,
    output reg [15:0] mshr_pipe_write_buffer_byte_mask_s2,
    
    input wire pipe_mshr_val_s3,
    input wire [3-1:0] pipe_mshr_op_s3,
    input wire [2-1:0] pipe_mshr_mshrid_s3,
    input wire [0:0] pipe_mshr_threadid_s3,
    input wire [2-1:0] pipe_mshr_write_update_state_s3,
    input wire [1:0] pipe_mshr_write_update_way_s3,
    
    
    
    
    
    input wire noc1buffer_mshr_homeid_write_val_s4,
    input wire [2-1:0] noc1buffer_mshr_homeid_write_mshrid_s4,
    input wire [0:0] noc1buffer_mshr_homeid_write_threadid_s4,
    input wire [(14+8+8)-1:0] noc1buffer_mshr_homeid_write_data_s4
    );
reg [39:0] ld_address [0:2-1];
reg [((((((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) + 1) + 1) + 1)-1:0] ld_control [0:2-1];
reg [2-1:0] ld_val;
reg [(14+8+8)-1:0] ld_homeid [0:2-1];
reg [((((((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) + 1) + 1) + 1)-1:0] ifill_control [0:2-1];
reg [2-1:0] ifill_val;
reg [39:0] st_address [0:2-1];
reg [((((((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) + 1) + 1) + 1)-1:0] st_control [0:2-1];
reg [2-1:0] st_val;
reg [(14+8+8)-1:0] st_homeid [0:2-1];
reg [2-1:0] st_state [0:2-1];
reg [1:0] st_way [0:2-1];
reg [127:0] st_write_buffer [0:2-1];
reg [15:0] st_write_buffer_byte_mask [0:2-1];
reg [3-1:0] op_s1;
reg [3-1:0] op_s3;
reg [0:0] threadid_s1;
reg [0:0] threadid_s3;
reg [2-1:0] mshrid_s1;
reg [2-1:0] mshrid_s3;
always @ *
begin
    op_s1 = pipe_mshr_writereq_op_s1;
    threadid_s1 = pipe_mshr_writereq_threadid_s1;
    mshrid_s1 = pipe_mshr_writereq_mshrid_s1;
    threadid_s3 = pipe_mshr_threadid_s3;
    op_s3 = pipe_mshr_op_s3;
    mshrid_s3 = pipe_mshr_mshrid_s3;
end
reg [4-1:0] tmp_vals [2-1:0];
reg [39:0] tmp_st_address [2-1:0];
reg [39:0] tmp_ld_address [2-1:0];
reg [2-1:0] tmp_st_way [2-1:0];
reg [2-1:0] tmp_st_state [2-1:0];
always @ *
begin
    
tmp_vals[0] = 0;
tmp_vals[0][2'd1] = ifill_val[0];
tmp_vals[0][2'd2] = ld_val[0];
tmp_vals[0][2'd3] = st_val[0];
tmp_st_address[0] = st_address[0];
tmp_ld_address[0] = ld_address[0];
tmp_st_way[0] = st_way[0];
tmp_st_state[0] =st_state[0];
tmp_vals[1] = 0;
tmp_vals[1][2'd1] = ifill_val[1];
tmp_vals[1][2'd2] = ld_val[1];
tmp_vals[1][2'd3] = st_val[1];
tmp_st_address[1] = st_address[1];
tmp_ld_address[1] = ld_address[1];
tmp_st_way[1] = st_way[1];
tmp_st_state[1] =st_state[1];
    mshr_pipe_vals_s1 = {tmp_vals[1], tmp_vals[0]};
    mshr_pipe_ld_address = {tmp_ld_address[1], tmp_ld_address[0]};
    mshr_pipe_st_address = {tmp_st_address[1], tmp_st_address[0]};
    mshr_pipe_st_way_s1 = {tmp_st_way[1], tmp_st_way[0]};
    mshr_pipe_st_state_s1 = {tmp_st_state[1], tmp_st_state[0]};
    
    mshr_pipe_readres_homeid_s1[(14+8+8)-1:0] = 0;
    mshr_pipe_readres_control_s1[((((((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) + 1) + 1) + 1)-1:0] = 0;
    case (pipe_mshr_readreq_mshrid_s1)
        2'd1:
        begin
            mshr_pipe_readres_control_s1 = ifill_control[pipe_mshr_readreq_threadid_s1];
        end
        2'd2:
        begin
            mshr_pipe_readres_control_s1 = ld_control[pipe_mshr_readreq_threadid_s1];
            mshr_pipe_readres_homeid_s1 = ld_homeid[pipe_mshr_readreq_threadid_s1];
        end
        2'd3:
        begin
            mshr_pipe_readres_control_s1 = st_control[pipe_mshr_readreq_threadid_s1];
            mshr_pipe_readres_homeid_s1 = st_homeid[pipe_mshr_readreq_threadid_s1];
        end
    endcase
    
    mshr_pipe_write_buffer_s2[127:0] = 128'b0;
    mshr_pipe_write_buffer_byte_mask_s2 = 16'b0;
    if (pipe_mshr_write_buffer_rd_en_s2)
    begin
        mshr_pipe_write_buffer_s2 = st_write_buffer[pipe_mshr_threadid_s2];
        mshr_pipe_write_buffer_byte_mask_s2 = st_write_buffer_byte_mask[pipe_mshr_threadid_s2];
    end
end
reg [127:0] bit_write_mask_s1;
always @ *
begin
    bit_write_mask_s1[0] = pipe_mshr_writereq_write_buffer_byte_mask_s1[0];
bit_write_mask_s1[1] = pipe_mshr_writereq_write_buffer_byte_mask_s1[0];
bit_write_mask_s1[2] = pipe_mshr_writereq_write_buffer_byte_mask_s1[0];
bit_write_mask_s1[3] = pipe_mshr_writereq_write_buffer_byte_mask_s1[0];
bit_write_mask_s1[4] = pipe_mshr_writereq_write_buffer_byte_mask_s1[0];
bit_write_mask_s1[5] = pipe_mshr_writereq_write_buffer_byte_mask_s1[0];
bit_write_mask_s1[6] = pipe_mshr_writereq_write_buffer_byte_mask_s1[0];
bit_write_mask_s1[7] = pipe_mshr_writereq_write_buffer_byte_mask_s1[0];
bit_write_mask_s1[8] = pipe_mshr_writereq_write_buffer_byte_mask_s1[1];
bit_write_mask_s1[9] = pipe_mshr_writereq_write_buffer_byte_mask_s1[1];
bit_write_mask_s1[10] = pipe_mshr_writereq_write_buffer_byte_mask_s1[1];
bit_write_mask_s1[11] = pipe_mshr_writereq_write_buffer_byte_mask_s1[1];
bit_write_mask_s1[12] = pipe_mshr_writereq_write_buffer_byte_mask_s1[1];
bit_write_mask_s1[13] = pipe_mshr_writereq_write_buffer_byte_mask_s1[1];
bit_write_mask_s1[14] = pipe_mshr_writereq_write_buffer_byte_mask_s1[1];
bit_write_mask_s1[15] = pipe_mshr_writereq_write_buffer_byte_mask_s1[1];
bit_write_mask_s1[16] = pipe_mshr_writereq_write_buffer_byte_mask_s1[2];
bit_write_mask_s1[17] = pipe_mshr_writereq_write_buffer_byte_mask_s1[2];
bit_write_mask_s1[18] = pipe_mshr_writereq_write_buffer_byte_mask_s1[2];
bit_write_mask_s1[19] = pipe_mshr_writereq_write_buffer_byte_mask_s1[2];
bit_write_mask_s1[20] = pipe_mshr_writereq_write_buffer_byte_mask_s1[2];
bit_write_mask_s1[21] = pipe_mshr_writereq_write_buffer_byte_mask_s1[2];
bit_write_mask_s1[22] = pipe_mshr_writereq_write_buffer_byte_mask_s1[2];
bit_write_mask_s1[23] = pipe_mshr_writereq_write_buffer_byte_mask_s1[2];
bit_write_mask_s1[24] = pipe_mshr_writereq_write_buffer_byte_mask_s1[3];
bit_write_mask_s1[25] = pipe_mshr_writereq_write_buffer_byte_mask_s1[3];
bit_write_mask_s1[26] = pipe_mshr_writereq_write_buffer_byte_mask_s1[3];
bit_write_mask_s1[27] = pipe_mshr_writereq_write_buffer_byte_mask_s1[3];
bit_write_mask_s1[28] = pipe_mshr_writereq_write_buffer_byte_mask_s1[3];
bit_write_mask_s1[29] = pipe_mshr_writereq_write_buffer_byte_mask_s1[3];
bit_write_mask_s1[30] = pipe_mshr_writereq_write_buffer_byte_mask_s1[3];
bit_write_mask_s1[31] = pipe_mshr_writereq_write_buffer_byte_mask_s1[3];
bit_write_mask_s1[32] = pipe_mshr_writereq_write_buffer_byte_mask_s1[4];
bit_write_mask_s1[33] = pipe_mshr_writereq_write_buffer_byte_mask_s1[4];
bit_write_mask_s1[34] = pipe_mshr_writereq_write_buffer_byte_mask_s1[4];
bit_write_mask_s1[35] = pipe_mshr_writereq_write_buffer_byte_mask_s1[4];
bit_write_mask_s1[36] = pipe_mshr_writereq_write_buffer_byte_mask_s1[4];
bit_write_mask_s1[37] = pipe_mshr_writereq_write_buffer_byte_mask_s1[4];
bit_write_mask_s1[38] = pipe_mshr_writereq_write_buffer_byte_mask_s1[4];
bit_write_mask_s1[39] = pipe_mshr_writereq_write_buffer_byte_mask_s1[4];
bit_write_mask_s1[40] = pipe_mshr_writereq_write_buffer_byte_mask_s1[5];
bit_write_mask_s1[41] = pipe_mshr_writereq_write_buffer_byte_mask_s1[5];
bit_write_mask_s1[42] = pipe_mshr_writereq_write_buffer_byte_mask_s1[5];
bit_write_mask_s1[43] = pipe_mshr_writereq_write_buffer_byte_mask_s1[5];
bit_write_mask_s1[44] = pipe_mshr_writereq_write_buffer_byte_mask_s1[5];
bit_write_mask_s1[45] = pipe_mshr_writereq_write_buffer_byte_mask_s1[5];
bit_write_mask_s1[46] = pipe_mshr_writereq_write_buffer_byte_mask_s1[5];
bit_write_mask_s1[47] = pipe_mshr_writereq_write_buffer_byte_mask_s1[5];
bit_write_mask_s1[48] = pipe_mshr_writereq_write_buffer_byte_mask_s1[6];
bit_write_mask_s1[49] = pipe_mshr_writereq_write_buffer_byte_mask_s1[6];
bit_write_mask_s1[50] = pipe_mshr_writereq_write_buffer_byte_mask_s1[6];
bit_write_mask_s1[51] = pipe_mshr_writereq_write_buffer_byte_mask_s1[6];
bit_write_mask_s1[52] = pipe_mshr_writereq_write_buffer_byte_mask_s1[6];
bit_write_mask_s1[53] = pipe_mshr_writereq_write_buffer_byte_mask_s1[6];
bit_write_mask_s1[54] = pipe_mshr_writereq_write_buffer_byte_mask_s1[6];
bit_write_mask_s1[55] = pipe_mshr_writereq_write_buffer_byte_mask_s1[6];
bit_write_mask_s1[56] = pipe_mshr_writereq_write_buffer_byte_mask_s1[7];
bit_write_mask_s1[57] = pipe_mshr_writereq_write_buffer_byte_mask_s1[7];
bit_write_mask_s1[58] = pipe_mshr_writereq_write_buffer_byte_mask_s1[7];
bit_write_mask_s1[59] = pipe_mshr_writereq_write_buffer_byte_mask_s1[7];
bit_write_mask_s1[60] = pipe_mshr_writereq_write_buffer_byte_mask_s1[7];
bit_write_mask_s1[61] = pipe_mshr_writereq_write_buffer_byte_mask_s1[7];
bit_write_mask_s1[62] = pipe_mshr_writereq_write_buffer_byte_mask_s1[7];
bit_write_mask_s1[63] = pipe_mshr_writereq_write_buffer_byte_mask_s1[7];
bit_write_mask_s1[64] = pipe_mshr_writereq_write_buffer_byte_mask_s1[8];
bit_write_mask_s1[65] = pipe_mshr_writereq_write_buffer_byte_mask_s1[8];
bit_write_mask_s1[66] = pipe_mshr_writereq_write_buffer_byte_mask_s1[8];
bit_write_mask_s1[67] = pipe_mshr_writereq_write_buffer_byte_mask_s1[8];
bit_write_mask_s1[68] = pipe_mshr_writereq_write_buffer_byte_mask_s1[8];
bit_write_mask_s1[69] = pipe_mshr_writereq_write_buffer_byte_mask_s1[8];
bit_write_mask_s1[70] = pipe_mshr_writereq_write_buffer_byte_mask_s1[8];
bit_write_mask_s1[71] = pipe_mshr_writereq_write_buffer_byte_mask_s1[8];
bit_write_mask_s1[72] = pipe_mshr_writereq_write_buffer_byte_mask_s1[9];
bit_write_mask_s1[73] = pipe_mshr_writereq_write_buffer_byte_mask_s1[9];
bit_write_mask_s1[74] = pipe_mshr_writereq_write_buffer_byte_mask_s1[9];
bit_write_mask_s1[75] = pipe_mshr_writereq_write_buffer_byte_mask_s1[9];
bit_write_mask_s1[76] = pipe_mshr_writereq_write_buffer_byte_mask_s1[9];
bit_write_mask_s1[77] = pipe_mshr_writereq_write_buffer_byte_mask_s1[9];
bit_write_mask_s1[78] = pipe_mshr_writereq_write_buffer_byte_mask_s1[9];
bit_write_mask_s1[79] = pipe_mshr_writereq_write_buffer_byte_mask_s1[9];
bit_write_mask_s1[80] = pipe_mshr_writereq_write_buffer_byte_mask_s1[10];
bit_write_mask_s1[81] = pipe_mshr_writereq_write_buffer_byte_mask_s1[10];
bit_write_mask_s1[82] = pipe_mshr_writereq_write_buffer_byte_mask_s1[10];
bit_write_mask_s1[83] = pipe_mshr_writereq_write_buffer_byte_mask_s1[10];
bit_write_mask_s1[84] = pipe_mshr_writereq_write_buffer_byte_mask_s1[10];
bit_write_mask_s1[85] = pipe_mshr_writereq_write_buffer_byte_mask_s1[10];
bit_write_mask_s1[86] = pipe_mshr_writereq_write_buffer_byte_mask_s1[10];
bit_write_mask_s1[87] = pipe_mshr_writereq_write_buffer_byte_mask_s1[10];
bit_write_mask_s1[88] = pipe_mshr_writereq_write_buffer_byte_mask_s1[11];
bit_write_mask_s1[89] = pipe_mshr_writereq_write_buffer_byte_mask_s1[11];
bit_write_mask_s1[90] = pipe_mshr_writereq_write_buffer_byte_mask_s1[11];
bit_write_mask_s1[91] = pipe_mshr_writereq_write_buffer_byte_mask_s1[11];
bit_write_mask_s1[92] = pipe_mshr_writereq_write_buffer_byte_mask_s1[11];
bit_write_mask_s1[93] = pipe_mshr_writereq_write_buffer_byte_mask_s1[11];
bit_write_mask_s1[94] = pipe_mshr_writereq_write_buffer_byte_mask_s1[11];
bit_write_mask_s1[95] = pipe_mshr_writereq_write_buffer_byte_mask_s1[11];
bit_write_mask_s1[96] = pipe_mshr_writereq_write_buffer_byte_mask_s1[12];
bit_write_mask_s1[97] = pipe_mshr_writereq_write_buffer_byte_mask_s1[12];
bit_write_mask_s1[98] = pipe_mshr_writereq_write_buffer_byte_mask_s1[12];
bit_write_mask_s1[99] = pipe_mshr_writereq_write_buffer_byte_mask_s1[12];
bit_write_mask_s1[100] = pipe_mshr_writereq_write_buffer_byte_mask_s1[12];
bit_write_mask_s1[101] = pipe_mshr_writereq_write_buffer_byte_mask_s1[12];
bit_write_mask_s1[102] = pipe_mshr_writereq_write_buffer_byte_mask_s1[12];
bit_write_mask_s1[103] = pipe_mshr_writereq_write_buffer_byte_mask_s1[12];
bit_write_mask_s1[104] = pipe_mshr_writereq_write_buffer_byte_mask_s1[13];
bit_write_mask_s1[105] = pipe_mshr_writereq_write_buffer_byte_mask_s1[13];
bit_write_mask_s1[106] = pipe_mshr_writereq_write_buffer_byte_mask_s1[13];
bit_write_mask_s1[107] = pipe_mshr_writereq_write_buffer_byte_mask_s1[13];
bit_write_mask_s1[108] = pipe_mshr_writereq_write_buffer_byte_mask_s1[13];
bit_write_mask_s1[109] = pipe_mshr_writereq_write_buffer_byte_mask_s1[13];
bit_write_mask_s1[110] = pipe_mshr_writereq_write_buffer_byte_mask_s1[13];
bit_write_mask_s1[111] = pipe_mshr_writereq_write_buffer_byte_mask_s1[13];
bit_write_mask_s1[112] = pipe_mshr_writereq_write_buffer_byte_mask_s1[14];
bit_write_mask_s1[113] = pipe_mshr_writereq_write_buffer_byte_mask_s1[14];
bit_write_mask_s1[114] = pipe_mshr_writereq_write_buffer_byte_mask_s1[14];
bit_write_mask_s1[115] = pipe_mshr_writereq_write_buffer_byte_mask_s1[14];
bit_write_mask_s1[116] = pipe_mshr_writereq_write_buffer_byte_mask_s1[14];
bit_write_mask_s1[117] = pipe_mshr_writereq_write_buffer_byte_mask_s1[14];
bit_write_mask_s1[118] = pipe_mshr_writereq_write_buffer_byte_mask_s1[14];
bit_write_mask_s1[119] = pipe_mshr_writereq_write_buffer_byte_mask_s1[14];
bit_write_mask_s1[120] = pipe_mshr_writereq_write_buffer_byte_mask_s1[15];
bit_write_mask_s1[121] = pipe_mshr_writereq_write_buffer_byte_mask_s1[15];
bit_write_mask_s1[122] = pipe_mshr_writereq_write_buffer_byte_mask_s1[15];
bit_write_mask_s1[123] = pipe_mshr_writereq_write_buffer_byte_mask_s1[15];
bit_write_mask_s1[124] = pipe_mshr_writereq_write_buffer_byte_mask_s1[15];
bit_write_mask_s1[125] = pipe_mshr_writereq_write_buffer_byte_mask_s1[15];
bit_write_mask_s1[126] = pipe_mshr_writereq_write_buffer_byte_mask_s1[15];
bit_write_mask_s1[127] = pipe_mshr_writereq_write_buffer_byte_mask_s1[15];
end
always @ (posedge clk)
begin
    if (pipe_mshr_writereq_val_s1 && (op_s1 == 3'b001))
    begin
        case (mshrid_s1)
            2'd1:
            begin
                
                ifill_control[threadid_s1] <= pipe_mshr_writereq_control_s1;
            end
            2'd2:
            begin
                ld_address[threadid_s1] <= pipe_mshr_writereq_address_s1;
                ld_control[threadid_s1] <= pipe_mshr_writereq_control_s1;
            end
            2'd3:
            begin
                st_address[threadid_s1] <= pipe_mshr_writereq_address_s1;
                st_control[threadid_s1] <= pipe_mshr_writereq_control_s1;
                st_write_buffer[threadid_s1] <= (pipe_mshr_writereq_write_buffer_data_s1 & bit_write_mask_s1);
                st_write_buffer_byte_mask[threadid_s1] <= pipe_mshr_writereq_write_buffer_byte_mask_s1;
            end
        endcase
    end 
    else if (pipe_mshr_writereq_val_s1 && op_s1 == 3'b100)
    begin
        st_write_buffer[threadid_s1] <= ((st_write_buffer[threadid_s1] & ~bit_write_mask_s1) | (pipe_mshr_writereq_write_buffer_data_s1 & bit_write_mask_s1));
        st_write_buffer_byte_mask[threadid_s1] <= (st_write_buffer_byte_mask[threadid_s1] | pipe_mshr_writereq_write_buffer_byte_mask_s1);
    end 
end
always @ (posedge clk)
begin
    if (pipe_mshr_val_s3 && op_s3 == 3'b011)
    begin
        st_state[threadid_s3] <= pipe_mshr_write_update_state_s3;
        st_way[threadid_s3] <= pipe_mshr_write_update_way_s3;
    end 
end 
reg [2-1:0] ld_val_next;
reg [2-1:0] st_val_next;
reg [2-1:0] ifill_val_next;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        ld_val <= 0;
        st_val <= 0;
        ifill_val <= 0;
    end
    else
    begin
        ld_val <= ld_val_next;
        st_val <= st_val_next;
        ifill_val <= ifill_val_next;
    end
end
reg [2-1:0] ld_alloc_mask;
reg [2-1:0] st_alloc_mask;
reg [2-1:0] ifill_alloc_mask;
reg [2-1:0] ld_dealloc_mask;
reg [2-1:0] st_dealloc_mask;
reg [2-1:0] ifill_dealloc_mask;
always @ *
begin
    
    
    
    
    
    
    
    
    
    
    
    
    ld_alloc_mask = 0;
    st_alloc_mask = 0;
    ifill_alloc_mask = 0;
    if (pipe_mshr_writereq_val_s1 && (op_s1 == 3'b001))
    begin
        if (mshrid_s1 == 2'd2)
            ld_alloc_mask[threadid_s1] = 1'b1;
        else if (mshrid_s1 == 2'd3)
            st_alloc_mask[threadid_s1] = 1'b1;
        else if (mshrid_s1 == 2'd1)
            ifill_alloc_mask[threadid_s1] = 1'b1;
    end
    ld_dealloc_mask = 0;
    st_dealloc_mask = 0;
    ifill_dealloc_mask = 0;
    if (pipe_mshr_val_s3 && (op_s3 == 3'b010))
    begin
        if (mshrid_s3 == 2'd2)
            ld_dealloc_mask[threadid_s3] = 1'b1;
        else if (mshrid_s3 == 2'd3)
            st_dealloc_mask[threadid_s3] = 1'b1;
        else if (mshrid_s3 == 2'd1)
            ifill_dealloc_mask[threadid_s3] = 1'b1;
    end
    ld_val_next = ld_val;
    st_val_next = st_val;
    ifill_val_next = ifill_val;
    ld_val_next = (ld_val & ~ld_dealloc_mask) | ld_alloc_mask;
    st_val_next = (st_val & ~st_dealloc_mask) | st_alloc_mask;
    ifill_val_next = (ifill_val & ~ifill_dealloc_mask) | ifill_alloc_mask;
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        st_homeid[0] <= 0;
        st_homeid[1] <= 0;
        ld_homeid[0] <= 0;
        ld_homeid[1] <= 0;
    end
    else
    begin
        if (noc1buffer_mshr_homeid_write_val_s4)
        begin
            if (noc1buffer_mshr_homeid_write_mshrid_s4 == 2'd2)
                ld_homeid[noc1buffer_mshr_homeid_write_threadid_s4] <= noc1buffer_mshr_homeid_write_data_s4;
            else if (noc1buffer_mshr_homeid_write_mshrid_s4 == 2'd3)
                st_homeid[noc1buffer_mshr_homeid_write_threadid_s4] <= noc1buffer_mshr_homeid_write_data_s4;
        end
    end
end
endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
module l15_pipeline(
    input wire clk,
    input wire rst_n,
    
    input wire [5-1:0] pcxdecoder_l15_rqtype,
    input wire [4-1:0] pcxdecoder_l15_amo_op,
    input wire pcxdecoder_l15_nc,
    input wire [3-1:0] pcxdecoder_l15_size,
    
    input wire [0:0] pcxdecoder_l15_threadid,
    input wire pcxdecoder_l15_prefetch,
    input wire pcxdecoder_l15_blockstore,
    input wire pcxdecoder_l15_blockinitstore,
    input wire [2-1:0] pcxdecoder_l15_l1rplway,
    input wire pcxdecoder_l15_val,
    input wire [39:0] pcxdecoder_l15_address,
    input wire [33-1:0] pcxdecoder_l15_csm_data,
    input wire [63:0] pcxdecoder_l15_data,
    input wire [63:0] pcxdecoder_l15_data_next_entry,
    input wire pcxdecoder_l15_invalidate_cacheline,
    
    input wire noc2decoder_l15_val,
    input wire [2-1:0] noc2decoder_l15_mshrid,
    input wire [0:0] noc2decoder_l15_threadid,
    input wire noc2decoder_l15_hmc_fill,
    input wire noc2decoder_l15_l2miss,
    input wire noc2decoder_l15_icache_type,
    input wire noc2decoder_l15_f4b, 
    input wire [8-1:0] noc2decoder_l15_reqtype, 
    input wire [2-1:0] noc2decoder_l15_ack_state,
    input wire [3:0] noc2decoder_l15_fwd_subcacheline_vector,
    input wire [63:0] noc2decoder_l15_data_0,
    input wire [63:0] noc2decoder_l15_data_1,
    input wire [63:0] noc2decoder_l15_data_2,
    input wire [63:0] noc2decoder_l15_data_3,
    input wire [39:0] noc2decoder_l15_address,
    input wire [(14+8+8)-1:0] noc2decoder_l15_src_homeid,
    input wire [3-1:0] noc2decoder_l15_csm_mshrid,
    
    input wire cpxencoder_l15_req_ack,
    
    input wire noc1encoder_l15_req_sent,
    input wire [2-1:0] noc1encoder_l15_req_data_sent,
    input wire noc3encoder_l15_req_ack,
    
    input wire [63:0] config_l15_read_res_data_s3,
    
    
    output reg l15_dtag_val_s1,
    output reg l15_dtag_rw_s1,
    output reg [((9-2))-1:0] l15_dtag_index_s1,
    output reg [33*4-1:0] l15_dtag_write_data_s1,
    output reg [33*4-1:0] l15_dtag_write_mask_s1,
    input wire [33*4-1:0] dtag_l15_dout_s2,
    
    output reg l15_dcache_val_s2,
    output reg l15_dcache_rw_s2,
    output reg [(((9-2))+2)-1:0] l15_dcache_index_s2,
    output reg [127:0] l15_dcache_write_data_s2,
    output reg [127:0] l15_dcache_write_mask_s2,
    input wire [127:0] dcache_l15_dout_s3,
    
    output reg l15_mesi_read_val_s1,
    output reg [((9-2))-1:0] l15_mesi_read_index_s1,
    input wire [7:0] mesi_l15_dout_s2,
    output reg l15_mesi_write_val_s2,
    output reg [((9-2))-1:0] l15_mesi_write_index_s2,
    output reg [7:0] l15_mesi_write_mask_s2,
    output reg [7:0] l15_mesi_write_data_s2,
    
    output reg l15_lrsc_flag_read_val_s1,
    output reg [((9-2))-1:0] l15_lrsc_flag_read_index_s1,
    input wire [3:0] lrsc_flag_l15_dout_s2,
    output reg l15_lrsc_flag_write_val_s2,
    output reg [((9-2))-1:0] l15_lrsc_flag_write_index_s2,
    output reg [3:0] l15_lrsc_flag_write_mask_s2,
    output reg [3:0] l15_lrsc_flag_write_data_s2,
    
    output reg l15_lruarray_read_val_s1,
    output reg [((9-2))-1:0] l15_lruarray_read_index_s1,
    input wire [(2 + 4)-1:0] lruarray_l15_dout_s2,
    output reg l15_lruarray_write_val_s3,
    output reg [((9-2))-1:0] l15_lruarray_write_index_s3,
    output reg [(2 + 4)-1:0] l15_lruarray_write_mask_s3,    
    output reg [(2 + 4)-1:0] l15_lruarray_write_data_s3,
    
    
    input wire [14 + 8 + 8-1:0] hmt_l15_dout_s3,
    output reg [14 + 8 + 8-1:0] l15_hmt_write_data_s2,
    output reg [14 + 8 + 8-1:0] l15_hmt_write_mask_s2,
    
    
    output reg l15_wmt_read_val_s2,
    output reg [6:0] l15_wmt_read_index_s2,
    input wire [4*((2+0)+1)-1:0] wmt_l15_data_s3,
    output reg l15_wmt_write_val_s3,
    output reg [6:0] l15_wmt_write_index_s3,
    output reg [4*((2+0)+1)-1:0] l15_wmt_write_mask_s3,
    output reg [4*((2+0)+1)-1:0] l15_wmt_write_data_s3,
    
    
    output reg pipe_mshr_writereq_val_s1,
    output reg [3-1:0] pipe_mshr_writereq_op_s1,   
    output reg [39:0] pipe_mshr_writereq_address_s1,
    output reg [127:0] pipe_mshr_writereq_write_buffer_data_s1,
    output reg [15:0] pipe_mshr_writereq_write_buffer_byte_mask_s1,
    output reg [((((((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) + 1) + 1) + 1)-1:0] pipe_mshr_writereq_control_s1,
    output reg [2-1:0] pipe_mshr_writereq_mshrid_s1,
    output reg [0:0] pipe_mshr_writereq_threadid_s1,
    
    output reg [0:0] pipe_mshr_readreq_threadid_s1,
    output reg [2-1:0] pipe_mshr_readreq_mshrid_s1,
    input wire [((((((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) + 1) + 1) + 1)-1:0] mshr_pipe_readres_control_s1,
    input wire [(14+8+8)-1:0] mshr_pipe_readres_homeid_s1,
    
        
    input wire [(4*2)-1:0] mshr_pipe_vals_s1,
    input wire [(40*2)-1:0] mshr_pipe_ld_address,
    input wire [(40*2)-1:0] mshr_pipe_st_address,
    input wire [(2*2)-1:0] mshr_pipe_st_way_s1,
    input wire [(2*2)-1:0] mshr_pipe_st_state_s1,
    
    output reg pipe_mshr_write_buffer_rd_en_s2,
    output reg [0:0] pipe_mshr_threadid_s2,
    input wire [127:0] mshr_pipe_write_buffer_s2,
    input wire [15:0] mshr_pipe_write_buffer_byte_mask_s2,
    
    output reg pipe_mshr_val_s3,
    output reg [3-1:0] pipe_mshr_op_s3,
    output reg [2-1:0] pipe_mshr_mshrid_s3,
    output reg [0:0] pipe_mshr_threadid_s3,
    output reg [2-1:0] pipe_mshr_write_update_state_s3,
    output reg [1:0] pipe_mshr_write_update_way_s3,
    
    
    output reg l15_cpxencoder_val,
    output reg [3:0] l15_cpxencoder_returntype,
    output reg l15_cpxencoder_l2miss,
    output reg [1:0] l15_cpxencoder_error,  
    output reg l15_cpxencoder_noncacheable,
    output reg l15_cpxencoder_atomic,
    output reg [0:0] l15_cpxencoder_threadid,
    output reg l15_cpxencoder_prefetch,
    output reg l15_cpxencoder_f4b,
    output reg [63:0] l15_cpxencoder_data_0,
    output reg [63:0] l15_cpxencoder_data_1,
    output reg [63:0] l15_cpxencoder_data_2,
    output reg [63:0] l15_cpxencoder_data_3,
    output reg l15_cpxencoder_inval_icache_all_way,
    output reg l15_cpxencoder_inval_dcache_all_way,         
    output reg [15:4] l15_cpxencoder_inval_address_15_4,
    output reg l15_cpxencoder_cross_invalidate,             
    output reg [1:0] l15_cpxencoder_cross_invalidate_way,   
    output reg l15_cpxencoder_inval_dcache_inval,
    output reg l15_cpxencoder_inval_icache_inval,           
    output reg l15_cpxencoder_blockinitstore,
    output reg [1:0] l15_cpxencoder_inval_way,
    
    output reg l15_noc1buffer_req_val,
    output reg [5-1:0] l15_noc1buffer_req_type,
    output reg [0:0] l15_noc1buffer_req_threadid,
    output reg [2-1:0] l15_noc1buffer_req_mshrid,
    output reg [39:0] l15_noc1buffer_req_address,
    output reg l15_noc1buffer_req_non_cacheable,
    output reg [2:0] l15_noc1buffer_req_size,
    output reg l15_noc1buffer_req_prefetch,
    output reg [33-1:0] l15_noc1buffer_req_csm_data,
    output reg [63:0] l15_noc1buffer_req_data_0,
    output reg [63:0] l15_noc1buffer_req_data_1,
    
    
    
    output reg l15_noc3encoder_req_val,
    output reg [3-1:0] l15_noc3encoder_req_type,
    output reg [63:0] l15_noc3encoder_req_data_0,
    output reg [63:0] l15_noc3encoder_req_data_1,
    output reg [2-1:0] l15_noc3encoder_req_mshrid,
    output reg [1:0] l15_noc3encoder_req_sequenceid,
    output reg [0:0] l15_noc3encoder_req_threadid,
    output reg [39:0] l15_noc3encoder_req_address,
    output reg l15_noc3encoder_req_with_data,
    output reg l15_noc3encoder_req_was_inval,
    output reg [3:0] l15_noc3encoder_req_fwdack_vector,
    output reg [(14+8+8)-1:0] l15_noc3encoder_req_homeid,
    
    output reg l15_pcxdecoder_ack,
    output reg l15_noc2decoder_ack,
    output reg l15_pcxdecoder_header_ack,
    output reg l15_noc2decoder_header_ack,
    
    output reg [40-1:0] l15_csm_req_address_s2,
    output reg l15_csm_req_val_s2,
    output reg l15_csm_stall_s3,
    output reg [3-1:0] l15_csm_req_ticket_s2,
    
    output reg  l15_csm_req_type_s2,     
    output reg [127:0] l15_csm_req_data_s2, 
    output reg [33-1:0] l15_csm_req_pcx_data_s2, 
    input wire csm_l15_res_val_s3,
    input wire [63:0] csm_l15_res_data_s3,
    
    output reg [3-1:0] l15_noc1buffer_req_csm_ticket,
    output reg [(14+8+8)-1:0] l15_noc1buffer_req_homeid,
    output reg l15_noc1buffer_req_homeid_val,
    
    output reg l15_config_req_val_s2,
    output reg l15_config_req_rw_s2,
    output reg [63:0] l15_config_write_req_data_s2,
    output reg [15:8] l15_config_req_address_s2
    );
reg stall_s1;
reg stall_s2;
reg stall_s3;
reg val_s1; 
reg val_s2;
reg val_s3;
reg pcx_ack_s1;
reg pcx_ack_s2;
reg pcx_ack_s3;
reg noc2_ack_s1;
reg noc2_ack_s2;
reg noc2_ack_s3;
reg [3-1:0] fetch_state_s1;
reg [3-1:0] fetch_state_next_s1;
reg [((9-2))-1:0] cache_index_s2;
reg [((6 + 4) - 4 + 1)-1:0] cache_index_l1d_s2;
reg [((9-2))-1:0] cache_index_s3;
reg [((6 + 4) - 4 + 1)-1:0] cache_index_l1d_s3;
reg [2-1:0] lru_way_s2;
always @ *
begin
    l15_pcxdecoder_ack = pcx_ack_s1 || pcx_ack_s2 || pcx_ack_s3;
    l15_noc2decoder_ack = noc2_ack_s1 || noc2_ack_s2 || noc2_ack_s3;
end
reg [(40 - 4 - ((9-2)))-1:0] predecode_dtag_write_data_s1;
reg [((9-2))-1:0] predecode_cache_index_s1;
reg [((((((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) + 1) + 1) + 1)-1:0] predecode_mshr_read_control_s1;
reg [(14+8+8)-1:0] predecode_mshr_read_homeid_s1;
reg [6-1:0] predecode_reqtype_s1;
reg [39:0] predecode_address_s1;
reg [39:0] predecode_address_plus0_s1;
reg [39:0] predecode_address_plus1_s1;
reg [39:0] predecode_address_plus2_s1;
reg [39:0] predecode_address_plus3_s1;
reg [2:0] predecode_size_s1;
reg [0:0] predecode_threadid_s1;
reg [2-1:0] predecode_l1_replacement_way_s1;
reg predecode_non_cacheable_s1;
reg predecode_is_last_inval_s1;
reg predecode_blockstore_bit_s1;
reg predecode_blockstore_init_s1;
reg predecode_prefetch_bit_s1;
reg predecode_l2_miss_s1;
reg predecode_f4b_s1;
reg predecode_dcache_load_s1;
reg predecode_atomic_s1;
reg predecode_dcache_noc2_store_im_s1;
reg predecode_dcache_noc2_store_sm_s1;
reg predecode_icache_bit_s1;
reg predecode_noc2_inval_s1;
reg predecode_val_s1;
reg [2-1:0] predecode_source_s1;
reg predecode_interrupt_broadcast_s1;
reg [3:0] predecode_fwd_subcacheline_vector_s1;
always @ *
begin
    predecode_source_s1 = 0;
    case (fetch_state_s1)
        3'd0:
            predecode_source_s1 = (noc2decoder_l15_val) ? 2'd2 :
                                    (pcxdecoder_l15_val) ? 2'd1 :
                                                            2'd0;
        3'd1:
            predecode_source_s1 = 2'd1;
        3'd5:
            predecode_source_s1 = 2'd2;
        3'd2,
        3'd3,
        3'd4:
            predecode_source_s1 = 2'd2;
        3'd6:
            predecode_source_s1 = 2'd2;
    endcase
end
reg [4-1:0] mshr_val_array [1:0];
reg [2-1:0] mshr_st_state_array [1:0];
reg [39:0] mshr_st_address_array [1:0];
reg [39:0] mshr_ld_address_array [1:0];
reg [2-1:0] mshr_st_way_array [1:0];
always @ *
begin
    pipe_mshr_readreq_mshrid_s1 = noc2decoder_l15_mshrid;
    pipe_mshr_readreq_threadid_s1 = noc2decoder_l15_threadid;
    predecode_mshr_read_control_s1 = mshr_pipe_readres_control_s1;
    
    predecode_mshr_read_homeid_s1 = mshr_pipe_readres_homeid_s1;
    
    mshr_val_array[0] = mshr_pipe_vals_s1[4*1 - 1 -: 4];
    mshr_st_state_array[0] = mshr_pipe_st_state_s1[2*1 - 1 -: 2];
    mshr_st_address_array[0] = mshr_pipe_st_address[40*1 - 1 -: 40];
    mshr_ld_address_array[0] = mshr_pipe_ld_address[40*1 - 1 -: 40];
    mshr_st_way_array[0] = mshr_pipe_st_way_s1[2*1 - 1 -: 2];
    mshr_val_array[1] = mshr_pipe_vals_s1[4*2 - 1 -: 4];
    mshr_st_state_array[1] = mshr_pipe_st_state_s1[2*2 - 1 -: 2];
    mshr_st_address_array[1] = mshr_pipe_st_address[40*2 - 1 -: 40];
    mshr_ld_address_array[1] = mshr_pipe_ld_address[40*2 - 1 -: 40];
    mshr_st_way_array[1] = mshr_pipe_st_way_s1[2*2 - 1 -: 2];
end
reg [8-1:0] predecode_special_access_s1;
reg predecode_is_pcx_config_asi_s1;
reg predecode_is_pcx_diag_data_access_s1;
reg predecode_is_pcx_diag_line_flush_s1;
reg predecode_is_hmc_diag_access_s1;
reg predecode_is_hmc_flush_s1;
always @ *
begin
    predecode_special_access_s1 = pcxdecoder_l15_address[39:32];
    predecode_is_pcx_config_asi_s1 = predecode_special_access_s1 == 8'hba;
    predecode_is_pcx_diag_data_access_s1 = predecode_special_access_s1 == 8'hb0;
    predecode_is_pcx_diag_line_flush_s1 = predecode_special_access_s1 == 8'hb3;
    predecode_is_hmc_diag_access_s1 = predecode_special_access_s1 == 8'hb2;
    predecode_is_hmc_flush_s1 = predecode_special_access_s1 == 8'hb5;
end
reg predecode_tagcheck_matched_t0ld_s1;
reg predecode_tagcheck_matched_t0st_s1;
reg predecode_tagcheck_matched_t1ld_s1;
reg predecode_tagcheck_matched_t1st_s1;
reg predecode_int_vec_dis_s1;
reg predecode_tagcheck_matched_s1;
reg [19:4] predecode_partial_tag_s1;
reg predecode_hit_stbuf_s1;
reg [0:0] predecode_hit_stbuf_threadid_s1;
wire [39:0] constant_int_vec_dis_address = 40'h9800000800;
always @ *
begin
    predecode_reqtype_s1 = 0;
    predecode_address_s1 = 0;
    predecode_address_plus0_s1 = 0;
    predecode_address_plus1_s1 = 0;
    predecode_address_plus2_s1 = 0;
    predecode_address_plus3_s1 = 0;
    predecode_is_last_inval_s1 = 0;
    
    predecode_size_s1 = 0;
    predecode_threadid_s1 = 0;
    predecode_l1_replacement_way_s1 = 0;
    predecode_non_cacheable_s1 = 0;
    predecode_blockstore_bit_s1 = 0;
    predecode_blockstore_init_s1 = 0;
    predecode_prefetch_bit_s1 = 0;
    
    predecode_l2_miss_s1 = 0;
    predecode_f4b_s1 = 0;
    predecode_icache_bit_s1 = 0;
    predecode_dcache_load_s1 = 0;
    predecode_atomic_s1 = 0;
    predecode_dcache_noc2_store_im_s1 = 0;
    predecode_dcache_noc2_store_sm_s1 = 0;
    predecode_noc2_inval_s1 = 0;
    predecode_fwd_subcacheline_vector_s1 = 0;
    predecode_interrupt_broadcast_s1 = 0;
    case (predecode_source_s1)
        2'd2:
        begin
            
            predecode_size_s1 = predecode_mshr_read_control_s1[(((((0 + 1) + 1) + 1) + 1) + 3) -: 3];
            
            predecode_threadid_s1[0:0] = noc2decoder_l15_threadid[0:0];
            predecode_l1_replacement_way_s1 = predecode_mshr_read_control_s1[(((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) -: 2];
            predecode_non_cacheable_s1 = predecode_mshr_read_control_s1[((((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) + 1) -: 1];
            
            predecode_blockstore_bit_s1 = predecode_mshr_read_control_s1[(((((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) + 1) + 1) -: 1];
            predecode_blockstore_init_s1 = predecode_mshr_read_control_s1[(0 + 1) -: 1];
            predecode_prefetch_bit_s1 = predecode_mshr_read_control_s1[0 -: 1];
            
            predecode_l2_miss_s1 = noc2decoder_l15_l2miss;
            predecode_f4b_s1 = noc2decoder_l15_f4b;
            predecode_atomic_s1 = predecode_mshr_read_control_s1[(((0 + 1) + 1) + 1)];
            predecode_dcache_load_s1 = predecode_mshr_read_control_s1[((0 + 1) + 1)];
            predecode_fwd_subcacheline_vector_s1 = noc2decoder_l15_fwd_subcacheline_vector;
            predecode_dcache_noc2_store_im_s1 = mshr_st_state_array[predecode_threadid_s1] == 2'b10;
            predecode_dcache_noc2_store_sm_s1 = mshr_st_state_array[predecode_threadid_s1] == 2'b01;
            predecode_address_plus0_s1 = {noc2decoder_l15_address[39:6], 2'b00, noc2decoder_l15_address[3:0]};
            predecode_address_plus1_s1 = {noc2decoder_l15_address[39:6], 2'b01, noc2decoder_l15_address[3:0]};
            predecode_address_plus2_s1 = {noc2decoder_l15_address[39:6], 2'b10, noc2decoder_l15_address[3:0]};
            predecode_address_plus3_s1 = {noc2decoder_l15_address[39:6], 2'b11, noc2decoder_l15_address[3:0]};
            if (noc2decoder_l15_icache_type)
                predecode_is_last_inval_s1 = ((fetch_state_s1 == 3'd6) && (predecode_fwd_subcacheline_vector_s1[3:2] == 2'b11)) ||
                                             ((fetch_state_s1 == 3'd0) && (predecode_fwd_subcacheline_vector_s1[3:0] == 4'b0011));
                
            else
                predecode_is_last_inval_s1 = ((fetch_state_s1 == 3'd4) && (predecode_fwd_subcacheline_vector_s1[3])) ||
                                             ((fetch_state_s1 == 3'd3) && (predecode_fwd_subcacheline_vector_s1[3:2] == 2'b01)) ||
                                             ((fetch_state_s1 == 3'd2) && (predecode_fwd_subcacheline_vector_s1[3:1] == 3'b001)) ||
                                             ((fetch_state_s1 == 3'd0) && (predecode_fwd_subcacheline_vector_s1[3:0] == 4'b0001));
            
            
            
            case(noc2decoder_l15_reqtype)
                8'd17:
                begin
                    predecode_icache_bit_s1 = noc2decoder_l15_icache_type;
                    if (predecode_icache_bit_s1)
                    begin
                        
                            predecode_reqtype_s1 = 6'd18;
                        
                        
                        predecode_address_s1 = (fetch_state_s1 == 3'd6) ? predecode_address_plus2_s1 :
                                                                                                predecode_address_plus0_s1;
                    end
                    else
                    begin
                        predecode_reqtype_s1 = 6'd6;
                        predecode_address_s1 = (fetch_state_s1 == 3'd2) ? predecode_address_plus1_s1 :
                                                (fetch_state_s1 == 3'd3) ? predecode_address_plus2_s1 :
                                                (fetch_state_s1 == 3'd4) ? predecode_address_plus3_s1 :
                                                                                                predecode_address_plus0_s1;
                    end
                end
                8'd18:
                begin
                    predecode_icache_bit_s1 = noc2decoder_l15_icache_type;
                    if (predecode_icache_bit_s1)
                    begin
                        
                            predecode_reqtype_s1 = 6'd18;
                        
                        
                        predecode_address_s1 = (fetch_state_s1 == 3'd6) ? predecode_address_plus2_s1 :
                                                                                                predecode_address_plus0_s1;
                    end
                    else
                    begin
                        predecode_reqtype_s1 = 6'd6;
                        predecode_noc2_inval_s1 = 1'b1;
                        predecode_address_s1 = (fetch_state_s1 == 3'd2) ? predecode_address_plus1_s1 :
                                                (fetch_state_s1 == 3'd3) ? predecode_address_plus2_s1 :
                                                (fetch_state_s1 == 3'd4) ? predecode_address_plus3_s1 :
                                                                                                predecode_address_plus0_s1;
                    end
                end
                8'd16:
                begin
                    predecode_icache_bit_s1 = noc2decoder_l15_icache_type;
                    if (predecode_icache_bit_s1)
                    begin
                        
                            predecode_reqtype_s1 = 6'd18;
                        
                        
                        predecode_address_s1 = (fetch_state_s1 == 3'd6) ? predecode_address_plus2_s1 :
                                                                                                predecode_address_plus0_s1;
                    end
                    else
                    begin
                        predecode_reqtype_s1 = 6'd7;
                        predecode_address_s1 = (fetch_state_s1 == 3'd2) ? predecode_address_plus1_s1 :
                                                (fetch_state_s1 == 3'd3) ? predecode_address_plus2_s1 :
                                                (fetch_state_s1 == 3'd4) ? predecode_address_plus3_s1 :
                                                                                                predecode_address_plus0_s1;
                    end
                end
                8'd29, 8'd26:
                begin
                    predecode_icache_bit_s1 = predecode_mshr_read_control_s1[((((0 + 1) + 1) + 1) + 1)];
                    if (noc2decoder_l15_mshrid == 2'd2)
                        predecode_address_s1 = mshr_ld_address_array[noc2decoder_l15_threadid];
                    else if (noc2decoder_l15_mshrid == 2'd3)
                        predecode_address_s1 = mshr_st_address_array[noc2decoder_l15_threadid];
                    if (noc2decoder_l15_hmc_fill)
                    begin
                        predecode_reqtype_s1 = 6'd28;
                        predecode_address_s1 = 0;   
                    end
                    else
                    if (predecode_non_cacheable_s1)
                    begin
                        if (predecode_icache_bit_s1)
                            predecode_reqtype_s1 = 6'd9;
                        else if (predecode_dcache_load_s1)
                            predecode_reqtype_s1 = 6'd8;
                        else if (predecode_atomic_s1)
                            predecode_reqtype_s1 = 6'd14;
                        else
                            predecode_reqtype_s1 = 6'd1; 
                    end
                    else
                    begin
                        if (predecode_icache_bit_s1)
                            predecode_reqtype_s1 = 6'd9;
                        else if (predecode_atomic_s1)
                            predecode_reqtype_s1 = 6'd46;
                            
                            
                        else if (predecode_dcache_load_s1)
                            predecode_reqtype_s1 = 6'd10;
                        else if (predecode_dcache_noc2_store_im_s1)
                            predecode_reqtype_s1 = 6'd11;
                        else if (predecode_dcache_noc2_store_sm_s1)
                            predecode_reqtype_s1 = 6'd12;
                        else
                            predecode_reqtype_s1 = 6'd1; 
                    end
                end
                8'd28, 8'd27:
                begin
                    predecode_icache_bit_s1 = predecode_mshr_read_control_s1[((((0 + 1) + 1) + 1) + 1)];
                    predecode_address_s1 = mshr_st_address_array[noc2decoder_l15_threadid];
                    
                    if (noc2decoder_l15_mshrid == 2'd3)
                        predecode_reqtype_s1 = 6'd13;
                    else
                    begin
                        predecode_reqtype_s1 = 6'd32;
                        predecode_address_s1 = 0; 
                    end
                end
                8'd33:
                begin
                    predecode_reqtype_s1 = 6'd20;
                end
            endcase
        end
        2'd1:
        begin
            predecode_address_s1 = pcxdecoder_l15_address;
            predecode_size_s1 = pcxdecoder_l15_size;
            predecode_threadid_s1[0:0] = pcxdecoder_l15_threadid[0:0];
            predecode_l1_replacement_way_s1 = pcxdecoder_l15_l1rplway;
            predecode_non_cacheable_s1 = pcxdecoder_l15_nc;
            predecode_blockstore_bit_s1 = pcxdecoder_l15_blockstore;
            predecode_blockstore_init_s1 = pcxdecoder_l15_blockinitstore;
            predecode_prefetch_bit_s1 = pcxdecoder_l15_prefetch;
            
            case(pcxdecoder_l15_rqtype)
                5'b00000:
                begin
                    if (predecode_is_pcx_config_asi_s1)
                        predecode_reqtype_s1 = 6'd24;
                    else if (predecode_is_pcx_diag_data_access_s1)
                        predecode_reqtype_s1 = 6'd25;
                    else if (predecode_is_hmc_diag_access_s1)
                        predecode_reqtype_s1 = 6'd29;
                    else if (predecode_prefetch_bit_s1)
                        predecode_reqtype_s1 = 6'd16;
                    else if (predecode_non_cacheable_s1)
                        predecode_reqtype_s1 = 6'd15;
                    else if (pcxdecoder_l15_invalidate_cacheline)
                        predecode_reqtype_s1 = 6'd34;
                    else
                        predecode_reqtype_s1 = 6'd21;
                    predecode_dcache_load_s1 = 1;
                end
                5'b10000:
                begin
                    if (pcxdecoder_l15_invalidate_cacheline)
                        predecode_reqtype_s1 = 6'd33;
                    else
                        predecode_reqtype_s1 = 6'd2;
                    predecode_icache_bit_s1 = 1;
                end
                5'b00001:
                    if (predecode_is_pcx_config_asi_s1)
                        predecode_reqtype_s1 = 6'd23;
                    else if (predecode_is_pcx_diag_data_access_s1)
                        predecode_reqtype_s1 = 6'd26;
                    else if (predecode_is_pcx_diag_line_flush_s1)
                        predecode_reqtype_s1 = 6'd27;
                    else if (predecode_is_hmc_diag_access_s1)
                        predecode_reqtype_s1 = 6'd30;
                    else if (predecode_is_hmc_flush_s1)
                        predecode_reqtype_s1 = 6'd31;
                    else if (predecode_non_cacheable_s1)
                    begin
                        predecode_reqtype_s1 = 6'd17;
                        
                        
                        
                        predecode_prefetch_bit_s1 = 1'b0;
                    end
                    else
                        predecode_reqtype_s1 = 6'd3;
                
                
                
                
                
                
                
                
                
                
                
                
                5'b00110:
                begin
                    case (pcxdecoder_l15_amo_op)
                    4'b0000:
                    begin
                        predecode_reqtype_s1 = 6'd1;
                    end
                    4'b0001:
                    begin
                        predecode_reqtype_s1 = 6'd35;
                        predecode_atomic_s1 = 1;
                    end
                    4'b0010:
                    begin
                        predecode_reqtype_s1 = 6'd36;
                        predecode_atomic_s1 = 1;
                    end
                    4'b0011:
                    begin
                        predecode_reqtype_s1 = 6'd5;
                        predecode_atomic_s1 = 1;
                    end
                    4'b0100:
                    begin
                        predecode_reqtype_s1 = 6'd38;
                        predecode_atomic_s1 = 1;
                    end
                    4'b0101:
                    begin
                        predecode_reqtype_s1 = 6'd39;
                        predecode_atomic_s1 = 1;
                    end
                    4'b0110:
                    begin
                        predecode_reqtype_s1 = 6'd40;
                        predecode_atomic_s1 = 1;
                    end
                    4'b0111:
                    begin
                        predecode_reqtype_s1 = 6'd41;
                        predecode_atomic_s1 = 1;
                    end
                    4'b1000:
                    begin
                        predecode_reqtype_s1 = 6'd42;
                        predecode_atomic_s1 = 1;
                    end
                    4'b1001:
                    begin
                        predecode_reqtype_s1 = 6'd43;
                        predecode_atomic_s1 = 1;
                    end
                    4'b1010:
                    begin
                        predecode_reqtype_s1 = 6'd44;
                        predecode_atomic_s1 = 1;
                    end
                    4'b1011:
                    begin
                        predecode_reqtype_s1 = 6'd45;
                        predecode_atomic_s1 = 1;
                    end
                    4'b1100:
                    begin
                        predecode_reqtype_s1 = 6'd4;
                        predecode_atomic_s1 = 1;
                    end
                    4'b1101:
                    begin
                        predecode_reqtype_s1 = 6'd1;
                    end
                    endcase
                end
                5'b01001:
                begin
                    predecode_reqtype_s1 = 6'd19;
                    predecode_interrupt_broadcast_s1 = predecode_non_cacheable_s1;
                end
                5'b01010:
                    predecode_reqtype_s1 = 6'd1;
                5'b01011:
                    predecode_reqtype_s1 = 6'd1;
                5'b00100:
                    predecode_reqtype_s1 = 6'd1;
                5'b00101:
                    predecode_reqtype_s1 = 6'd1;
                5'b01101:
                    predecode_reqtype_s1 = 6'd1;
                5'b01110:
                    predecode_reqtype_s1 = 6'd1;
            endcase
        end
    endcase
    predecode_val_s1 = (predecode_source_s1 != 2'd0);
    val_s1 = predecode_val_s1;
    predecode_cache_index_s1[((9-2))-1:0]
         = predecode_address_s1[(((9-2))+4-1):4]; 
    predecode_dtag_write_data_s1[(40 - 4 - ((9-2)))-1:0] = predecode_address_s1[(39):((((9-2))+4-1) + 1)];
    
    
    
    predecode_int_vec_dis_s1 = (pcxdecoder_l15_address[39:32] == constant_int_vec_dis_address[39:32] 
                              && pcxdecoder_l15_address[11:8] == constant_int_vec_dis_address[11:8]); 
    
    predecode_partial_tag_s1[19:4] = pcxdecoder_l15_address[19:4]; 
    predecode_tagcheck_matched_t0ld_s1 = mshr_val_array[0][2'd2] 
                                        && (predecode_partial_tag_s1[19:4] == mshr_ld_address_array[0][19:4]);
    predecode_tagcheck_matched_t1ld_s1 = mshr_val_array[1][2'd2] 
                                        && (predecode_partial_tag_s1[19:4] == mshr_ld_address_array[1][19:4]);
    predecode_tagcheck_matched_t0st_s1 = mshr_val_array[0][2'd3] 
                                        && (pcxdecoder_l15_address[39:4] == mshr_st_address_array[0][39:4]);
    predecode_tagcheck_matched_t1st_s1 = mshr_val_array[1][2'd3] 
                                        && (pcxdecoder_l15_address[39:4] == mshr_st_address_array[1][39:4]);
    predecode_tagcheck_matched_s1 = predecode_tagcheck_matched_t0ld_s1 || predecode_tagcheck_matched_t1ld_s1
                                    || predecode_tagcheck_matched_t0st_s1 || predecode_tagcheck_matched_t1st_s1;
    
    predecode_hit_stbuf_s1 = predecode_tagcheck_matched_t0st_s1 || predecode_tagcheck_matched_t1st_s1;
    predecode_hit_stbuf_threadid_s1 = predecode_tagcheck_matched_t1st_s1 ? 1'b1 : 1'b0;
    
end
reg [3:0] creditman_noc1_avail;
reg [3:0] creditman_noc1_data_avail;
reg [3:0] creditman_noc1_avail_next;
reg [3:0] creditman_noc1_data_avail_next;
reg [3:0] creditman_noc1_reserve;
reg [3:0] creditman_noc1_reserve_next;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        creditman_noc1_avail <= 8;
        creditman_noc1_data_avail <= 2;
        creditman_noc1_reserve <= 0;
    end
    else
    begin
        creditman_noc1_avail <= creditman_noc1_avail_next;
        creditman_noc1_data_avail <= creditman_noc1_data_avail_next;
        creditman_noc1_reserve <= creditman_noc1_reserve_next;
    end
end
reg creditman_noc1_data_add1;
reg creditman_noc1_data_add2;
reg creditman_noc1_data_minus1;
reg creditman_noc1_data_minus2;
reg creditman_noc1_add2;
reg creditman_noc1_add1;
reg creditman_noc1_minus1;
reg creditman_noc1_minus2;
reg creditman_noc1_reserve_add1;
reg creditman_noc1_reserve_minus1;
always @ *
begin
    creditman_noc1_avail_next = creditman_noc1_add2 ? creditman_noc1_avail + 2 :
                             creditman_noc1_add1 ? creditman_noc1_avail + 1 :
                             creditman_noc1_minus1 ? creditman_noc1_avail - 1 :
                             creditman_noc1_minus2 ? creditman_noc1_avail - 2 :
                                                creditman_noc1_avail;
    creditman_noc1_data_avail_next = creditman_noc1_data_add1 ? creditman_noc1_data_avail + 1 :
                                    creditman_noc1_data_add2 ? creditman_noc1_data_avail + 2 :
                                    creditman_noc1_data_minus1 ? creditman_noc1_data_avail - 1 :
                                    creditman_noc1_data_minus2 ? creditman_noc1_data_avail - 2 :
                                                            creditman_noc1_data_avail;
    creditman_noc1_reserve_next = creditman_noc1_reserve_add1 ? creditman_noc1_reserve + 1 :
                                  creditman_noc1_reserve_minus1 ? creditman_noc1_reserve - 1 :
                                                                creditman_noc1_reserve;
end
reg creditman_noc1_mispredicted_s3;
reg creditman_noc1_reserve_s3;
reg creditman_noc1_req;
reg creditman_noc1_upX;
reg creditman_noc1_up1;
reg creditman_noc1_up2;
reg creditman_noc1_down1;
reg creditman_noc1_down2;
reg creditman_noc1_data_up1;
reg creditman_noc1_data_up2;
reg creditman_noc1_data_down1;
reg creditman_noc1_data_down2;
reg decoder_creditman_req_8B_s1;
reg decoder_creditman_req_16B_s1;
reg [1:0] decoder_creditman_noc1_needed;
reg decoder_creditman_noc1_unreserve_s1;
always @ *
begin
    creditman_noc1_req = val_s1 && !stall_s1 && (decoder_creditman_noc1_needed != 2'd0);
    
    
    creditman_noc1_upX = noc1encoder_l15_req_sent || creditman_noc1_mispredicted_s3;
    creditman_noc1_up1 = noc1encoder_l15_req_sent ^ creditman_noc1_mispredicted_s3;
    creditman_noc1_up2 = noc1encoder_l15_req_sent && creditman_noc1_mispredicted_s3;
    creditman_noc1_down1 = creditman_noc1_req && decoder_creditman_noc1_needed == 2'd1;
    creditman_noc1_down2 = creditman_noc1_req && decoder_creditman_noc1_needed == 2'd2;
    creditman_noc1_add2 = creditman_noc1_up2 && ~creditman_noc1_req;
    creditman_noc1_add1 = (creditman_noc1_up2 && creditman_noc1_down1) || (creditman_noc1_up1 && ~creditman_noc1_req);
    creditman_noc1_minus1 = (creditman_noc1_down2 && creditman_noc1_up1) || (creditman_noc1_down1 && !creditman_noc1_upX);
    creditman_noc1_minus2 = creditman_noc1_down2 && !creditman_noc1_upX;
    creditman_noc1_data_up1 = noc1encoder_l15_req_sent && (noc1encoder_l15_req_data_sent == 2'd1);
    
    creditman_noc1_data_up2 = noc1encoder_l15_req_sent && (noc1encoder_l15_req_data_sent == 2'd2);
    creditman_noc1_data_down1 = creditman_noc1_req && decoder_creditman_req_8B_s1;
    creditman_noc1_data_down2 = creditman_noc1_req && decoder_creditman_req_16B_s1;
    creditman_noc1_data_add2 = creditman_noc1_data_up2 && !creditman_noc1_data_down1 && !creditman_noc1_data_down2;
    creditman_noc1_data_add1 = creditman_noc1_data_up1 &&  !creditman_noc1_data_down1 && !creditman_noc1_data_down2 ||
                            creditman_noc1_data_up2 && creditman_noc1_data_down1;
    creditman_noc1_data_minus2 = creditman_noc1_data_down2 && !creditman_noc1_data_up1 && !creditman_noc1_data_up2;
    creditman_noc1_data_minus1 = creditman_noc1_data_down1 &&  !creditman_noc1_data_up1 && !creditman_noc1_data_up2 ||
                            creditman_noc1_data_down2 && creditman_noc1_data_up1;
    creditman_noc1_reserve_add1 = (creditman_noc1_reserve_s3 && !stall_s3 && val_s3) 
                                    && !(val_s1 && !stall_s1 && decoder_creditman_noc1_unreserve_s1);
    creditman_noc1_reserve_minus1 = !(creditman_noc1_reserve_s3 && !stall_s3 && val_s3) 
                                    && (val_s1 && !stall_s1 && decoder_creditman_noc1_unreserve_s1);
end
reg fetch_is_pcx_atomic_instruction_s1;
reg fetch_is_pcx_storenc_instruction_s1;
reg fetch_is_pcx_loadnc_instruction_s1;
reg fetch_is_noc2_data_invalidation_s1;
reg fetch_is_noc2_instruction_invalidation_s1;
reg fetch_is_noc2_ackdt_s1;
reg fetch_is_pcx_flush_s1;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        fetch_state_s1 <= 3'd0;
    end
    else
    begin
        fetch_state_s1 <= fetch_state_next_s1;
    end
end
always @ *
begin
    fetch_is_pcx_atomic_instruction_s1 =
        (predecode_reqtype_s1 == 6'd4 ||
         predecode_reqtype_s1 == 6'd5 ||
         predecode_reqtype_s1 == 6'd35 ||
         predecode_reqtype_s1 == 6'd36 ||
         predecode_reqtype_s1 == 6'd38 ||
         predecode_reqtype_s1 == 6'd39 ||
         predecode_reqtype_s1 == 6'd40 ||
         predecode_reqtype_s1 == 6'd41 ||
         predecode_reqtype_s1 == 6'd42 ||
         predecode_reqtype_s1 == 6'd43 ||
         predecode_reqtype_s1 == 6'd44 ||
         predecode_reqtype_s1 == 6'd45);
    
    fetch_is_pcx_storenc_instruction_s1 = (predecode_reqtype_s1 == 6'd17) && !predecode_int_vec_dis_s1;
    fetch_is_pcx_loadnc_instruction_s1 = (predecode_reqtype_s1 == 6'd15);
    fetch_is_noc2_data_invalidation_s1 = (predecode_reqtype_s1 == 6'd6 ||
                                    predecode_reqtype_s1 == 6'd7);
    fetch_is_noc2_instruction_invalidation_s1 = (predecode_reqtype_s1 == 6'd18);
    fetch_is_noc2_ackdt_s1 = (predecode_reqtype_s1 == 6'd10 || predecode_reqtype_s1 == 6'd11 || predecode_reqtype_s1 == 6'd46);
    fetch_state_next_s1 = 3'd0;
    fetch_is_pcx_flush_s1 = predecode_reqtype_s1 == 6'd27;
    case (fetch_state_s1)
        3'd0:
        begin
            fetch_state_next_s1 = 3'd0;
            if (!stall_s1)
            begin
                
                if ((fetch_is_pcx_atomic_instruction_s1 && (predecode_reqtype_s1 != 6'd36))
                    || fetch_is_pcx_storenc_instruction_s1 || fetch_is_pcx_loadnc_instruction_s1 || fetch_is_pcx_flush_s1)
                    fetch_state_next_s1 = 3'd1;
                else if (fetch_is_noc2_data_invalidation_s1)
                    fetch_state_next_s1 = 3'd2;
                else if (fetch_is_noc2_instruction_invalidation_s1)
                    fetch_state_next_s1 = 3'd6;
                else if (fetch_is_noc2_ackdt_s1)
                    fetch_state_next_s1 = 3'd5;
            end
        end
        3'd1:
        begin
            fetch_state_next_s1 = 3'd1;
            if (!stall_s1)
                fetch_state_next_s1 = 3'd0;
        end
        3'd5:
        begin
            fetch_state_next_s1 = 3'd5;
            if (!stall_s1)
                fetch_state_next_s1 = 3'd0;
        end
        3'd2:
        begin
            fetch_state_next_s1 = 3'd2;
            if (!stall_s1)
                fetch_state_next_s1 = 3'd3;
        end
        3'd3:
        begin
            fetch_state_next_s1 = 3'd3;
            if (!stall_s1)
                fetch_state_next_s1 = 3'd4;
        end
        3'd4:
        begin
            fetch_state_next_s1 = 3'd4;
            if (!stall_s1)
                fetch_state_next_s1 = 3'd0;
        end
        3'd6:
        begin
            fetch_state_next_s1 = 3'd6;
            if (!stall_s1)
                fetch_state_next_s1 = 3'd0;
        end
    endcase
end
reg [2-1:0] decoder_pcx_ack_stage_s1;
reg [2-1:0] decoder_noc2_ack_stage_s1;
reg decoder_stall_on_mshr_allocation_s1;
reg [2-1:0] decoder_mshr_allocation_type_s1;
reg decoder_stall_on_matched_bypassed_index_s1;
reg [2-1:0]decoder_s1_mshr_operation_s1;
reg [2-1:0]decoder_dtag_operation_s1;
reg [1-1:0]decoder_s2_mshr_operation_s1;
reg [1-1:0]decoder_mesi_read_op_s1;
reg [4-1:0]decoder_dcache_operation_s1;
reg [3-1:0]decoder_s3_mshr_operation_s1;
reg [3-1:0]decoder_mesi_write_op_s1;
reg [1-1:0]decoder_wmt_read_op_s1;
reg [3-1:0]decoder_wmt_write_op_s1;
reg [3-1:0]decoder_wmt_compare_op_s1;
reg [3-1:0]decoder_lruarray_write_op_s1;
reg [5-1:0]decoder_cpx_operation_s1;
reg [1-1:0]decoder_hmt_op_s1;
reg [5-1:0]decoder_noc1_operation_s1;
reg [4-1:0]decoder_noc3_operation_s1;
reg [4-1:0]decoder_csm_op_s1;
reg [2-1:0]decoder_config_op_s1;
reg decoder_no_free_mshr_s1;
reg decoder_stall_on_matched_mshr_s1;
reg [2-1:0]decoder_mshrid_s1;
reg decoder_lrsc_flag_read_op_s1;
reg [3-1:0] decoder_lrsc_flag_write_op_s1;
always @ *
begin
    decoder_pcx_ack_stage_s1 = 1'b0;
    decoder_noc2_ack_stage_s1 = 1'b0;
    decoder_stall_on_mshr_allocation_s1 = 1'b0;
    decoder_stall_on_matched_bypassed_index_s1 = 1'b0;
    
    
    decoder_s1_mshr_operation_s1 = 1'b0;
    decoder_dtag_operation_s1 = 1'b0;
    decoder_s2_mshr_operation_s1 = 1'b0;
    decoder_mesi_read_op_s1 = 1'b0;
    decoder_dcache_operation_s1 = 1'b0;
    decoder_s3_mshr_operation_s1 = 1'b0;
    decoder_mesi_write_op_s1 = 1'b0;
    decoder_wmt_read_op_s1 = 1'b0;
    decoder_wmt_write_op_s1 = 1'b0;
    decoder_wmt_compare_op_s1 = 1'b0;
    decoder_lruarray_write_op_s1 = 1'b0;
    decoder_cpx_operation_s1 = 1'b0;
    decoder_noc1_operation_s1 = 1'b0;
    decoder_noc3_operation_s1 = 1'b0;
    decoder_csm_op_s1 = 1'b0;
    decoder_config_op_s1 = 1'b0;
    decoder_creditman_noc1_needed = 2'b0;
    decoder_creditman_noc1_unreserve_s1 = 1'b0;
    decoder_creditman_req_8B_s1 = 1'b0;
    decoder_creditman_req_16B_s1 = 1'b0;
    decoder_stall_on_matched_mshr_s1 = 1'b0;
    decoder_mshr_allocation_type_s1 = 0; 
    decoder_lrsc_flag_read_op_s1 = 1'b0;
    decoder_lrsc_flag_write_op_s1 = 2'b0;
    decoder_no_free_mshr_s1 = 0;
    
    decoder_hmt_op_s1 = 0;
    
    case (predecode_reqtype_s1)
        6'd15:
        begin
            if (fetch_state_s1 == 3'd0)
            begin 
                decoder_stall_on_matched_bypassed_index_s1 = 1;
                decoder_stall_on_matched_mshr_s1 = 1;
                decoder_stall_on_mshr_allocation_s1 = 1'b1;
                decoder_mshr_allocation_type_s1 = 2'd2;
                decoder_dtag_operation_s1 = 2'd1;
                decoder_mesi_read_op_s1 = 1'd1;
                decoder_mesi_write_op_s1 = 3'd3;
                decoder_lrsc_flag_write_op_s1 = 3'd2;
                decoder_wmt_read_op_s1 = 1'd1;
                decoder_wmt_write_op_s1 = 3'd1;
                decoder_wmt_compare_op_s1 = 3'd2;
                decoder_dcache_operation_s1 = 4'd1;
                
                decoder_lruarray_write_op_s1 = 3'd4;
                decoder_cpx_operation_s1 = 5'd1;
                decoder_noc1_operation_s1 = 5'd9;
                decoder_creditman_noc1_needed = 2'd2; 
                decoder_noc3_operation_s1 = 4'd5;
                decoder_csm_op_s1 = 4'd10;
            end
            else
            begin 
                decoder_pcx_ack_stage_s1 = 2'd1;
                decoder_s1_mshr_operation_s1 = 2'd1;
                decoder_mshr_allocation_type_s1 = 2'd2;
                decoder_csm_op_s1 = 4'd1;
                decoder_noc1_operation_s1 = 5'd1;
            end
        end
        6'd16:
        begin
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            decoder_pcx_ack_stage_s1 = 2'd1;
            
            decoder_cpx_operation_s1 = 5'd2;
            
            
        end
        6'd21:
        begin 
            decoder_pcx_ack_stage_s1 = 2'd1;
            decoder_stall_on_matched_bypassed_index_s1 = 1;
            decoder_stall_on_matched_mshr_s1 = 1;
            decoder_stall_on_mshr_allocation_s1 = 1'b1;
            decoder_mshr_allocation_type_s1 = 2'd2;
            decoder_s1_mshr_operation_s1 = 2'd1;
            decoder_dtag_operation_s1 = 2'd1;
            decoder_mesi_read_op_s1 = 1'd1;
            decoder_dcache_operation_s1 = 4'd2;
            decoder_s3_mshr_operation_s1 = 3'd2;
            decoder_cpx_operation_s1 = 5'd4;
            decoder_wmt_read_op_s1 = 1'd1;
            decoder_wmt_write_op_s1 = 3'd4;
            decoder_wmt_compare_op_s1 = 3'd2;
            decoder_csm_op_s1 = 4'd6;
            decoder_lruarray_write_op_s1 = 3'd1;
            decoder_noc1_operation_s1 = 5'd2;
            decoder_creditman_noc1_needed = 2'd1;
        end
        6'd25:
        begin 
            decoder_pcx_ack_stage_s1 = 2'd1;
            decoder_dcache_operation_s1 = 4'd8;
            decoder_cpx_operation_s1 = 5'd16;
        end
        6'd2:
        begin
            decoder_pcx_ack_stage_s1 = 2'd1;
            decoder_stall_on_mshr_allocation_s1 = 1'b1;
            decoder_mshr_allocation_type_s1 = 2'd1;
            decoder_s1_mshr_operation_s1 = 2'd1;
            decoder_csm_op_s1 = 4'd1;
            decoder_noc1_operation_s1 = 5'd3;
            decoder_creditman_noc1_needed = 2'd1;
        end
        6'd17:
        begin
            if (predecode_int_vec_dis_s1)
            begin
                
                
                decoder_pcx_ack_stage_s1 = 2'd3;
                decoder_cpx_operation_s1 = 5'd6;
                decoder_noc1_operation_s1 = 5'd10;
                decoder_creditman_req_8B_s1 = 1'b1;
                decoder_creditman_noc1_needed = 2'd1;
            end
            else
            begin
                if (fetch_state_s1 == 3'd0)
                begin 
                    decoder_stall_on_matched_bypassed_index_s1 = 1;
                    decoder_stall_on_matched_mshr_s1 = 1;
                    decoder_stall_on_mshr_allocation_s1 = 1'b1;
                    decoder_mshr_allocation_type_s1 = 2'd3;
                    decoder_dtag_operation_s1 = 2'd1;
                    decoder_mesi_read_op_s1 = 1'd1;
                    decoder_dcache_operation_s1 = 4'd1;
                    decoder_mesi_write_op_s1 = 3'd3;
                    decoder_lrsc_flag_write_op_s1 = 3'd2;
                    
                    decoder_wmt_read_op_s1 = 1'd1;
                    decoder_wmt_write_op_s1 = 3'd1;
                    decoder_wmt_compare_op_s1 = 3'd2;
                    decoder_lruarray_write_op_s1 = 3'd4;
                    decoder_cpx_operation_s1 = 5'd1;
                    decoder_noc1_operation_s1 = 5'd9;
                    
                    decoder_creditman_noc1_needed = 2'd2; 
                    decoder_noc3_operation_s1 = 4'd5;
                    
                    decoder_creditman_req_8B_s1 = 1'b1;
                    decoder_csm_op_s1 = 4'd10;
                end
                else
                begin 
                    decoder_pcx_ack_stage_s1 = 2'd3;
                    decoder_s1_mshr_operation_s1 = 2'd1;
                    decoder_mshr_allocation_type_s1 = 2'd3;
                    decoder_csm_op_s1 = 4'd1;
                    decoder_noc1_operation_s1 = 5'd5;
                    decoder_s3_mshr_operation_s1 = 3'd6;
                    
                    
                    
                end
            end
        end
        6'd3:
        begin
            if (predecode_hit_stbuf_s1)
            begin 
                decoder_pcx_ack_stage_s1 = 2'd1;
                decoder_stall_on_matched_bypassed_index_s1 = 1'b1;
                decoder_stall_on_mshr_allocation_s1 = 1'b1;
                decoder_mshr_allocation_type_s1 = 2'd3;
                decoder_s1_mshr_operation_s1 = 2'd2;
                decoder_mesi_read_op_s1 = 1'd1;
                decoder_wmt_read_op_s1 = 1'd1;
                decoder_wmt_compare_op_s1 = 3'd4;
                decoder_cpx_operation_s1 = 5'd11;
            end
            else
            begin 
                decoder_pcx_ack_stage_s1 = 2'd1;
                decoder_stall_on_matched_bypassed_index_s1 = 1'b1;
                decoder_stall_on_matched_mshr_s1 = 1'b1;
                decoder_stall_on_mshr_allocation_s1 = 1'b1;
                decoder_s1_mshr_operation_s1 = 2'd1;
                decoder_mshr_allocation_type_s1 = 2'd3;
                decoder_dtag_operation_s1 = 2'd1;
                decoder_mesi_read_op_s1 = 1'd1;
                decoder_s2_mshr_operation_s1 = 1'd1;
                decoder_dcache_operation_s1 = 4'd4;
                decoder_wmt_read_op_s1 = 1'd1;
                decoder_wmt_compare_op_s1 = 3'd2;
                decoder_lruarray_write_op_s1 = 3'd1;
                decoder_csm_op_s1 = 4'd2;
                decoder_s3_mshr_operation_s1 = 3'd3;
                decoder_mesi_write_op_s1 = 3'd2;
                decoder_cpx_operation_s1 = 5'd7;
                decoder_noc1_operation_s1 = 5'd4;
                decoder_creditman_noc1_needed = 2'd1;
            end
        end
        6'd26:
        begin
            
            decoder_pcx_ack_stage_s1 = 2'd2; 
            decoder_dcache_operation_s1 = 4'd9;
            decoder_cpx_operation_s1 = 5'd6;
        end
        6'd27:
        begin
            
            if (fetch_state_s1 == 3'd0)
            begin 
                decoder_stall_on_matched_bypassed_index_s1 = 1;
                decoder_cpx_operation_s1 = 5'd6;
            end
            else
            begin
                decoder_pcx_ack_stage_s1 = 2'd1;
                decoder_dtag_operation_s1 = 2'd1;
                decoder_mesi_read_op_s1 = 1'd1;
                decoder_dcache_operation_s1 = 4'd10;
                decoder_mesi_write_op_s1 = 3'd6;
                decoder_lrsc_flag_write_op_s1 = 3'd4;
                decoder_wmt_read_op_s1 = 1'd1;
                decoder_wmt_write_op_s1 = 3'd5;
                decoder_wmt_compare_op_s1 = 3'd3;
                decoder_lruarray_write_op_s1 = 3'd5;
                decoder_cpx_operation_s1 = 5'd17;
                decoder_noc1_operation_s1 = 5'd12;
                decoder_creditman_noc1_needed = 2'd1;
                decoder_noc3_operation_s1 = 4'd8;
                decoder_csm_op_s1 = 4'd9;
            end
        end
        6'd36: 
        begin
            begin 
            
                decoder_pcx_ack_stage_s1 = 2'd1;
                decoder_stall_on_matched_bypassed_index_s1 = 1'b1;
                decoder_stall_on_matched_mshr_s1 = 1'b1;
                decoder_stall_on_mshr_allocation_s1 = 1'b1;
                decoder_s1_mshr_operation_s1 = 2'd1;
                decoder_mshr_allocation_type_s1 = 2'd3;
                decoder_dtag_operation_s1 = 2'd1;
                decoder_mesi_read_op_s1 = 1'd1;
                decoder_lrsc_flag_read_op_s1 = 1'd1;
                decoder_s2_mshr_operation_s1 = 1'd1;
                decoder_dcache_operation_s1 = 4'd11;
                decoder_wmt_read_op_s1 = 1'd1;
                decoder_wmt_compare_op_s1 = 3'd2;
                decoder_lruarray_write_op_s1 = 3'd6;
                
                decoder_s3_mshr_operation_s1 = 3'd1;  
                
                decoder_lrsc_flag_write_op_s1 = 3'd2;
                decoder_cpx_operation_s1 = 5'd20;
                
                
            end
        end
        6'd4,
        6'd5,
        6'd35,
        6'd38,
        6'd39,
        6'd40,
        6'd41,
        6'd42,
        6'd43,
        6'd44,
        6'd45:
        begin
            if (fetch_state_s1 == 3'd0)
            begin 
                decoder_stall_on_matched_bypassed_index_s1 = 1;
                decoder_stall_on_matched_mshr_s1 = 1;
                decoder_stall_on_mshr_allocation_s1 = 1'b1;
                decoder_mshr_allocation_type_s1 = 2'd2;
                decoder_dtag_operation_s1 = 2'd1;
                decoder_mesi_read_op_s1 = 1'd1;
                decoder_dcache_operation_s1 = 4'd1;
                decoder_mesi_write_op_s1 = 3'd3;
                decoder_lrsc_flag_write_op_s1 = 3'd2;
                
                decoder_wmt_read_op_s1 = 1'd1;
                decoder_wmt_write_op_s1 = 3'd1;
                decoder_wmt_compare_op_s1 = 3'd2;
                decoder_lruarray_write_op_s1 = 3'd4;
                decoder_cpx_operation_s1 = 5'd1;
                decoder_noc1_operation_s1 = 5'd9;
                decoder_creditman_noc1_needed = 2'd2;
                decoder_noc3_operation_s1 = 4'd5;
                decoder_csm_op_s1 = 4'd10;
                
                if (predecode_reqtype_s1 == 6'd4)
                begin
                    decoder_creditman_req_16B_s1 = 1'b1;
                end
                else if (predecode_reqtype_s1 != 6'd35)
                begin
                    
                    decoder_creditman_req_8B_s1 = 1'b1;
                end
            end
            else
            begin
                
                decoder_pcx_ack_stage_s1 = 2'd3;
                decoder_s1_mshr_operation_s1 = 2'd1;
                decoder_mshr_allocation_type_s1 = 2'd2;
                decoder_csm_op_s1 = 4'd1;
                
                
                
                
                
                
                
                
                
                
                case (predecode_reqtype_s1)
                    6'd35:
                    begin
                        decoder_noc1_operation_s1 = 5'd21;
                    end
                    6'd4:
                        decoder_noc1_operation_s1 = 5'd6;
                    6'd5:
                        decoder_noc1_operation_s1 = 5'd7;
                    6'd38:
                        decoder_noc1_operation_s1 = 5'd13;
                    6'd39:
                        decoder_noc1_operation_s1 = 5'd14;
                    6'd40:
                        decoder_noc1_operation_s1 = 5'd15;
                    6'd41:
                        decoder_noc1_operation_s1 = 5'd16;
                    6'd42:
                        decoder_noc1_operation_s1 = 5'd17;
                    6'd43:
                        decoder_noc1_operation_s1 = 5'd18;
                    6'd44:
                        decoder_noc1_operation_s1 = 5'd19;
                    6'd45:
                        decoder_noc1_operation_s1 = 5'd20;
                endcase
                
            end
        end
        6'd18:
        begin
            
            decoder_cpx_operation_s1 = 5'd14;
            if (predecode_is_last_inval_s1)
            begin
                decoder_noc2_ack_stage_s1 = 2'd1;
                decoder_noc3_operation_s1 = 4'd7;
            end
        end
        6'd33:
        begin
            decoder_pcx_ack_stage_s1 = 2'd1;
            decoder_cpx_operation_s1 = 5'd14;
        end
        6'd34:
        begin
            decoder_pcx_ack_stage_s1 = 2'd1;
            decoder_stall_on_matched_bypassed_index_s1 = 1;
            decoder_dtag_operation_s1 = 2'd1;
            decoder_wmt_read_op_s1 = 1'd1;
            decoder_wmt_write_op_s1 = 3'd1;
            
            decoder_wmt_compare_op_s1 = 3'd2; 
            
            decoder_cpx_operation_s1 = 5'd19;
        end 
        6'd6:
        begin
            if (fetch_state_s1 == 3'd0)
            begin 
                decoder_noc2_ack_stage_s1 = 2'd0;
                decoder_stall_on_matched_bypassed_index_s1 = 1;
            end
            else if (fetch_state_s1 == 3'd4)
            begin 
                decoder_noc2_ack_stage_s1 = 2'd1;
                decoder_stall_on_matched_bypassed_index_s1 = 1;
            end
            else
            begin 
                decoder_noc2_ack_stage_s1 = 2'd0;
                decoder_stall_on_matched_bypassed_index_s1 = 1;
            end
            decoder_dtag_operation_s1 = 2'd1;
            decoder_mesi_read_op_s1 = 1'd1;
            decoder_dcache_operation_s1 = 4'd1;
            decoder_s3_mshr_operation_s1 = 3'd4;
            decoder_mesi_write_op_s1 = 3'd3;
            decoder_lrsc_flag_write_op_s1 = 3'd2;
            
            decoder_wmt_read_op_s1 = 1'd1;
            decoder_wmt_write_op_s1 = 3'd1;
            decoder_wmt_compare_op_s1 = 3'd2;
            decoder_lruarray_write_op_s1 = 3'd4;
            decoder_cpx_operation_s1 = 5'd1;
            if (predecode_is_last_inval_s1)
                decoder_noc3_operation_s1 = 4'd1;
            else
                decoder_noc3_operation_s1 = 4'd2;
            decoder_csm_op_s1 = 4'd10;
        end
        6'd7:
        begin
            if (fetch_state_s1 == 3'd0)
            begin 
                decoder_noc2_ack_stage_s1 = 2'd0;
                decoder_stall_on_matched_bypassed_index_s1 = 1;
            end
            else if (fetch_state_s1 == 3'd4)
            begin 
                decoder_noc2_ack_stage_s1 = 2'd1;
                decoder_stall_on_matched_bypassed_index_s1 = 1;
            end
            else
            begin 
                decoder_noc2_ack_stage_s1 = 2'd0;
                decoder_stall_on_matched_bypassed_index_s1 = 1;
            end
            decoder_dtag_operation_s1 = 2'd1;
            decoder_mesi_read_op_s1 = 1'd1;
            decoder_dcache_operation_s1 = 4'd1;
            decoder_mesi_write_op_s1 = 3'd1;
            decoder_lrsc_flag_write_op_s1 = 3'd2;
            if (predecode_is_last_inval_s1)
                decoder_noc3_operation_s1 = 4'd3;
            else
                decoder_noc3_operation_s1 = 4'd4;
        end
        6'd10:
        begin
            if (fetch_state_s1 == 3'd0)
            begin 
                decoder_stall_on_matched_bypassed_index_s1 = 1;
                decoder_dtag_operation_s1 = 2'd1;
                decoder_mesi_read_op_s1 = 1'd1;
                decoder_dcache_operation_s1 = 4'd3;
                decoder_s3_mshr_operation_s1 = 3'd5;
                
                decoder_wmt_read_op_s1 = 1'd1;
                decoder_wmt_write_op_s1 = 3'd2;
                decoder_wmt_compare_op_s1 = 3'd1;
                decoder_lruarray_write_op_s1 = 3'd2;
                decoder_lrsc_flag_write_op_s1 = 3'd3;
                decoder_cpx_operation_s1 = 5'd8;
                decoder_noc1_operation_s1 = 5'd8;
                decoder_creditman_noc1_needed = 2'd1;
                decoder_noc3_operation_s1 = 4'd6;
                decoder_creditman_noc1_unreserve_s1 = 1'b1;
                decoder_csm_op_s1 = 4'd8;
            end
            else 
            begin
                decoder_noc2_ack_stage_s1 = 2'd3;
                decoder_dtag_operation_s1 = 2'd2;
                decoder_dcache_operation_s1 = 4'd5;
                decoder_s3_mshr_operation_s1 = 3'd1;
                decoder_mesi_write_op_s1 = 3'd4;
                
                decoder_wmt_read_op_s1 = 1'd1;
                decoder_wmt_write_op_s1 = 3'd3;
                
                decoder_wmt_compare_op_s1 = 3'd1;
                
                decoder_lruarray_write_op_s1 = 3'd3;
                decoder_cpx_operation_s1 = 5'd5;
                
                decoder_hmt_op_s1 = 1'd1;
                
            end
        end
        6'd8:
        begin
            decoder_noc2_ack_stage_s1 = 2'd3;
            decoder_stall_on_matched_bypassed_index_s1 = 1;
            decoder_s3_mshr_operation_s1 = 3'd1;
            decoder_cpx_operation_s1 = 5'd5;
            
        end
        6'd9:
        begin
            decoder_noc2_ack_stage_s1 = 2'd3;
            decoder_s3_mshr_operation_s1 = 3'd1;
            decoder_cpx_operation_s1 = 5'd9;
        end
        6'd11:
        begin
            if (fetch_state_s1 == 3'd0)
            begin 
                decoder_stall_on_matched_bypassed_index_s1 = 1;
                decoder_dtag_operation_s1 = 2'd1;
                decoder_mesi_read_op_s1 = 1'd1;
                decoder_dcache_operation_s1 = 4'd3;
                decoder_s3_mshr_operation_s1 = 3'd5;
                
                decoder_wmt_read_op_s1 = 1'd1;
                decoder_wmt_write_op_s1 = 3'd2;
                decoder_wmt_compare_op_s1 = 3'd1;
                decoder_lruarray_write_op_s1 = 3'd2;
                decoder_lrsc_flag_write_op_s1 = 3'd3;
                decoder_cpx_operation_s1 = 5'd8;
                decoder_noc1_operation_s1 = 5'd8;
                decoder_creditman_noc1_needed = 2'd1;
                decoder_noc3_operation_s1 = 4'd6;
                decoder_creditman_noc1_unreserve_s1 = 1'b1;
                decoder_csm_op_s1 = 4'd8;
            end
            else 
            begin
                decoder_noc2_ack_stage_s1 = 2'd3;
                decoder_dtag_operation_s1 = 2'd2;
                decoder_s2_mshr_operation_s1 = 1'd1;
                decoder_dcache_operation_s1 = 4'd6;
                decoder_s3_mshr_operation_s1 = 3'd1;
                decoder_mesi_write_op_s1 = 3'd4;
                decoder_lruarray_write_op_s1 = 3'd3;
                decoder_cpx_operation_s1 = 5'd6;
                
                decoder_hmt_op_s1 = 1'd1;
                
            end
        end
        6'd12:
        begin
            decoder_noc2_ack_stage_s1 = 2'd1;
            decoder_stall_on_matched_bypassed_index_s1 = 1;
            decoder_s2_mshr_operation_s1 = 1'd1;
            decoder_dcache_operation_s1 = 4'd7;
            decoder_s3_mshr_operation_s1 = 3'd1;
            decoder_mesi_write_op_s1 = 3'd5;
            decoder_wmt_read_op_s1 = 1'd1;
            decoder_wmt_compare_op_s1 = 3'd4; 
            decoder_cpx_operation_s1 = 5'd11;
            decoder_creditman_noc1_unreserve_s1 = 1'b1;
        end
        6'd13:
        begin
            decoder_noc2_ack_stage_s1 = 2'd1;
            decoder_stall_on_matched_bypassed_index_s1 = 1;
            decoder_s3_mshr_operation_s1 = 3'd1;
            decoder_cpx_operation_s1 = 5'd6;
        end
        6'd32:
        begin
           decoder_noc2_ack_stage_s1 = 2'd1;
           
           
           
        end
        6'd14:
        begin
            decoder_noc2_ack_stage_s1 = 2'd3;
            decoder_stall_on_matched_bypassed_index_s1 = 1;
            decoder_s3_mshr_operation_s1 = 3'd1;
            decoder_cpx_operation_s1 = 5'd10;
        end
        6'd46:
        begin
            if (fetch_state_s1 == 3'd0)
            begin 
                decoder_stall_on_matched_bypassed_index_s1 = 1;
                decoder_dtag_operation_s1 = 2'd1;
                decoder_mesi_read_op_s1 = 1'd1;
                decoder_dcache_operation_s1 = 4'd3;
                decoder_s3_mshr_operation_s1 = 3'd5;
                
                decoder_wmt_read_op_s1 = 1'd1;
                decoder_wmt_write_op_s1 = 3'd2;
                decoder_wmt_compare_op_s1 = 3'd1;
                decoder_lruarray_write_op_s1 = 3'd2;
                decoder_cpx_operation_s1 = 5'd8;
                decoder_noc1_operation_s1 = 5'd8;
                decoder_creditman_noc1_needed = 2'd1;
                decoder_noc3_operation_s1 = 4'd6;
                decoder_creditman_noc1_unreserve_s1 = 1'b1;
                decoder_csm_op_s1 = 4'd8;
            end
            else 
            begin
                decoder_noc2_ack_stage_s1 = 2'd3;
                decoder_dtag_operation_s1 = 2'd2;
                decoder_dcache_operation_s1 = 4'd5;
                decoder_s3_mshr_operation_s1 = 3'd1;
                decoder_mesi_write_op_s1 = 3'd4; 
                decoder_lrsc_flag_write_op_s1 = 3'd1;
                
                decoder_wmt_read_op_s1 = 1'd1;
                
                
   
                
                decoder_wmt_compare_op_s1 = 3'd1;
                decoder_lruarray_write_op_s1 = 3'd3;
                decoder_cpx_operation_s1 = 5'd10;
                
                decoder_hmt_op_s1 = 1'd1;
                
            end
        end
        6'd20:
        begin
            decoder_noc2_ack_stage_s1 = 2'd3;
            decoder_cpx_operation_s1 = 5'd13;
        end
        6'd19:
        begin
            if (predecode_interrupt_broadcast_s1)
            begin
                decoder_pcx_ack_stage_s1 = 2'd1;
                decoder_cpx_operation_s1 = 5'd12;
            end
            else
            begin
                decoder_pcx_ack_stage_s1 = 2'd3;
                decoder_noc1_operation_s1 = 5'd10;
                decoder_creditman_noc1_needed = 2'd1;
                decoder_creditman_req_8B_s1 = 1'b1;
            end
        end
        6'd24:
        begin
            decoder_pcx_ack_stage_s1 = 2'd1;
            decoder_cpx_operation_s1 = 5'd15;
            decoder_config_op_s1 = 2'd1;
        end
        6'd23:
        begin
            decoder_pcx_ack_stage_s1 = 2'd2;
            decoder_cpx_operation_s1 = 5'd6;
            decoder_config_op_s1 = 2'd2;
        end
        6'd28:
        begin
            decoder_noc2_ack_stage_s1 = 2'd2;
            decoder_csm_op_s1 = 4'd3;
            
        end
        6'd29:
        begin
            decoder_pcx_ack_stage_s1 = 2'd1;
            decoder_csm_op_s1 = 4'd5;
            decoder_cpx_operation_s1 = 5'd18;
        end
        6'd30:
        begin
            decoder_pcx_ack_stage_s1 = 2'd2;
            decoder_csm_op_s1 = 4'd4;
            decoder_cpx_operation_s1 = 5'd6;
        end
        6'd31:
        begin
            decoder_pcx_ack_stage_s1 = 2'd1;
            decoder_csm_op_s1 = 4'd7;
            decoder_cpx_operation_s1 = 5'd6;
        end
        6'd1:
        begin 
            decoder_pcx_ack_stage_s1 = 2'd1;
        end
    endcase
    
    decoder_no_free_mshr_s1 = mshr_val_array[predecode_threadid_s1][decoder_mshr_allocation_type_s1];
    decoder_mshrid_s1 =
        (predecode_source_s1 == 2'd2) ? noc2decoder_l15_mshrid : decoder_mshr_allocation_type_s1;
end
reg stall_tag_match_stall_s1;
reg stall_index_bypass_match_s1;
reg stall_index_conflict_stall_s1;
reg stall_mshr_allocation_busy_s1;
reg stall_noc1_data_buffer_unavail_s1;
reg stall_noc1_command_buffer_1_unavail_s1;
reg stall_noc1_command_buffer_2_unavail_s1;
reg stall_noc1_command_buffer_unavail_s1;
reg stall_pcx_noc1_buffer_s1;
reg [4:0] stall_tmp_operand1;
reg [4:0] stall_tmp_operand2;
reg [4:0] stall_tmp_result;
always @ *
begin
    
    stall_noc1_data_buffer_unavail_s1 = decoder_creditman_req_8B_s1  ? creditman_noc1_data_avail == 4'd0 :
                                                    decoder_creditman_req_16B_s1 ? creditman_noc1_data_avail < 4'd2 :
                                                                                            1'b0;
    
    
    
    
    stall_tmp_operand1 = {1'b1, creditman_noc1_avail[3:0]};
    stall_tmp_operand2 = {1'b0, creditman_noc1_reserve[3:0]};
    stall_tmp_result = stall_tmp_operand1 - stall_tmp_operand2;
    stall_noc1_command_buffer_1_unavail_s1 = (stall_tmp_result[3:0] == 4'b0) || stall_tmp_result[4] == 1'b0;
    stall_noc1_command_buffer_2_unavail_s1 = stall_noc1_command_buffer_1_unavail_s1 || (stall_tmp_result[3:0] == 4'b1);
    stall_noc1_command_buffer_unavail_s1 = (decoder_creditman_noc1_needed == 2'd1 && stall_noc1_command_buffer_1_unavail_s1)
                                        || (decoder_creditman_noc1_needed == 2'd2 && stall_noc1_command_buffer_2_unavail_s1);
    
    stall_pcx_noc1_buffer_s1 = (stall_noc1_command_buffer_unavail_s1 || stall_noc1_data_buffer_unavail_s1)
                                            && (predecode_source_s1 == 2'd1)
                                            && (fetch_state_s1 == 3'd0);
    
    stall_tag_match_stall_s1 = predecode_tagcheck_matched_s1 && decoder_stall_on_matched_mshr_s1;
    
    stall_index_bypass_match_s1 = (val_s2 && (predecode_cache_index_s1 == cache_index_s2))
                                     || (val_s3 && (predecode_cache_index_s1 == cache_index_s3));
    stall_index_conflict_stall_s1 = decoder_stall_on_matched_bypassed_index_s1 && stall_index_bypass_match_s1;
    stall_mshr_allocation_busy_s1 = decoder_no_free_mshr_s1 && decoder_stall_on_mshr_allocation_s1;
    
    stall_s1 = val_s1 && (stall_tag_match_stall_s1 || stall_index_conflict_stall_s1 || stall_s2 || stall_mshr_allocation_busy_s1
                    || stall_pcx_noc1_buffer_s1);
end
reg dtag_val_s1;
reg dtag_rw_s1;
reg [((9-2))-1:0] dtag_index_s1;
reg [2-1:0] dtag_write_way_s1;
reg [33-1:0] dtag_write_tag_s1;
reg [3:0] dtag_write_way_mask;
always @ *
begin
    dtag_val_s1 = 0;
    dtag_rw_s1 = 0;
    dtag_index_s1 = 0;
    dtag_write_way_s1 = 0;
    dtag_write_tag_s1[33-1:0]  = 0;
    dtag_write_way_mask = 0;
    case (decoder_dtag_operation_s1)
        2'd1:
        begin
            dtag_val_s1 = val_s1;
            dtag_rw_s1 = 1'b1;
            dtag_index_s1 = predecode_cache_index_s1;
        end
        2'd2:
        begin
            dtag_val_s1 = val_s1;
            dtag_rw_s1 = 1'b0;
            dtag_index_s1 = predecode_cache_index_s1;
            dtag_write_way_s1 = lru_way_s2; 
            
            dtag_write_tag_s1[33-1:0]  = {{33-(40 - 4 - ((9-2))){1'b0}},predecode_dtag_write_data_s1[(40 - 4 - ((9-2)))-1:0]} ;
        end
    endcase
    dtag_write_way_mask = (dtag_write_way_s1 == 2'b00) ? 4'b0_0_0_1 :
                            (dtag_write_way_s1 == 2'b01) ? 4'b0_0_1_0 :
                            (dtag_write_way_s1 == 2'b10) ? 4'b0_1_0_0 :
                                                        4'b1_0_0_0 ;
    
    l15_dtag_val_s1 = dtag_val_s1 && !stall_s1;
    l15_dtag_rw_s1 = dtag_rw_s1;
    l15_dtag_index_s1[((9-2))-1:0] = dtag_index_s1;
    l15_dtag_write_data_s1[33*4-1:0] = {4{dtag_write_tag_s1[33-1:0]}} ;
    l15_dtag_write_mask_s1[33*4-1:0] =
                                                                    {{33{dtag_write_way_mask[3]}},
                                                                     {33{dtag_write_way_mask[2]}},
                                                                     {33{dtag_write_way_mask[1]}},
                                                                     {33{dtag_write_way_mask[0]}}};
end
reg mesi_read_val_s1;
reg [((9-2))-1:0] mesi_read_index_s1;
always @ *
begin
    mesi_read_val_s1 = 0;
    mesi_read_index_s1 = 0;
    case (decoder_mesi_read_op_s1)
        1'd1:
        begin
            mesi_read_val_s1 = 1'b1;
            mesi_read_index_s1 = predecode_cache_index_s1;
        end
    endcase
    l15_mesi_read_val_s1 = mesi_read_val_s1 && val_s1 && !stall_s1;
    l15_mesi_read_index_s1[((9-2))-1:0] = mesi_read_index_s1;
end
reg lrsc_flag_read_val_s1;
reg [((9-2))-1:0] lrsc_flag_read_index_s1;
always @ *
begin
    lrsc_flag_read_val_s1 = 0;
    lrsc_flag_read_index_s1 = 0;
    case (decoder_lrsc_flag_read_op_s1)
        1'd1:
        begin
            lrsc_flag_read_val_s1 = 1'b1;
            lrsc_flag_read_index_s1 = predecode_cache_index_s1;
        end
    endcase
    l15_lrsc_flag_read_val_s1 = lrsc_flag_read_val_s1 && val_s1 && !stall_s1;
    l15_lrsc_flag_read_index_s1[((9-2))-1:0] = lrsc_flag_read_index_s1;
end
reg [((((((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) + 1) + 1) + 1)-1:0] mshr_control_bits_write_s1;
always @ *
begin
    
    
    mshr_control_bits_write_s1 = 0;
    mshr_control_bits_write_s1 [(((((0 + 1) + 1) + 1) + 1) + 3) -: 3] = predecode_size_s1;
    mshr_control_bits_write_s1 [((((((0 + 1) + 1) + 1) + 1) + 3) + 1) -: 1] = predecode_threadid_s1;
    mshr_control_bits_write_s1 [(((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) -: 2] = predecode_l1_replacement_way_s1;
    
    mshr_control_bits_write_s1 [((((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) + 1) -: 1] = (predecode_reqtype_s1 == 6'd35) ? 1'b0 : predecode_non_cacheable_s1;
    mshr_control_bits_write_s1 [(((((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) + 1) + 1) -: 1] = predecode_blockstore_bit_s1;
    mshr_control_bits_write_s1 [(0 + 1) -: 1] = predecode_blockstore_init_s1;
    mshr_control_bits_write_s1 [0 -: 1] = predecode_prefetch_bit_s1;
    
    mshr_control_bits_write_s1 [((((0 + 1) + 1) + 1) + 1) -: 1] = predecode_icache_bit_s1;
    mshr_control_bits_write_s1 [((0 + 1) + 1) -: 1] = predecode_dcache_load_s1;
    mshr_control_bits_write_s1 [(((0 + 1) + 1) + 1) -: 1] = predecode_atomic_s1;
end
reg s1_mshr_write_val_s1;
reg [3-1:0] s1_mshr_write_type_s1;
reg [39:0] s1_mshr_write_address_s1;
reg [((((((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) + 1) + 1) + 1)-1:0] s1_mshr_write_control_s1;
reg [2-1:0] s1_mshr_write_mshrid_s1;
reg [0:0] s1_mshr_write_threadid_s1;
reg [15:0] unshifted_write_mask_s1;
reg [15:0] write_mask_s1;
reg [15:0] write_mask_1B_s1;
reg [15:0] write_mask_2B_s1;
reg [15:0] write_mask_4B_s1;
reg [15:0] write_mask_8B_s1;
reg [15:0] write_mask_16B_s1;
always @ *
begin
    s1_mshr_write_val_s1 = 0;
    s1_mshr_write_type_s1 = 0;
    s1_mshr_write_address_s1 = 0;
    s1_mshr_write_control_s1 = 0;
    s1_mshr_write_mshrid_s1 = 0;
    
    
    write_mask_s1 = 0;
    s1_mshr_write_threadid_s1 = 0;
    case (decoder_s1_mshr_operation_s1)
        2'd1:
        begin
            s1_mshr_write_val_s1 = 1'b1; 
            s1_mshr_write_type_s1 = 3'b001;
            s1_mshr_write_address_s1 = pcxdecoder_l15_address;
            s1_mshr_write_control_s1 = mshr_control_bits_write_s1;
            s1_mshr_write_mshrid_s1 = decoder_mshr_allocation_type_s1;
            s1_mshr_write_threadid_s1[0:0] = predecode_threadid_s1[0:0];
        end
        2'd2:
        begin
            s1_mshr_write_val_s1 = 1'b1;
            s1_mshr_write_type_s1 = 3'b100;
            
            s1_mshr_write_threadid_s1 = predecode_hit_stbuf_threadid_s1;
        end
    endcase
    unshifted_write_mask_s1 =   (predecode_size_s1 == 3'b001) ? 16'b1000_0000_0000_0000 :
                                (predecode_size_s1 == 3'b010) ? 16'b1100_0000_0000_0000 :
                                (predecode_size_s1 == 3'b011) ? 16'b1111_0000_0000_0000 :
                                                                    16'b1111_1111_0000_0000 ;
    write_mask_1B_s1 = unshifted_write_mask_s1 >> (pcxdecoder_l15_address & 4'b1111);
    write_mask_2B_s1 = unshifted_write_mask_s1 >> (pcxdecoder_l15_address & 4'b1110);
    write_mask_4B_s1 = unshifted_write_mask_s1 >> (pcxdecoder_l15_address & 4'b1100);
    write_mask_8B_s1 = unshifted_write_mask_s1 >> (pcxdecoder_l15_address & 4'b1000);
    write_mask_16B_s1 = {16{1'b1}};
    case(predecode_size_s1)
        3'b001:
        begin
            write_mask_s1 = write_mask_1B_s1;
        end
        3'b010:
        begin
            write_mask_s1 = write_mask_2B_s1;
        end
        3'b011:
        begin
            write_mask_s1 = write_mask_4B_s1;
        end
        3'b100:
        begin
            write_mask_s1 = write_mask_8B_s1;
        end
        3'b101:
        begin
            write_mask_s1 = write_mask_16B_s1;
        end
        default:
        begin
            write_mask_s1 = write_mask_16B_s1;
        end
    endcase
    
    pipe_mshr_writereq_val_s1 = s1_mshr_write_val_s1 && !stall_s1 && val_s1;
    pipe_mshr_writereq_op_s1[3-1:0] = s1_mshr_write_type_s1[3-1:0];
    pipe_mshr_writereq_address_s1[39:0] = s1_mshr_write_address_s1[39:0];
    pipe_mshr_writereq_control_s1[((((((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) + 1) + 1) + 1)-1:0] = s1_mshr_write_control_s1[((((((((((0 + 1) + 1) + 1) + 1) + 3) + 1) + 2) + 1) + 1) + 1)-1:0];
    pipe_mshr_writereq_write_buffer_data_s1[127:0] = {pcxdecoder_l15_data, pcxdecoder_l15_data};
    pipe_mshr_writereq_write_buffer_byte_mask_s1[15:0] = write_mask_s1[15:0];
    pipe_mshr_writereq_mshrid_s1[2-1:0] = s1_mshr_write_mshrid_s1[2-1:0];
    pipe_mshr_writereq_threadid_s1 = s1_mshr_write_threadid_s1;
end
always @ *
begin
    l15_lruarray_read_val_s1 = val_s1 && !stall_s1;
    l15_lruarray_read_index_s1 = predecode_cache_index_s1;
end
reg acklogic_pcx_s1;
reg acklogic_noc2_s1;
always @ *
begin
    acklogic_pcx_s1 = 0;
    acklogic_noc2_s1 = 0;
    if (decoder_pcx_ack_stage_s1 == 2'd1)
        acklogic_pcx_s1 = 1;
    if (decoder_noc2_ack_stage_s1 == 2'd1)
        acklogic_noc2_s1 = 1;
    
    pcx_ack_s1 = val_s1 && !stall_s1 && acklogic_pcx_s1;
    noc2_ack_s1 = val_s1 && !stall_s1 && acklogic_noc2_s1;
    
    
    l15_pcxdecoder_header_ack = (predecode_source_s1 == 2'd1) && !stall_s1 && val_s1
                                                && (fetch_state_s1 == 3'd0);
    
    l15_noc2decoder_header_ack = (predecode_source_s1 == 2'd2) && !stall_s1 && val_s1
                                                && (fetch_state_s1 == 3'd0);
end
reg val_s2_next;
reg [1-1:0] threadid_s2;
reg [1-1:0] threadid_s2_next;
reg [2-1:0] mshrid_s2;
reg [2-1:0] mshrid_s2_next;
reg [40-1:0] address_s2;
reg [40-1:0] address_s2_next;
reg [1-1:0] non_cacheable_s2;
reg [1-1:0] non_cacheable_s2_next;
reg [3-1:0] size_s2;
reg [3-1:0] size_s2_next;
reg [1-1:0] prefetch_s2;
reg [1-1:0] prefetch_s2_next;
reg [2-1:0] l1_replacement_way_s2;
reg [2-1:0] l1_replacement_way_s2_next;
reg [1-1:0] l2_miss_s2;
reg [1-1:0] l2_miss_s2_next;
reg [1-1:0] f4b_s2;
reg [1-1:0] f4b_s2_next;
reg [1-1:0] predecode_noc2_inval_s2;
reg [1-1:0] predecode_noc2_inval_s2_next;
reg [4-1:0] predecode_fwd_subcacheline_vector_s2;
reg [4-1:0] predecode_fwd_subcacheline_vector_s2_next;
reg [3-1:0] lrsc_flag_write_op_s2;
reg [3-1:0] lrsc_flag_write_op_s2_next;
reg [1-1:0] blockstore_s2;
reg [1-1:0] blockstore_s2_next;
reg [1-1:0] blockstoreinit_s2;
reg [1-1:0] blockstoreinit_s2_next;
reg [6-1:0] predecode_reqtype_s2;
reg [6-1:0] predecode_reqtype_s2_next;
reg [2-1:0] decoder_dtag_operation_s2;
reg [2-1:0] decoder_dtag_operation_s2_next;
reg [3-1:0] wmt_write_op_s2;
reg [3-1:0] wmt_write_op_s2_next;
reg [3-1:0] wmt_compare_op_s2;
reg [3-1:0] wmt_compare_op_s2_next;
reg [3-1:0] lruarray_write_op_s2;
reg [3-1:0] lruarray_write_op_s2_next;
reg [4-1:0] csm_op_s2;
reg [4-1:0] csm_op_s2_next;
reg [2-1:0] config_op_s2;
reg [2-1:0] config_op_s2_next;
reg [1-1:0] wmt_read_op_s2;
reg [1-1:0] wmt_read_op_s2_next;
reg [(14+8+8)-1:0] noc2_src_homeid_s2;
reg [(14+8+8)-1:0] noc2_src_homeid_s2_next;
reg [(14+8+8)-1:0] hmt_fill_homeid_s2;
reg [(14+8+8)-1:0] hmt_fill_homeid_s2_next;
reg [3-1:0] s3_mshr_operation_s2;
reg [3-1:0] s3_mshr_operation_s2_next;
reg [5-1:0] cpx_operation_s2;
reg [5-1:0] cpx_operation_s2_next;
reg [5-1:0] noc1_operation_s2;
reg [5-1:0] noc1_operation_s2_next;
reg [4-1:0] noc3_operations_s2;
reg [4-1:0] noc3_operations_s2_next;
reg [1-1:0] mesi_read_op_s2;
reg [1-1:0] mesi_read_op_s2_next;
reg [3-1:0] mesi_write_op_s2;
reg [3-1:0] mesi_write_op_s2_next;
reg [4-1:0] dcache_operation_s2;
reg [4-1:0] dcache_operation_s2_next;
reg [1-1:0] s2_mshr_operation_s2;
reg [1-1:0] s2_mshr_operation_s2_next;
reg [2-1:0] pcx_ack_stage_s2;
reg [2-1:0] pcx_ack_stage_s2_next;
reg [2-1:0] noc2_ack_stage_s2;
reg [2-1:0] noc2_ack_stage_s2_next;
reg [2-1:0] noc2_ack_state_s2;
reg [2-1:0] noc2_ack_state_s2_next;
reg [33-1:0] csm_pcx_data_s2;
reg [33-1:0] csm_pcx_data_s2_next;
reg [33-1:0] hmt_op_s2;
reg [33-1:0] hmt_op_s2_next;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        val_s2 <= 1'b0;
        threadid_s2 <= 0;
mshrid_s2 <= 0;
address_s2 <= 0;
non_cacheable_s2 <= 0;
size_s2 <= 0;
prefetch_s2 <= 0;
l1_replacement_way_s2 <= 0;
l2_miss_s2 <= 0;
f4b_s2 <= 0;
predecode_noc2_inval_s2 <= 0;
predecode_fwd_subcacheline_vector_s2 <= 0;
lrsc_flag_write_op_s2 <= 0;
blockstore_s2 <= 0;
blockstoreinit_s2 <= 0;
predecode_reqtype_s2 <= 0;
decoder_dtag_operation_s2 <= 0;
wmt_write_op_s2 <= 0;
wmt_compare_op_s2 <= 0;
lruarray_write_op_s2 <= 0;
csm_op_s2 <= 0;
config_op_s2 <= 0;
wmt_read_op_s2 <= 0;
noc2_src_homeid_s2 <= 0;
hmt_fill_homeid_s2 <= 0;
s3_mshr_operation_s2 <= 0;
cpx_operation_s2 <= 0;
noc1_operation_s2 <= 0;
noc3_operations_s2 <= 0;
mesi_read_op_s2 <= 0;
mesi_write_op_s2 <= 0;
dcache_operation_s2 <= 0;
s2_mshr_operation_s2 <= 0;
pcx_ack_stage_s2 <= 0;
noc2_ack_stage_s2 <= 0;
noc2_ack_state_s2 <= 0;
csm_pcx_data_s2 <= 0;
hmt_op_s2 <= 0;
    end
    else
    begin
        val_s2 <= val_s2_next;
        threadid_s2 <= threadid_s2_next;
mshrid_s2 <= mshrid_s2_next;
address_s2 <= address_s2_next;
non_cacheable_s2 <= non_cacheable_s2_next;
size_s2 <= size_s2_next;
prefetch_s2 <= prefetch_s2_next;
l1_replacement_way_s2 <= l1_replacement_way_s2_next;
l2_miss_s2 <= l2_miss_s2_next;
f4b_s2 <= f4b_s2_next;
predecode_noc2_inval_s2 <= predecode_noc2_inval_s2_next;
predecode_fwd_subcacheline_vector_s2 <= predecode_fwd_subcacheline_vector_s2_next;
lrsc_flag_write_op_s2 <= lrsc_flag_write_op_s2_next;
blockstore_s2 <= blockstore_s2_next;
blockstoreinit_s2 <= blockstoreinit_s2_next;
predecode_reqtype_s2 <= predecode_reqtype_s2_next;
decoder_dtag_operation_s2 <= decoder_dtag_operation_s2_next;
wmt_write_op_s2 <= wmt_write_op_s2_next;
wmt_compare_op_s2 <= wmt_compare_op_s2_next;
lruarray_write_op_s2 <= lruarray_write_op_s2_next;
csm_op_s2 <= csm_op_s2_next;
config_op_s2 <= config_op_s2_next;
wmt_read_op_s2 <= wmt_read_op_s2_next;
noc2_src_homeid_s2 <= noc2_src_homeid_s2_next;
hmt_fill_homeid_s2 <= hmt_fill_homeid_s2_next;
s3_mshr_operation_s2 <= s3_mshr_operation_s2_next;
cpx_operation_s2 <= cpx_operation_s2_next;
noc1_operation_s2 <= noc1_operation_s2_next;
noc3_operations_s2 <= noc3_operations_s2_next;
mesi_read_op_s2 <= mesi_read_op_s2_next;
mesi_write_op_s2 <= mesi_write_op_s2_next;
dcache_operation_s2 <= dcache_operation_s2_next;
s2_mshr_operation_s2 <= s2_mshr_operation_s2_next;
pcx_ack_stage_s2 <= pcx_ack_stage_s2_next;
noc2_ack_stage_s2 <= noc2_ack_stage_s2_next;
noc2_ack_state_s2 <= noc2_ack_state_s2_next;
csm_pcx_data_s2 <= csm_pcx_data_s2_next;
hmt_op_s2 <= hmt_op_s2_next;
    end
end
reg [1:0] way_mshr_st_s2;
reg [(40 - 4 - ((9-2)))-1:0] address_cache_tag_s2;
always @ *
begin
    cache_index_s2 = address_s2[(((9-2))+4-1):4];
    cache_index_l1d_s2 = address_s2[(6 + 4):4];
    address_cache_tag_s2 = address_s2[(39):((((9-2))+4-1) + 1)];
    way_mshr_st_s2 = mshr_st_way_array[threadid_s2];
    
    if (stall_s2)
    begin
        val_s2_next = val_s2;
        
        threadid_s2_next = threadid_s2;
mshrid_s2_next = mshrid_s2;
address_s2_next = address_s2;
non_cacheable_s2_next = non_cacheable_s2;
size_s2_next = size_s2;
prefetch_s2_next = prefetch_s2;
l1_replacement_way_s2_next = l1_replacement_way_s2;
l2_miss_s2_next = l2_miss_s2;
f4b_s2_next = f4b_s2;
predecode_noc2_inval_s2_next = predecode_noc2_inval_s2;
predecode_fwd_subcacheline_vector_s2_next = predecode_fwd_subcacheline_vector_s2;
lrsc_flag_write_op_s2_next = lrsc_flag_write_op_s2;
blockstore_s2_next = blockstore_s2;
blockstoreinit_s2_next = blockstoreinit_s2;
predecode_reqtype_s2_next = predecode_reqtype_s2;
decoder_dtag_operation_s2_next = decoder_dtag_operation_s2;
wmt_write_op_s2_next = wmt_write_op_s2;
wmt_compare_op_s2_next = wmt_compare_op_s2;
lruarray_write_op_s2_next = lruarray_write_op_s2;
csm_op_s2_next = csm_op_s2;
config_op_s2_next = config_op_s2;
wmt_read_op_s2_next = wmt_read_op_s2;
noc2_src_homeid_s2_next = noc2_src_homeid_s2;
hmt_fill_homeid_s2_next = hmt_fill_homeid_s2;
s3_mshr_operation_s2_next = s3_mshr_operation_s2;
cpx_operation_s2_next = cpx_operation_s2;
noc1_operation_s2_next = noc1_operation_s2;
noc3_operations_s2_next = noc3_operations_s2;
mesi_read_op_s2_next = mesi_read_op_s2;
mesi_write_op_s2_next = mesi_write_op_s2;
dcache_operation_s2_next = dcache_operation_s2;
s2_mshr_operation_s2_next = s2_mshr_operation_s2;
pcx_ack_stage_s2_next = pcx_ack_stage_s2;
noc2_ack_stage_s2_next = noc2_ack_stage_s2;
noc2_ack_state_s2_next = noc2_ack_state_s2;
csm_pcx_data_s2_next = csm_pcx_data_s2;
hmt_op_s2_next = hmt_op_s2;
        
        
    end
    else
    begin
        val_s2_next = val_s1 && !stall_s1;
        threadid_s2_next = predecode_threadid_s1;
        mshrid_s2_next = decoder_mshrid_s1;
        address_s2_next = predecode_address_s1;
        non_cacheable_s2_next = predecode_non_cacheable_s1;
        size_s2_next = predecode_size_s1;
        prefetch_s2_next = predecode_prefetch_bit_s1;
        l1_replacement_way_s2_next = predecode_l1_replacement_way_s1;
        l2_miss_s2_next = predecode_l2_miss_s1;
        f4b_s2_next = predecode_f4b_s1;
        
        wmt_write_op_s2_next = decoder_wmt_write_op_s1;
        wmt_compare_op_s2_next = decoder_wmt_compare_op_s1;
        lruarray_write_op_s2_next = decoder_lruarray_write_op_s1;
        csm_op_s2_next = decoder_csm_op_s1;
        config_op_s2_next = decoder_config_op_s1;
        s3_mshr_operation_s2_next = decoder_s3_mshr_operation_s1;
        cpx_operation_s2_next = decoder_cpx_operation_s1;
        noc1_operation_s2_next = decoder_noc1_operation_s1;
        noc3_operations_s2_next = decoder_noc3_operation_s1;
        mesi_read_op_s2_next = decoder_mesi_read_op_s1;
        mesi_write_op_s2_next = decoder_mesi_write_op_s1;
        dcache_operation_s2_next = decoder_dcache_operation_s1;
        s2_mshr_operation_s2_next = decoder_s2_mshr_operation_s1;
        pcx_ack_stage_s2_next = decoder_pcx_ack_stage_s1;
        noc2_ack_stage_s2_next = decoder_noc2_ack_stage_s1;
        noc2_ack_state_s2_next = noc2decoder_l15_ack_state;
        predecode_reqtype_s2_next = predecode_reqtype_s1;
        predecode_fwd_subcacheline_vector_s2_next = predecode_fwd_subcacheline_vector_s1;
        predecode_noc2_inval_s2_next = predecode_noc2_inval_s1;
        blockstore_s2_next = predecode_blockstore_bit_s1;
        blockstoreinit_s2_next = predecode_blockstore_init_s1;
        noc2_src_homeid_s2_next = noc2decoder_l15_src_homeid;
        lrsc_flag_write_op_s2_next = decoder_lrsc_flag_write_op_s1;
        
        hmt_fill_homeid_s2_next = predecode_mshr_read_homeid_s1;
        
        csm_pcx_data_s2_next = pcxdecoder_l15_csm_data;
        decoder_dtag_operation_s2_next = decoder_dtag_operation_s1;
        wmt_read_op_s2_next = decoder_wmt_read_op_s1;
        
        hmt_op_s2_next = decoder_hmt_op_s1;
        
    end
end
always @ *
begin
    
    
    stall_s2 = val_s2 && stall_s3;
end
always @ *
begin
    
    
    pcx_ack_s2 = val_s2 && !stall_s2 && (pcx_ack_stage_s2 == 2'd2);
    noc2_ack_s2 = val_s2 && !stall_s2 && (noc2_ack_stage_s2 == 2'd2);
end
reg [33-1:0] dtag_tag_way0_s2;
reg [33-1:0] dtag_tag_way1_s2;
reg [33-1:0] dtag_tag_way2_s2;
reg [33-1:0] dtag_tag_way3_s2;
reg [2-1:0] mesi_state_way0_s2;
reg [2-1:0] mesi_state_way1_s2;
reg [2-1:0] mesi_state_way2_s2;
reg [2-1:0] mesi_state_way3_s2;
reg [7:0] mesi_read_data_s2;
reg tagcheck_way0_equals;
reg tagcheck_way1_equals;
reg tagcheck_way2_equals;
reg tagcheck_way3_equals;
reg [1:0] tagcheck_state_s2;
reg tagcheck_state_me_s2;
reg tagcheck_state_mes_s2;
reg tagcheck_state_s_s2;
reg tagcheck_state_m_s2;
reg tagcheck_state_e_s2;
reg [1:0] tagcheck_way_s2;
reg tagcheck_val_s2;
reg tagcheck_lrsc_flag_s2;
reg [1:0] lru_state_s2;
reg lru_state_m_s2;
reg lru_state_mes_s2;
reg [(40 - 4 - ((9-2)))-1:0] lru_way_tag_s2;
reg [39:0] lru_way_address_s2;
reg [1:0] flush_state_s2;
reg flush_state_m_s2;
reg flush_state_me_s2;
reg flush_state_mes_s2;
reg [1:0] flush_way_s2;
reg [(40 - 4 - ((9-2)))-1:0] flush_way_tag_s2;
reg [39:0] flush_way_address_s2;
always @ *
begin
    
    dtag_tag_way0_s2 = dtag_l15_dout_s2[0*33 +: 33];
    dtag_tag_way1_s2 = dtag_l15_dout_s2[1*33 +: 33];
    dtag_tag_way2_s2 = dtag_l15_dout_s2[2*33 +: 33];
    dtag_tag_way3_s2 = dtag_l15_dout_s2[3*33 +: 33];
    mesi_state_way0_s2 = mesi_l15_dout_s2[1:0];
    mesi_state_way1_s2 = mesi_l15_dout_s2[3:2];
    mesi_state_way2_s2 = mesi_l15_dout_s2[5:4];
    mesi_state_way3_s2 = mesi_l15_dout_s2[7:6];
    mesi_read_data_s2 = mesi_l15_dout_s2;
    
    lru_state_s2 =   (lru_way_s2 == 0) ? mesi_state_way0_s2 :
                        (lru_way_s2 == 1) ? mesi_state_way1_s2 :
                        (lru_way_s2 == 2) ? mesi_state_way2_s2 :
                                                mesi_state_way3_s2;
    lru_way_tag_s2[(40 - 4 - ((9-2)))-1:0] =
                        (lru_way_s2 == 0) ? dtag_tag_way0_s2[(40 - 4 - ((9-2)))-1:0] :
                        (lru_way_s2 == 1) ? dtag_tag_way1_s2[(40 - 4 - ((9-2)))-1:0] :
                        (lru_way_s2 == 2) ? dtag_tag_way2_s2[(40 - 4 - ((9-2)))-1:0] :
                                                dtag_tag_way3_s2[(40 - 4 - ((9-2)))-1:0];
    lru_way_address_s2 = {lru_way_tag_s2, address_s2[(((9-2))+4-1):4], 4'b0};
    
    
    tagcheck_way0_equals = (address_cache_tag_s2[(40 - 4 - ((9-2)))-1:0] == dtag_tag_way0_s2[(40 - 4 - ((9-2)))-1:0]);
    tagcheck_way1_equals = (address_cache_tag_s2[(40 - 4 - ((9-2)))-1:0] == dtag_tag_way1_s2[(40 - 4 - ((9-2)))-1:0]);
    tagcheck_way2_equals = (address_cache_tag_s2[(40 - 4 - ((9-2)))-1:0] == dtag_tag_way2_s2[(40 - 4 - ((9-2)))-1:0]);
    tagcheck_way3_equals = (address_cache_tag_s2[(40 - 4 - ((9-2)))-1:0] == dtag_tag_way3_s2[(40 - 4 - ((9-2)))-1:0]);
    {tagcheck_val_s2, tagcheck_way_s2} = tagcheck_way0_equals && (mesi_state_way0_s2 != 2'd0) ? {1'b1, 2'd0} :
                                                    tagcheck_way1_equals && (mesi_state_way1_s2 != 2'd0) ?  {1'b1, 2'd1} :
                                                    tagcheck_way2_equals && (mesi_state_way2_s2 != 2'd0) ?  {1'b1, 2'd2} :
                                                    tagcheck_way3_equals && (mesi_state_way3_s2 != 2'd0) ?  {1'b1, 2'd3} : 3'b0;
    
    
    
    
    tagcheck_lrsc_flag_s2 = (tagcheck_val_s2 == 1'b0) ? 1'b0 :
                                (tagcheck_way_s2 == 2'd0) ? lrsc_flag_l15_dout_s2[0] :
                                (tagcheck_way_s2 == 2'd1) ? lrsc_flag_l15_dout_s2[1] :
                                (tagcheck_way_s2 == 2'd2) ? lrsc_flag_l15_dout_s2[2] :
                                                            lrsc_flag_l15_dout_s2[3] ;
    tagcheck_state_s2 = (tagcheck_val_s2 == 1'b0) ? 2'd0 :
                                (tagcheck_way_s2 == 2'd0) ? mesi_state_way0_s2 :
                                (tagcheck_way_s2 == 2'd1) ? mesi_state_way1_s2 :
                                (tagcheck_way_s2 == 2'd2) ? mesi_state_way2_s2 :
                                                                     mesi_state_way3_s2 ;
    flush_way_s2 = address_s2[25:24];
    flush_state_s2 =  (flush_way_s2 == 2'd0) ? mesi_state_way0_s2 :
                            (flush_way_s2 == 2'd1) ? mesi_state_way1_s2 :
                            (flush_way_s2 == 2'd2) ? mesi_state_way2_s2 :
                                                             mesi_state_way3_s2 ;
    flush_way_tag_s2[(40 - 4 - ((9-2)))-1:0] =
                        (flush_way_s2 == 0) ? dtag_tag_way0_s2[(40 - 4 - ((9-2)))-1:0] :
                        (flush_way_s2 == 1) ? dtag_tag_way1_s2[(40 - 4 - ((9-2)))-1:0] :
                        (flush_way_s2 == 2) ? dtag_tag_way2_s2[(40 - 4 - ((9-2)))-1:0] :
                                                        dtag_tag_way3_s2[(40 - 4 - ((9-2)))-1:0];
    flush_way_address_s2 = {flush_way_tag_s2, address_s2[(((9-2))+4-1):4], 4'b0};
    
    tagcheck_state_me_s2 = tagcheck_state_s2 == 2'd3 || tagcheck_state_s2 == 2'd2;
    tagcheck_state_mes_s2 = tagcheck_state_s2 == 2'd3 || tagcheck_state_s2 == 2'd2
                                                        || tagcheck_state_s2 == 2'd1;
    tagcheck_state_s_s2 = tagcheck_state_s2 == 2'd1;
    tagcheck_state_m_s2 = tagcheck_state_s2 == 2'd3;
    tagcheck_state_e_s2 = tagcheck_state_s2 == 2'd2;
    lru_state_m_s2 = lru_state_s2 == 2'd3;
    lru_state_mes_s2 = lru_state_s2 == 2'd3 || lru_state_s2 == 2'd2
                                                        || lru_state_s2 == 2'd1;
    flush_state_m_s2 = flush_state_s2 == 2'd3;
    flush_state_me_s2 = flush_state_s2 == 2'd3 || flush_state_s2 == 2'd2;
    flush_state_mes_s2 = flush_state_s2 == 2'd3 || flush_state_s2 == 2'd2
                                                        || flush_state_s2 == 2'd1;
end
reg [4-1:0] lru_used_bits_s2;
reg [2-1:0] lru_round_robin_turn_s2;
always @ *
begin
    lru_used_bits_s2[4-1:0] = lruarray_l15_dout_s2[4-1:0];
    lru_round_robin_turn_s2[2-1:0] = lruarray_l15_dout_s2[4+2-1 -: 2];
    lru_way_s2 = 0;
    if (&lru_used_bits_s2 == 1'b1)
    begin
        
        lru_way_s2[2-1:0] = lru_round_robin_turn_s2;
    end
    else
    begin
        case (lru_round_robin_turn_s2)
            2'd0:
            begin
                lru_way_s2[2-1:0] = (lru_used_bits_s2[2'd0] == 1'b0) ? 2'd0 :
                                            (lru_used_bits_s2[2'd1] == 1'b0) ? 2'd1 :
                                            (lru_used_bits_s2[2'd2] == 1'b0) ? 2'd2 :
                                                                      2'd3 ;
            end
            2'd1:
            begin
                lru_way_s2[2-1:0] = (lru_used_bits_s2[2'd1] == 1'b0) ? 2'd1 :
                                            (lru_used_bits_s2[2'd2] == 1'b0) ? 2'd2 :
                                            (lru_used_bits_s2[2'd3] == 1'b0) ? 2'd3 :
                                                                      2'd0 ;
            end
            2'd2:
            begin
                lru_way_s2[2-1:0] = (lru_used_bits_s2[2'd2] == 1'b0) ? 2'd2 :
                                            (lru_used_bits_s2[2'd3] == 1'b0) ? 2'd3 :
                                            (lru_used_bits_s2[2'd0] == 1'b0) ? 2'd0 :
                                                                      2'd1 ;
            end
            2'd3:
            begin
                lru_way_s2[2-1:0] = (lru_used_bits_s2[2'd3] == 1'b0) ? 2'd3 :
                                            (lru_used_bits_s2[2'd0] == 1'b0) ? 2'd0 :
                                            (lru_used_bits_s2[2'd1] == 1'b0) ? 2'd1 :
                                                                      2'd2 ;
            end
        endcase
    end
end
reg s2_mshr_val_s2;
reg [2-1:0] s2_mshr_mshrid_s2;
always @ *
begin
    s2_mshr_val_s2 = 0;
    s2_mshr_mshrid_s2 = 0;
    case (s2_mshr_operation_s2)
        1'd1:
        begin
            s2_mshr_val_s2 = 1;
            s2_mshr_mshrid_s2 = mshrid_s2;
        end
    endcase
    
    
    pipe_mshr_write_buffer_rd_en_s2 = s2_mshr_val_s2;
    pipe_mshr_threadid_s2 = threadid_s2;
end
reg dcache_val_s2;
reg dcache_rw_s2;
reg [((9-2))-1:0] dcache_index_s2;
reg [1:0] dcache_way_s2;
reg [127:0] dcache_mshr_write_mask_s2;
reg [127:0] dcache_write_merge_mshr_noc2_s2;
reg [3-1:0] dcache_source_s2;
reg [127:0] dcache_write_mask_s2;
reg [127:0] dcache_write_data_s2;
reg [((9-2))-1:0] dcache_diag_index_s2;
reg [1:0] dcache_diag_way_s2;
reg [0:0] dcache_diag_offset_s2;
reg [1:0] lru_way_s3_bypassed;
always @ *
begin
    dcache_val_s2 = 0;
    dcache_rw_s2 = 0;
    dcache_index_s2 = 0;
    dcache_way_s2 = 0;
    dcache_mshr_write_mask_s2 = 0;
    dcache_write_merge_mshr_noc2_s2 = 0;
    dcache_source_s2 = 0;
    dcache_write_mask_s2 = 0;
    dcache_write_data_s2 = 0;
    dcache_diag_way_s2 = address_s2[25:24];
    dcache_diag_index_s2 = address_s2[(((9-2))+4-1):4];
    dcache_diag_offset_s2 = address_s2[3];
    case (dcache_operation_s2)
        4'd1:
        begin
            dcache_val_s2 = tagcheck_state_m_s2;
            dcache_rw_s2 = 1'b1;
            dcache_index_s2 = cache_index_s2;
            dcache_way_s2 = tagcheck_way_s2;
        end
        4'd2:
        begin
            dcache_val_s2 = tagcheck_state_mes_s2;
            dcache_rw_s2 = 1'b1;
            dcache_index_s2 = cache_index_s2;
            dcache_way_s2 = tagcheck_way_s2;
        end
        4'd3:
        begin
            dcache_val_s2 = lru_state_m_s2;
            dcache_rw_s2 = 1'b1;
            dcache_index_s2 = cache_index_s2;
            dcache_way_s2 = lru_way_s2;
        end
        4'd10:
        begin
            dcache_val_s2 = flush_state_m_s2;
            dcache_rw_s2 = 1'b1;
            dcache_index_s2 = cache_index_s2;
            dcache_way_s2 = flush_way_s2;
        end
        4'd4:
        begin
            dcache_val_s2 = tagcheck_state_me_s2;
            dcache_rw_s2 = 1'b0;
            dcache_index_s2 = cache_index_s2;
            dcache_way_s2 = tagcheck_way_s2;
            dcache_source_s2 = 3'd1;
        end
        4'd11:
        begin
            dcache_val_s2 = (tagcheck_state_m_s2 & tagcheck_lrsc_flag_s2); 
            dcache_rw_s2 = 1'b0;
            dcache_index_s2 = cache_index_s2;
            dcache_way_s2 = tagcheck_way_s2;
            dcache_source_s2 = 3'd1;
        end
        4'd5:
        begin
            dcache_val_s2 = 1'b1;
            dcache_rw_s2 = 1'b0;
            dcache_index_s2 = cache_index_s2;
            dcache_way_s2 = lru_way_s3_bypassed; 
            dcache_source_s2 = 3'd2;
        end
        4'd6:
        begin
            dcache_val_s2 = 1'b1;
            dcache_rw_s2 = 1'b0;
            dcache_index_s2 = cache_index_s2;
            dcache_way_s2 = lru_way_s3_bypassed; 
            dcache_source_s2 = 3'd3;
        end
        4'd7:
        begin
            
            dcache_val_s2 = 1'b1;
            dcache_rw_s2 = 1'b0;
            dcache_index_s2 = cache_index_s2;
            dcache_way_s2 = way_mshr_st_s2;
            dcache_source_s2 = 3'd1;
        end
        4'd8:
        begin
            dcache_val_s2 = 1'b1;
            dcache_rw_s2 = 1'b1;
            dcache_index_s2 = dcache_diag_index_s2;
            dcache_way_s2 = dcache_diag_way_s2;
        end
        4'd9:
        begin
            dcache_val_s2 = 1'b1;
            dcache_rw_s2 = 1'b0;
            dcache_index_s2 = dcache_diag_index_s2;
            dcache_way_s2 = dcache_diag_way_s2;
            dcache_source_s2 = 3'd4;
        end
    endcase
    dcache_mshr_write_mask_s2 = {
        {8{mshr_pipe_write_buffer_byte_mask_s2[15]}},
        {8{mshr_pipe_write_buffer_byte_mask_s2[14]}},
        {8{mshr_pipe_write_buffer_byte_mask_s2[13]}},
        {8{mshr_pipe_write_buffer_byte_mask_s2[12]}},
        {8{mshr_pipe_write_buffer_byte_mask_s2[11]}},
        {8{mshr_pipe_write_buffer_byte_mask_s2[10]}},
        {8{mshr_pipe_write_buffer_byte_mask_s2[9]}},
        {8{mshr_pipe_write_buffer_byte_mask_s2[8]}},
        {8{mshr_pipe_write_buffer_byte_mask_s2[7]}},
        {8{mshr_pipe_write_buffer_byte_mask_s2[6]}},
        {8{mshr_pipe_write_buffer_byte_mask_s2[5]}},
        {8{mshr_pipe_write_buffer_byte_mask_s2[4]}},
        {8{mshr_pipe_write_buffer_byte_mask_s2[3]}},
        {8{mshr_pipe_write_buffer_byte_mask_s2[2]}},
        {8{mshr_pipe_write_buffer_byte_mask_s2[1]}},
        {8{mshr_pipe_write_buffer_byte_mask_s2[0]}}
    };
    dcache_write_merge_mshr_noc2_s2[127:0] =
                    {(~dcache_mshr_write_mask_s2[127:64] & noc2decoder_l15_data_0[63:0]),
                    (~dcache_mshr_write_mask_s2[63:0] & noc2decoder_l15_data_1[63:0])}
                        | (dcache_mshr_write_mask_s2[127:0] & mshr_pipe_write_buffer_s2[127:0]);
    case (dcache_source_s2)
        3'd1:
        begin
            dcache_write_mask_s2[127:0] = dcache_mshr_write_mask_s2[127:0];
            dcache_write_data_s2[127:0] = mshr_pipe_write_buffer_s2[127:0];
        end
        3'd2:
        begin
            dcache_write_mask_s2[127:0] = {128{1'b1}};
            dcache_write_data_s2[127:0] = {noc2decoder_l15_data_0[63:0], noc2decoder_l15_data_1[63:0]};
        end
        3'd3:
        begin
            dcache_write_mask_s2[127:0] = {128{1'b1}};
            dcache_write_data_s2[127:0] = dcache_write_merge_mshr_noc2_s2[127:0];
        end
        3'd4:
        begin
            dcache_write_mask_s2[127:0] = dcache_diag_offset_s2 == 1'b0 ? {{64{1'b1}},64'b0} : {64'b0,{64{1'b1}}};
            dcache_write_data_s2[127:0] = {pcxdecoder_l15_data[63:0],pcxdecoder_l15_data[63:0]};
        end
    endcase
    l15_dcache_val_s2 = dcache_val_s2 && val_s2 && !stall_s2;
    l15_dcache_rw_s2 = dcache_rw_s2;
    l15_dcache_index_s2 = {dcache_index_s2, dcache_way_s2};
    l15_dcache_write_mask_s2[127:0] = dcache_write_mask_s2;
    l15_dcache_write_data_s2[127:0] = dcache_write_data_s2;
    
    
    
    
    
    l15_hmt_write_data_s2[14 + 8 + 8-1:0] = 0;
    l15_hmt_write_data_s2[14 + 8 + 8 - 1 -:  14] = hmt_fill_homeid_s2[((14+8+8)-1):(8+8)];
    l15_hmt_write_data_s2[8 + 8 - 1 -: 8] = hmt_fill_homeid_s2[8-1:0];
    l15_hmt_write_data_s2[8 - 1 -: 8] = hmt_fill_homeid_s2[8+8-1:8];
    
    
    
    l15_hmt_write_mask_s2 = 0;
    if (hmt_op_s2 == 1'd1)
      l15_hmt_write_mask_s2[14 + 8 + 8-1:0] = {14 + 8 + 8{1'b1}};
    
end
reg mesi_write_val_s2;
reg [((9-2))-1:0] mesi_write_index_s2;
reg [1:0] mesi_write_way_s2;
reg [1:0] mesi_write_state_s2;
always @ *
begin
    mesi_write_val_s2 = 0;
    mesi_write_index_s2 = 0;
    mesi_write_way_s2 = 0;
    mesi_write_state_s2 = 0;
    case (mesi_write_op_s2)
        3'd3:
        begin
            mesi_write_val_s2 = tagcheck_state_mes_s2;
            mesi_write_index_s2 = cache_index_s2;
            mesi_write_way_s2 = tagcheck_way_s2;
            mesi_write_state_s2 = 2'd0;
        end
        3'd6:
        begin
            mesi_write_val_s2 = flush_state_mes_s2;
            mesi_write_index_s2 = cache_index_s2;
            mesi_write_way_s2 = flush_way_s2;
            mesi_write_state_s2 = 2'd0;
        end
        3'd1:
        begin
            mesi_write_val_s2 = tagcheck_state_me_s2;
            mesi_write_index_s2 = cache_index_s2;
            mesi_write_way_s2 = tagcheck_way_s2;
            mesi_write_state_s2 = 2'd1;
        end
        3'd2:
        begin
            mesi_write_val_s2 = tagcheck_state_e_s2;
            mesi_write_index_s2 = cache_index_s2;
            mesi_write_way_s2 = tagcheck_way_s2;
            mesi_write_state_s2 = 2'd3;
        end
        3'd4:
        begin
            mesi_write_val_s2 = 1'b1;
            mesi_write_index_s2 = cache_index_s2;
            mesi_write_way_s2 = lru_way_s2;
            mesi_write_state_s2 = noc2_ack_state_s2;
        end
        3'd5:
        begin
            mesi_write_val_s2 = 1'b1;
            mesi_write_index_s2 = cache_index_s2;
            mesi_write_way_s2 = way_mshr_st_s2;
            mesi_write_state_s2 = noc2_ack_state_s2;
        end
    endcase
    
    
    l15_mesi_write_val_s2 = mesi_write_val_s2 && val_s2 && !stall_s2;
    l15_mesi_write_index_s2[((9-2))-1:0] = mesi_write_index_s2;
    l15_mesi_write_mask_s2[7:0] =  (mesi_write_way_s2 == 0) ? 8'b00_00_00_11 :
                            (mesi_write_way_s2 == 1) ? 8'b00_00_11_00 :
                            (mesi_write_way_s2 == 2) ? 8'b00_11_00_00 :
                                                    8'b11_00_00_00 ;
    l15_mesi_write_data_s2[7:0] = {4{mesi_write_state_s2}};
end
reg lrsc_flag_write_val_s2;
reg [((9-2))-1:0] lrsc_flag_write_index_s2;
reg [1:0] lrsc_flag_write_way_s2;
reg lrsc_flag_write_state_s2;
always @ *
begin
    lrsc_flag_write_val_s2 = 0;
    lrsc_flag_write_index_s2 = 0;
    lrsc_flag_write_way_s2 = 0;
    lrsc_flag_write_state_s2 = 0;
    case (lrsc_flag_write_op_s2)
        3'd1:
        begin
            lrsc_flag_write_val_s2 = 1'b1;
            lrsc_flag_write_index_s2 = cache_index_s2;
            lrsc_flag_write_way_s2 = lru_way_s2;
            lrsc_flag_write_state_s2 = 1'b1;
        end
        3'd2:  
        begin
            lrsc_flag_write_val_s2 = tagcheck_state_m_s2;  
            lrsc_flag_write_index_s2 = cache_index_s2;
            lrsc_flag_write_way_s2 = tagcheck_way_s2;
            lrsc_flag_write_state_s2 = 1'b0;
        end
        3'd3:  
        begin
            lrsc_flag_write_val_s2 = 1'b1;
            lrsc_flag_write_index_s2 = cache_index_s2;
            lrsc_flag_write_way_s2 = lru_way_s2;
            lrsc_flag_write_state_s2 = 1'b0;
        end
        3'd4:  
        begin
            lrsc_flag_write_val_s2 = flush_state_m_s2;
            lrsc_flag_write_index_s2 = cache_index_s2;
            lrsc_flag_write_way_s2 = flush_way_s2;
            lrsc_flag_write_state_s2 = 1'b0;
        end
    endcase
    
    
    l15_lrsc_flag_write_val_s2 = lrsc_flag_write_val_s2 && val_s2 && !stall_s2;
    l15_lrsc_flag_write_index_s2[((9-2))-1:0] = lrsc_flag_write_index_s2;
    l15_lrsc_flag_write_mask_s2[3:0] =  (lrsc_flag_write_way_s2 == 0) ? 4'b0001 :
                            (lrsc_flag_write_way_s2 == 1) ? 4'b0010 :
                            (lrsc_flag_write_way_s2 == 2) ? 4'b0100 :
                                                    4'b1000 ;
    l15_lrsc_flag_write_data_s2[3:0] = {4{lrsc_flag_write_state_s2}};
end
reg [3-1:0] csm_ticket_s2;
reg [127:0] csm_fill_data;
reg csm_req_val_s2;
reg csm_req_type_s2;
reg csm_req_lru_address_s2;
reg [39:0] csm_address_s2;
always @ *
begin
    
    
    csm_fill_data = 0;
    csm_req_val_s2 = 0;
    csm_req_type_s2 = 0;
    csm_req_lru_address_s2 = 0;
    csm_address_s2 = 0;
    
    csm_ticket_s2 = {threadid_s2, mshrid_s2};
    l15_csm_req_ticket_s2 = csm_ticket_s2;
    case (csm_op_s2)
        4'd1:
        begin
            csm_req_val_s2 = 1'b1;
            csm_req_type_s2 = 1'b0;
            
            csm_address_s2 = address_s2;
            
        end
        4'd2:
        begin
            csm_req_val_s2 = (tagcheck_state_me_s2 == 1'b0);
            csm_req_type_s2 = 1'b0;
            
            csm_address_s2 = address_s2;
            
        end
        4'd6:
        begin
            csm_req_val_s2 = (tagcheck_state_mes_s2 == 1'b0);
            csm_req_type_s2 = 1'b0;
            
            csm_address_s2 = address_s2;
            
        end
        4'd3:
        begin
            csm_req_val_s2 = 1'b1;
            csm_req_type_s2 = 1'b1;
            csm_fill_data = {noc2decoder_l15_data_1[63:0], noc2decoder_l15_data_0[63:0]};
            
            l15_csm_req_ticket_s2 = noc2decoder_l15_csm_mshrid[3-1:0];
        end
        4'd4:
        begin
            csm_req_val_s2 = 1'b1;
            csm_req_type_s2 = 1'b1;
            csm_fill_data = {pcxdecoder_l15_data[63:0],pcxdecoder_l15_data[63:0]};
            
            csm_address_s2 = address_s2;
        end
        4'd5:
        begin
            csm_req_val_s2 = 1'b1;
            csm_req_type_s2 = 1'b0;
            
            csm_address_s2 = address_s2;
        end
        4'd7:
        begin
            csm_req_val_s2 = 1'b1;
            
            
            csm_address_s2 = address_s2;
        end
        
        
        
    endcase
    l15_csm_req_address_s2 = csm_address_s2;
    l15_csm_req_val_s2 = csm_req_val_s2 && !stall_s2 && val_s2;
    l15_csm_req_type_s2 = csm_req_type_s2;
    
    
    l15_csm_req_data_s2 = csm_fill_data[127:0];
    l15_csm_req_pcx_data_s2 = csm_pcx_data_s2;
end
reg wmt_read_val_s2;
reg [6:0] wmt_read_index_s2;
always @ *
begin
    wmt_read_val_s2 = 0;
    wmt_read_index_s2 = 0;
    case(wmt_read_op_s2)
        1'd1:
        begin
            wmt_read_val_s2 = 1'b1;
            wmt_read_index_s2 = cache_index_l1d_s2[6:0];
            
        end
    endcase
    l15_wmt_read_val_s2 = wmt_read_val_s2 && val_s2 && !stall_s2;
    l15_wmt_read_index_s2 = wmt_read_index_s2;
end
reg config_req_val_s2;
reg config_req_rw_s2;
reg [63:0] config_write_req_data_s2;
reg [39:0] config_req_address_s2;
always @ *
begin
    config_req_val_s2 = 0;
    config_req_rw_s2 = 0;
    config_write_req_data_s2 = 0;
    config_req_address_s2 = 0;
    case (config_op_s2)
        2'd1:
        begin
            config_req_val_s2 = 1'b1;
            config_req_rw_s2 = 1'b0;
            config_req_address_s2 = address_s2;
        end
        2'd2:
        begin
            config_req_val_s2 = 1'b1;
            config_req_rw_s2 = 1'b1;
            config_req_address_s2 = address_s2;
            config_write_req_data_s2[63:0] = pcxdecoder_l15_data[63:0];
        end
    endcase
    l15_config_req_val_s2 = config_req_val_s2 && val_s2 && !stall_s2;
    l15_config_req_rw_s2 = config_req_rw_s2;
    l15_config_write_req_data_s2 = config_write_req_data_s2;
    l15_config_req_address_s2 = config_req_address_s2[15:8];
end
reg [2-1:0] tagcheck_way_s3;
reg [2-1:0] tagcheck_way_s3_next;
reg [2-1:0] tagcheck_state_s3;
reg [2-1:0] tagcheck_state_s3_next;
reg [1-1:0] tagcheck_lrsc_flag_s3;
reg [1-1:0] tagcheck_lrsc_flag_s3_next;
reg [2-1:0] flush_way_s3;
reg [2-1:0] flush_way_s3_next;
reg [2-1:0] flush_state_s3;
reg [2-1:0] flush_state_s3_next;
reg [2-1:0] lru_way_s3;
reg [2-1:0] lru_way_s3_next;
reg [2-1:0] lru_state_s3;
reg [2-1:0] lru_state_s3_next;
reg [2-1:0] mshrid_s3;
reg [2-1:0] mshrid_s3_next;
reg [40-1:0] address_s3;
reg [40-1:0] address_s3_next;
reg [1-1:0] threadid_s3;
reg [1-1:0] threadid_s3_next;
reg [1-1:0] non_cacheable_s3;
reg [1-1:0] non_cacheable_s3_next;
reg [3-1:0] size_s3;
reg [3-1:0] size_s3_next;
reg [1-1:0] prefetch_s3;
reg [1-1:0] prefetch_s3_next;
reg [2-1:0] l1_replacement_way_s3;
reg [2-1:0] l1_replacement_way_s3_next;
reg [1-1:0] l2_miss_s3;
reg [1-1:0] l2_miss_s3_next;
reg [1-1:0] f4b_s3;
reg [1-1:0] f4b_s3_next;
reg [1-1:0] blockstore_s3;
reg [1-1:0] blockstore_s3_next;
reg [1-1:0] blockstoreinit_s3;
reg [1-1:0] blockstoreinit_s3_next;
reg [(14+8+8)-1:0] noc2_src_homeid_s3;
reg [(14+8+8)-1:0] noc2_src_homeid_s3_next;
reg [3-1:0] lruarray_write_op_s3;
reg [3-1:0] lruarray_write_op_s3_next;
reg [1-1:0] predecode_noc2_inval_s3;
reg [1-1:0] predecode_noc2_inval_s3_next;
reg [4-1:0] predecode_fwd_subcacheline_vector_s3;
reg [4-1:0] predecode_fwd_subcacheline_vector_s3_next;
reg [6-1:0] predecode_reqtype_s3;
reg [6-1:0] predecode_reqtype_s3_next;
reg [3-1:0] wmt_write_op_s3;
reg [3-1:0] wmt_write_op_s3_next;
reg [3-1:0] wmt_compare_op_s3;
reg [3-1:0] wmt_compare_op_s3_next;
reg [3-1:0] csm_ticket_s3;
reg [3-1:0] csm_ticket_s3_next;
reg [3-1:0] s3_mshr_operation_s3;
reg [3-1:0] s3_mshr_operation_s3_next;
reg [5-1:0] cpx_operation_s3;
reg [5-1:0] cpx_operation_s3_next;
reg [5-1:0] noc1_operation_s3;
reg [5-1:0] noc1_operation_s3_next;
reg [4-1:0] noc3_operations_s3;
reg [4-1:0] noc3_operations_s3_next;
reg [2-1:0] pcx_ack_stage_s3;
reg [2-1:0] pcx_ack_stage_s3_next;
reg [2-1:0] noc2_ack_stage_s3;
reg [2-1:0] noc2_ack_stage_s3_next;
reg [2-1:0] noc2_ack_state_s3;
reg [2-1:0] noc2_ack_state_s3_next;
reg [(40 - 4 - ((9-2)))-1:0] lru_way_tag_s3;
reg [(40 - 4 - ((9-2)))-1:0] lru_way_tag_s3_next;
reg [(40 - 4 - ((9-2)))-1:0] flush_way_tag_s3;
reg [(40 - 4 - ((9-2)))-1:0] flush_way_tag_s3_next;
reg [33-1:0] csm_pcx_data_s3;
reg [33-1:0] csm_pcx_data_s3_next;
reg val_s3_next;
reg [(2 + 4)-1:0] lru_data_s3;
reg cpxencoder_req_staled_s3;
reg cpxencoder_req_staled_s3_next;
reg noc1encoder_req_staled_s3;
reg noc1encoder_req_staled_s3_next;
reg noc3encoder_req_staled_s3;
reg noc3encoder_req_staled_s3_next;
reg stall_for_cpx_s3;
reg stall_for_noc3_s3;
reg tagcheck_state_me_s3;
reg tagcheck_state_mes_s3;
reg tagcheck_state_s_s3;
reg tagcheck_state_e_s3;
reg tagcheck_state_m_s3;
reg lru_state_m_s3;
reg lru_state_mes_s3;
reg flush_state_m_s3;
reg flush_state_mes_s3;
reg [39:0] lru_way_address_s3;
reg [39:0] flush_way_address_s3;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        cpxencoder_req_staled_s3 <= 0;
        noc1encoder_req_staled_s3 <= 0;
        noc3encoder_req_staled_s3 <= 0;
        val_s3 <= 0;
        lru_data_s3 <= 0;
        tagcheck_way_s3 <= 0;
tagcheck_state_s3 <= 0;
tagcheck_lrsc_flag_s3 <= 0;
flush_way_s3 <= 0;
flush_state_s3 <= 0;
lru_way_s3 <= 0;
lru_state_s3 <= 0;
mshrid_s3 <= 0;
address_s3 <= 0;
threadid_s3 <= 0;
non_cacheable_s3 <= 0;
size_s3 <= 0;
prefetch_s3 <= 0;
l1_replacement_way_s3 <= 0;
l2_miss_s3 <= 0;
f4b_s3 <= 0;
blockstore_s3 <= 0;
blockstoreinit_s3 <= 0;
noc2_src_homeid_s3 <= 0;
lruarray_write_op_s3 <= 0;
predecode_noc2_inval_s3 <= 0;
predecode_fwd_subcacheline_vector_s3 <= 0;
predecode_reqtype_s3 <= 0;
wmt_write_op_s3 <= 0;
wmt_compare_op_s3 <= 0;
csm_ticket_s3 <= 0;
s3_mshr_operation_s3 <= 0;
cpx_operation_s3 <= 0;
noc1_operation_s3 <= 0;
noc3_operations_s3 <= 0;
pcx_ack_stage_s3 <= 0;
noc2_ack_stage_s3 <= 0;
noc2_ack_state_s3 <= 0;
lru_way_tag_s3 <= 0;
flush_way_tag_s3 <= 0;
csm_pcx_data_s3 <= 0;
    end
    else
    begin
        cpxencoder_req_staled_s3 <= cpxencoder_req_staled_s3_next;
        noc1encoder_req_staled_s3 <= noc1encoder_req_staled_s3_next;
        noc3encoder_req_staled_s3 <= noc3encoder_req_staled_s3_next;
        val_s3 <= val_s3_next;
        lru_data_s3 <= lruarray_l15_dout_s2;
        tagcheck_way_s3 <= tagcheck_way_s3_next;
tagcheck_state_s3 <= tagcheck_state_s3_next;
tagcheck_lrsc_flag_s3 <= tagcheck_lrsc_flag_s3_next;
flush_way_s3 <= flush_way_s3_next;
flush_state_s3 <= flush_state_s3_next;
lru_way_s3 <= lru_way_s3_next;
lru_state_s3 <= lru_state_s3_next;
mshrid_s3 <= mshrid_s3_next;
address_s3 <= address_s3_next;
threadid_s3 <= threadid_s3_next;
non_cacheable_s3 <= non_cacheable_s3_next;
size_s3 <= size_s3_next;
prefetch_s3 <= prefetch_s3_next;
l1_replacement_way_s3 <= l1_replacement_way_s3_next;
l2_miss_s3 <= l2_miss_s3_next;
f4b_s3 <= f4b_s3_next;
blockstore_s3 <= blockstore_s3_next;
blockstoreinit_s3 <= blockstoreinit_s3_next;
noc2_src_homeid_s3 <= noc2_src_homeid_s3_next;
lruarray_write_op_s3 <= lruarray_write_op_s3_next;
predecode_noc2_inval_s3 <= predecode_noc2_inval_s3_next;
predecode_fwd_subcacheline_vector_s3 <= predecode_fwd_subcacheline_vector_s3_next;
predecode_reqtype_s3 <= predecode_reqtype_s3_next;
wmt_write_op_s3 <= wmt_write_op_s3_next;
wmt_compare_op_s3 <= wmt_compare_op_s3_next;
csm_ticket_s3 <= csm_ticket_s3_next;
s3_mshr_operation_s3 <= s3_mshr_operation_s3_next;
cpx_operation_s3 <= cpx_operation_s3_next;
noc1_operation_s3 <= noc1_operation_s3_next;
noc3_operations_s3 <= noc3_operations_s3_next;
pcx_ack_stage_s3 <= pcx_ack_stage_s3_next;
noc2_ack_stage_s3 <= noc2_ack_stage_s3_next;
noc2_ack_state_s3 <= noc2_ack_state_s3_next;
lru_way_tag_s3 <= lru_way_tag_s3_next;
flush_way_tag_s3 <= flush_way_tag_s3_next;
csm_pcx_data_s3 <= csm_pcx_data_s3_next;
    end
end
reg [1:0] stbuf_compare_address_match_s3;
reg [1:0] stbuf_compare_match_s3;
reg [1:0] stbuf_compare_lru_match_s3;
reg [0:0] stbuf_compare_threadid_s3;
reg [0:0] stbuf_compare_lru_threadid_s3;
reg stbuf_compare_match_val_s3;
reg stbuf_compare_lru_match_val_s3;
reg [1:0] stbuf_way_s3; 
always @ *
begin
    stbuf_compare_address_match_s3[0] = mshr_st_address_array[0][39:4] == address_s3[39:4];
    stbuf_compare_match_s3[0] = mshr_val_array[0][2'd3] 
                                && (mshr_st_state_array[0] == 2'b01) 
                                && (stbuf_compare_address_match_s3[0] == 1'b1);
    stbuf_compare_lru_match_s3[0] = stbuf_compare_match_s3[0] && (mshr_st_way_array[0] == lru_way_s3);
    stbuf_compare_address_match_s3[1] = mshr_st_address_array[1][39:4] == address_s3[39:4];
    stbuf_compare_match_s3[1] = mshr_val_array[1][2'd3] 
                                && (mshr_st_state_array[1] == 2'b01) 
                                && (stbuf_compare_address_match_s3[1] == 1'b1);
    stbuf_compare_lru_match_s3[1] = stbuf_compare_match_s3[1] && (mshr_st_way_array[1] == lru_way_s3);
    stbuf_compare_threadid_s3 = stbuf_compare_match_s3[1] ? 1'b1 : 1'b0;
    stbuf_compare_lru_threadid_s3 = stbuf_compare_lru_match_s3[1] ? 1'b1 : 1'b0;
    stbuf_compare_match_val_s3 = stbuf_compare_match_s3[0] || stbuf_compare_match_s3[1];
    stbuf_compare_lru_match_val_s3 = stbuf_compare_lru_match_s3[0] || stbuf_compare_lru_match_s3[1];
    stbuf_way_s3 = mshr_st_way_array[stbuf_compare_threadid_s3];
    
    
    
end
reg [3:0] tagcheck_way_mask_s3;
always @ *
begin
    
    tagcheck_way_mask_s3[3:0] = tagcheck_way_s3 == 2'd0 ? 4'b0001 :
                                                  2'd1 ? 4'b0010 :
                                                  2'd2 ? 4'b0100 :
                                                        4'b1000 ;
    tagcheck_state_me_s3 = tagcheck_state_s3 == 2'd3 || tagcheck_state_s3 == 2'd2;
    tagcheck_state_mes_s3 = tagcheck_state_s3 == 2'd3 || tagcheck_state_s3 == 2'd2
                                                        || tagcheck_state_s3 == 2'd1;
    tagcheck_state_s_s3 = tagcheck_state_s3 == 2'd1;
    tagcheck_state_m_s3 = tagcheck_state_s3 == 2'd3;
    tagcheck_state_e_s3 = tagcheck_state_s3 == 2'd2;
    lru_state_m_s3 = lru_state_s3 == 2'd3;
    lru_state_mes_s3 = lru_state_s3 == 2'd3 || lru_state_s3 == 2'd2
                                                        || lru_state_s3 == 2'd1;
    flush_state_m_s3 = flush_state_s3 == 2'd3;
    flush_state_mes_s3 = flush_state_s3 == 2'd3 || flush_state_s3 == 2'd2
                                                        || flush_state_s3 == 2'd1;
    cache_index_s3 = address_s3[(((9-2))+4-1):4];
    cache_index_l1d_s3 = address_s3[(6 + 4):4];
    lru_way_address_s3 = {lru_way_tag_s3, cache_index_s3, 4'b0};
    flush_way_address_s3 = {flush_way_tag_s3, cache_index_s3, 4'b0};
end
always @* begin
    
    if (stall_s3)
    begin
        val_s3_next = val_s3;
        tagcheck_way_s3_next = tagcheck_way_s3;
tagcheck_state_s3_next = tagcheck_state_s3;
tagcheck_lrsc_flag_s3_next = tagcheck_lrsc_flag_s3;
flush_way_s3_next = flush_way_s3;
flush_state_s3_next = flush_state_s3;
lru_way_s3_next = lru_way_s3;
lru_state_s3_next = lru_state_s3;
mshrid_s3_next = mshrid_s3;
address_s3_next = address_s3;
threadid_s3_next = threadid_s3;
non_cacheable_s3_next = non_cacheable_s3;
size_s3_next = size_s3;
prefetch_s3_next = prefetch_s3;
l1_replacement_way_s3_next = l1_replacement_way_s3;
l2_miss_s3_next = l2_miss_s3;
f4b_s3_next = f4b_s3;
blockstore_s3_next = blockstore_s3;
blockstoreinit_s3_next = blockstoreinit_s3;
noc2_src_homeid_s3_next = noc2_src_homeid_s3;
lruarray_write_op_s3_next = lruarray_write_op_s3;
predecode_noc2_inval_s3_next = predecode_noc2_inval_s3;
predecode_fwd_subcacheline_vector_s3_next = predecode_fwd_subcacheline_vector_s3;
predecode_reqtype_s3_next = predecode_reqtype_s3;
wmt_write_op_s3_next = wmt_write_op_s3;
wmt_compare_op_s3_next = wmt_compare_op_s3;
csm_ticket_s3_next = csm_ticket_s3;
s3_mshr_operation_s3_next = s3_mshr_operation_s3;
cpx_operation_s3_next = cpx_operation_s3;
noc1_operation_s3_next = noc1_operation_s3;
noc3_operations_s3_next = noc3_operations_s3;
pcx_ack_stage_s3_next = pcx_ack_stage_s3;
noc2_ack_stage_s3_next = noc2_ack_stage_s3;
noc2_ack_state_s3_next = noc2_ack_state_s3;
lru_way_tag_s3_next = lru_way_tag_s3;
flush_way_tag_s3_next = flush_way_tag_s3;
csm_pcx_data_s3_next = csm_pcx_data_s3;
    end
    else
    begin
        val_s3_next = val_s2 && !stall_s2;
        tagcheck_way_s3_next = tagcheck_way_s2;
tagcheck_state_s3_next = tagcheck_state_s2;
tagcheck_lrsc_flag_s3_next = tagcheck_lrsc_flag_s2;
flush_way_s3_next = flush_way_s2;
flush_state_s3_next = flush_state_s2;
lru_way_s3_next = lru_way_s2;
lru_state_s3_next = lru_state_s2;
mshrid_s3_next = mshrid_s2;
address_s3_next = address_s2;
threadid_s3_next = threadid_s2;
non_cacheable_s3_next = non_cacheable_s2;
size_s3_next = size_s2;
prefetch_s3_next = prefetch_s2;
l1_replacement_way_s3_next = l1_replacement_way_s2;
l2_miss_s3_next = l2_miss_s2;
f4b_s3_next = f4b_s2;
blockstore_s3_next = blockstore_s2;
blockstoreinit_s3_next = blockstoreinit_s2;
noc2_src_homeid_s3_next = noc2_src_homeid_s2;
lruarray_write_op_s3_next = lruarray_write_op_s2;
predecode_noc2_inval_s3_next = predecode_noc2_inval_s2;
predecode_fwd_subcacheline_vector_s3_next = predecode_fwd_subcacheline_vector_s2;
predecode_reqtype_s3_next = predecode_reqtype_s2;
wmt_write_op_s3_next = wmt_write_op_s2;
wmt_compare_op_s3_next = wmt_compare_op_s2;
csm_ticket_s3_next = csm_ticket_s2;
s3_mshr_operation_s3_next = s3_mshr_operation_s2;
cpx_operation_s3_next = cpx_operation_s2;
noc1_operation_s3_next = noc1_operation_s2;
noc3_operations_s3_next = noc3_operations_s2;
pcx_ack_stage_s3_next = pcx_ack_stage_s2;
noc2_ack_stage_s3_next = noc2_ack_stage_s2;
noc2_ack_state_s3_next = noc2_ack_state_s2;
lru_way_tag_s3_next = lru_way_tag_s2;
flush_way_tag_s3_next = flush_way_tag_s2;
csm_pcx_data_s3_next = csm_pcx_data_s2;
    end
end
always @* begin
    
    if (!cpxencoder_req_staled_s3)
        cpxencoder_req_staled_s3_next = (!stall_for_cpx_s3 && stall_for_noc3_s3) ? 1'b1 : 1'b0;
    else
        cpxencoder_req_staled_s3_next = stall_s3 ? 1'b1 : 1'b0;
end
always @* begin
    if (!noc1encoder_req_staled_s3)
        noc1encoder_req_staled_s3_next = (stall_for_cpx_s3 || stall_for_noc3_s3) ? 1'b1 : 1'b0;
    else
        noc1encoder_req_staled_s3_next = stall_s3 ? 1'b1 : 1'b0;
end
always @* begin
    if (!noc3encoder_req_staled_s3)
        noc3encoder_req_staled_s3_next = (!stall_for_noc3_s3 && stall_for_cpx_s3) ? 1'b1 : 1'b0;
    else
        noc3encoder_req_staled_s3_next = stall_s3 ? 1'b1 : 1'b0;
end
always @* begin
    
    
    
    
    
    stall_for_cpx_s3 = !cpxencoder_req_staled_s3 && l15_cpxencoder_val && !cpxencoder_l15_req_ack;
    
    stall_for_noc3_s3 = !noc3encoder_req_staled_s3 && l15_noc3encoder_req_val && !noc3encoder_l15_req_ack;
    stall_s3 = val_s3 && (stall_for_cpx_s3 || stall_for_noc3_s3);
    
    pcx_ack_s3 = val_s3 && !stall_s3 && (pcx_ack_stage_s3 == 2'd3);
    noc2_ack_s3 = val_s3 && !stall_s3 && (noc2_ack_stage_s3 == 2'd3);
    
    l15_csm_stall_s3 = stall_s3;
    
    lru_way_s3_bypassed = lru_way_s3;
end
reg [(2+0)-1:0] wmt_compare_data_s3;
reg [2-1:0] wmt_compare_way_s3;
reg [((2+0)+1)-1:0] wmt_data_s3 [0:4-1];
reg [4-1:0] wmt_compare_mask_s3;
reg wmt_compare_match_s3;
reg [2-1:0] wmt_compare_match_way_s3;
always @ *
begin
    
    
    
    
    
    
  wmt_data_s3[0] = wmt_l15_data_s3[(0+1)*((2+0)+1)-1 -: ((2+0)+1)];
  wmt_data_s3[1] = wmt_l15_data_s3[(1+1)*((2+0)+1)-1 -: ((2+0)+1)];
  wmt_data_s3[2] = wmt_l15_data_s3[(2+1)*((2+0)+1)-1 -: ((2+0)+1)];
  wmt_data_s3[3] = wmt_l15_data_s3[(3+1)*((2+0)+1)-1 -: ((2+0)+1)];
    wmt_compare_data_s3 = 0;
    wmt_compare_way_s3 = 0;
    case (wmt_compare_op_s3)
        3'd1:
        begin
            wmt_compare_way_s3 = lru_way_s3;
        end
        3'd2:
        begin
            wmt_compare_way_s3 = tagcheck_way_s3;
        end
        3'd3:
        begin
            wmt_compare_way_s3 = flush_way_s3;
        end
        3'd4:
        begin
            wmt_compare_way_s3 = stbuf_way_s3;
        end
    endcase
    wmt_compare_data_s3 = wmt_compare_way_s3;
    
    
    
    
    
    
    
    
  wmt_compare_mask_s3[0] = wmt_data_s3[0][(2+0)] && (wmt_compare_data_s3[(2+0)-1:0] == wmt_data_s3[0][(2+0)-1:0]);
  wmt_compare_mask_s3[1] = wmt_data_s3[1][(2+0)] && (wmt_compare_data_s3[(2+0)-1:0] == wmt_data_s3[1][(2+0)-1:0]);
  wmt_compare_mask_s3[2] = wmt_data_s3[2][(2+0)] && (wmt_compare_data_s3[(2+0)-1:0] == wmt_data_s3[2][(2+0)-1:0]);
  wmt_compare_mask_s3[3] = wmt_data_s3[3][(2+0)] && (wmt_compare_data_s3[(2+0)-1:0] == wmt_data_s3[3][(2+0)-1:0]);
    
    wmt_compare_match_s3 = |wmt_compare_mask_s3;
    
                               
                               
                                                        
    wmt_compare_match_way_s3 = 0;
if (wmt_compare_mask_s3[0])
   wmt_compare_match_way_s3 = 0;
else if (wmt_compare_mask_s3[1])
   wmt_compare_match_way_s3 = 1;
else if (wmt_compare_mask_s3[2])
   wmt_compare_match_way_s3 = 2;
else if (wmt_compare_mask_s3[3])
   wmt_compare_match_way_s3 = 3;
end
reg [(2 + 4)-1:0] lruarray_write_data_s3;
reg lruarray_write_val_s3;
reg [3:0] lruarray_lru_mask_s3;
reg [3:0] lruarray_tagcheck_mask_s3;
reg [3:0] lruarray_flush_mask_s3;
reg [((9-2))-1:0] lruarray_write_index_s3;
always @ *
begin
    lruarray_write_data_s3 = 0;
    lruarray_write_val_s3 = 0;
    lruarray_lru_mask_s3 = lru_way_s3[1:0] == 2'd0 ? 4'b0001 :
                                  lru_way_s3[1:0] == 2'd1 ? 4'b0010 :
                                  lru_way_s3[1:0] == 2'd2 ? 4'b0100 :
                                                                     4'b1000 ;
    lruarray_flush_mask_s3 =   flush_way_s3[1:0] == 2'd0 ? 4'b0001 :
                                        flush_way_s3[1:0] == 2'd1 ? 4'b0010 :
                                        flush_way_s3[1:0] == 2'd2 ? 4'b0100 :
                                                                            4'b1000 ;
    lruarray_tagcheck_mask_s3 = tagcheck_way_mask_s3;
    case (lruarray_write_op_s3)
        3'd1:
        begin
            lruarray_write_val_s3 = tagcheck_state_mes_s3;
            if ((lru_data_s3[3:0] | lruarray_tagcheck_mask_s3) == 4'b1111)
                lruarray_write_data_s3[3:0] = 4'b0000;
            else
                lruarray_write_data_s3[3:0] = lru_data_s3[3:0] | lruarray_tagcheck_mask_s3;
            lruarray_write_data_s3[5:4] = lru_data_s3[5:4]; 
        end
        3'd6:
        begin
            lruarray_write_val_s3 = tagcheck_lrsc_flag_s3;
            if ((lru_data_s3[3:0] | lruarray_tagcheck_mask_s3) == 4'b1111)
                lruarray_write_data_s3[3:0] = 4'b0000;
            else
                lruarray_write_data_s3[3:0] = lru_data_s3[3:0] | lruarray_tagcheck_mask_s3;
            lruarray_write_data_s3[5:4] = lru_data_s3[5:4]; 
        end
        3'd2:
        begin
            
            
            
            
        end
        3'd3:
        begin
            
            
            
            
            lruarray_write_val_s3 = 1'b1; 
            lruarray_write_data_s3[3:0] = lru_data_s3[3:0] | lruarray_lru_mask_s3;
            lruarray_write_data_s3[5:4] = lru_data_s3[5:4] + 2'b1;
        end
        3'd4:
        begin
            lruarray_write_val_s3 = tagcheck_state_mes_s3;
            lruarray_write_data_s3[3:0] = lru_data_s3[3:0] & ~lruarray_tagcheck_mask_s3;
                
            lruarray_write_data_s3[5:4] = lru_data_s3[5:4];
        end
        3'd5:
        begin
            lruarray_write_val_s3 = flush_state_mes_s3;
            lruarray_write_data_s3[3:0] = lru_data_s3[3:0] & ~lruarray_flush_mask_s3;
                
            lruarray_write_data_s3[5:4] = lru_data_s3[5:4];
        end
    endcase
    lruarray_write_index_s3 = cache_index_s3;
    l15_lruarray_write_val_s3 = lruarray_write_val_s3 && val_s3;
    l15_lruarray_write_data_s3 = lruarray_write_data_s3;
    l15_lruarray_write_mask_s3 = 6'b111111;
    
    l15_lruarray_write_index_s3 = lruarray_write_index_s3;
end
reg wmt_write_val_s3;
reg [6:0] wmt_write_index_s3;
reg [4*((2+0)+1)-1:0] wmt_write_data_s3;
reg wmt_write_inval_val_s3;
reg wmt_write_update_val_s3;
reg wmt_write_dedup_l1way_val_s3;
reg [2-1:0] wmt_write_update_way_s3;
reg [4*((2+0)+1)-1:0] wmt_write_inval_mask_s3;
reg [4*((2+0)+1)-1:0] wmt_write_update_mask_s3;
reg [4*((2+0)+1)-1:0] wmt_write_dedup_mask_s3;
reg [4*((2+0)+1)-1:0] wmt_write_mask_s3;
reg [(2+0)-1:0] wmt_write_update_data_s3;
reg [0-1:0] wmt_alias_bits;
always @ *
begin
    wmt_write_val_s3 = 0;
    wmt_write_index_s3 = 0;
    wmt_write_inval_val_s3 = 0;
    wmt_write_update_val_s3 = 0;
    wmt_write_dedup_l1way_val_s3 = 0;
    wmt_write_update_way_s3 = 0;
    wmt_write_update_data_s3 = 0;
    
    
    wmt_write_inval_mask_s3 = 0;
    wmt_write_update_mask_s3 = 0;
    wmt_write_dedup_mask_s3 = 0;
    case(wmt_write_op_s3)
        3'd1:
        begin
            wmt_write_val_s3 = tagcheck_state_mes_s3;
            wmt_write_index_s3 = cache_index_l1d_s3[6:0];
            wmt_write_inval_val_s3 = 1'b1;
            
        end
        3'd2:
        begin
            wmt_write_val_s3 = lru_state_mes_s3;
            wmt_write_index_s3 = cache_index_l1d_s3[6:0];
            wmt_write_inval_val_s3 = 1'b1;
            
        end
        3'd5:
        begin
            wmt_write_val_s3 = val_s3 && flush_state_mes_s3;
            wmt_write_index_s3 = cache_index_l1d_s3[6:0];
            wmt_write_inval_val_s3 = 1'b1;
            
        end
        3'd3: 
        begin
            wmt_write_val_s3 = 1'b1;
            wmt_write_index_s3 = cache_index_l1d_s3[6:0];
            wmt_write_update_val_s3 = 1'b1;
            wmt_write_update_way_s3 = lru_way_s3;
            wmt_write_inval_val_s3 = 1'b1;
        end
        3'd4:
        begin
            wmt_write_val_s3 = tagcheck_state_mes_s3;
            wmt_write_index_s3 = cache_index_l1d_s3[6:0];
            wmt_write_update_val_s3 = 1'b1;
            wmt_write_update_way_s3 = tagcheck_way_s3;
            wmt_write_inval_val_s3 = 1'b1;
        end
    endcase
    
    
    
    
    
    
    
    
    wmt_write_update_mask_s3[4*((2+0)+1)-1:0] = 0;
    if (wmt_write_update_val_s3 == 1'b1)
    begin
        
        
        
        
        
        
        
        
        
  if (l1_replacement_way_s3 == 0)
      wmt_write_update_mask_s3[(0+1)*((2+0)+1)-1 -: ((2+0)+1)] = {((2+0)+1){1'b1}};
  if (l1_replacement_way_s3 == 1)
      wmt_write_update_mask_s3[(1+1)*((2+0)+1)-1 -: ((2+0)+1)] = {((2+0)+1){1'b1}};
  if (l1_replacement_way_s3 == 2)
      wmt_write_update_mask_s3[(2+1)*((2+0)+1)-1 -: ((2+0)+1)] = {((2+0)+1){1'b1}};
  if (l1_replacement_way_s3 == 3)
      wmt_write_update_mask_s3[(3+1)*((2+0)+1)-1 -: ((2+0)+1)] = {((2+0)+1){1'b1}};
    end
    
                                                        
                                                        
                                                        
    
    
    
    
    
    
    
    
    wmt_write_inval_mask_s3[4*((2+0)+1)-1:0] = 0;
    if (wmt_write_inval_val_s3 == 1'b1)
    begin
        
        
        
        
        
  wmt_write_inval_mask_s3[(0+1)*((2+0)+1)-1 -: ((2+0)+1)] = {((2+0)+1){wmt_compare_mask_s3[0]}};
  wmt_write_inval_mask_s3[(1+1)*((2+0)+1)-1 -: ((2+0)+1)] = {((2+0)+1){wmt_compare_mask_s3[1]}};
  wmt_write_inval_mask_s3[(2+1)*((2+0)+1)-1 -: ((2+0)+1)] = {((2+0)+1){wmt_compare_mask_s3[2]}};
  wmt_write_inval_mask_s3[(3+1)*((2+0)+1)-1 -: ((2+0)+1)] = {((2+0)+1){wmt_compare_mask_s3[3]}};
    end
    wmt_write_update_data_s3 = wmt_write_update_way_s3;
    
    wmt_write_mask_s3[4*((2+0)+1)-1:0] = wmt_write_inval_mask_s3 | wmt_write_update_mask_s3;
    wmt_write_data_s3[4*((2+0)+1)-1:0] = {4{{1'b1,wmt_write_update_data_s3}}} & wmt_write_update_mask_s3;
    
    
    
    l15_wmt_write_val_s3 = wmt_write_val_s3 && val_s3;
    l15_wmt_write_index_s3 = wmt_write_index_s3;
    l15_wmt_write_mask_s3 = wmt_write_mask_s3;
    l15_wmt_write_data_s3 = wmt_write_data_s3;
end
reg lru_eviction_matched_st1_s3;
reg lru_eviction_matched_st2_s3;
reg tagcheck_matched_st1_s3;
reg tagcheck_matched_st2_s3;
reg s3_mshr_val_s3;
reg [3-1:0] s3_mshr_write_type_s3;
reg [2-1:0] s3_mshr_update_state_s3;
reg [2-1:0] s3_mshr_write_mshrid_s3;
reg [1:0] s3_mshr_update_way_s3;
reg [0:0] s3_mshr_write_threadid_s3;
always @ *
begin
    s3_mshr_val_s3 = 0;
    s3_mshr_write_type_s3 = 0;
    s3_mshr_write_mshrid_s3 = 0;
    s3_mshr_update_state_s3 = 0;
    s3_mshr_update_way_s3 = 0;
    s3_mshr_write_threadid_s3[0:0] = threadid_s3[0:0];
    case (s3_mshr_operation_s3)
        3'd1:
        begin
            s3_mshr_val_s3 = val_s3;
            s3_mshr_write_type_s3 = 3'b010;
            s3_mshr_write_mshrid_s3 = mshrid_s3;
        end
        3'd2:
        begin
            s3_mshr_val_s3 = val_s3 && tagcheck_state_mes_s3;
            s3_mshr_write_type_s3 = 3'b010;
            s3_mshr_write_mshrid_s3 = mshrid_s3;
        end
        3'd3:
        begin
            s3_mshr_val_s3 = val_s3;
            s3_mshr_write_type_s3 = tagcheck_state_me_s3 ?  3'b010 :
                                                                            3'b011;
            s3_mshr_write_mshrid_s3 = mshrid_s3;
            s3_mshr_update_state_s3 = tagcheck_state_mes_s3 ?
                                                    2'b01 : 2'b10;
            s3_mshr_update_way_s3 = tagcheck_way_s3;
        end
        3'd4:
        begin
            s3_mshr_val_s3 = val_s3 && stbuf_compare_match_val_s3;
            s3_mshr_write_type_s3 = 3'b011;
            
            s3_mshr_update_state_s3 = 2'b10;
            
            s3_mshr_write_threadid_s3[0:0] = stbuf_compare_threadid_s3[0:0];
        end
        3'd5:
        begin
            s3_mshr_val_s3 = val_s3 && stbuf_compare_lru_match_val_s3;
            s3_mshr_write_type_s3 = 3'b011;
            
            s3_mshr_update_state_s3 = 2'b10;
            s3_mshr_write_threadid_s3[0:0] = stbuf_compare_lru_threadid_s3[0:0];
            
        end
        3'd6:
        begin
            s3_mshr_val_s3 = val_s3;
            s3_mshr_write_type_s3 = 3'b011;
            
            s3_mshr_update_state_s3 = 2'b11;
            
            
        end
    endcase
    
    pipe_mshr_val_s3 = s3_mshr_val_s3;
    pipe_mshr_op_s3 = s3_mshr_write_type_s3;
    pipe_mshr_mshrid_s3 = s3_mshr_write_mshrid_s3;
    pipe_mshr_threadid_s3[0:0] = s3_mshr_write_threadid_s3[0:0];
    pipe_mshr_write_update_state_s3 = s3_mshr_update_state_s3;
    pipe_mshr_write_update_way_s3 = s3_mshr_update_way_s3;
end
reg cpx_req_val_s3;
reg [4-1:0] cpx_type_s3;
reg cpx_invalidate_l1_s3;
reg [1:0] cpx_inval_way_s3;
reg [3-1:0] cpx_data_source_s3;
reg cpx_atomic_bit_s3;
reg cpx_icache_inval_s3;
always @ *
begin
    cpx_req_val_s3 = 0;
    cpx_type_s3 = 0;
    cpx_invalidate_l1_s3 = 0;
    
    cpx_inval_way_s3 = 0;
    cpx_data_source_s3 = 0;
    cpx_atomic_bit_s3 = 0;
    cpx_icache_inval_s3 = 0;
    case(cpx_operation_s3)
        5'd14:
        begin
            cpx_req_val_s3 = 1'b1;
            cpx_type_s3 = 4'b0011;
            cpx_icache_inval_s3 = 1;
        end
        5'd19:
        begin
            cpx_req_val_s3 = 1'b1;
            cpx_type_s3 = 4'b0011;
            cpx_invalidate_l1_s3 = 1;
            cpx_inval_way_s3 = wmt_compare_match_way_s3;
        end
        5'd1:
        begin
            cpx_req_val_s3 = tagcheck_state_mes_s3 && wmt_compare_match_s3;
            cpx_type_s3 = 4'b0011;
            cpx_invalidate_l1_s3 = 1;
            cpx_inval_way_s3 = wmt_compare_match_way_s3;
        end
        5'd8:
        begin
            cpx_req_val_s3 = lru_state_mes_s3 && wmt_compare_match_s3;
            cpx_type_s3 = 4'b0011;
            cpx_invalidate_l1_s3 = 1;
            cpx_inval_way_s3 = wmt_compare_match_way_s3;
        end
        5'd17:
        begin
            cpx_req_val_s3 = flush_state_mes_s3 && wmt_compare_match_s3;
            cpx_type_s3 = 4'b0011;
            cpx_invalidate_l1_s3 = 1;
            cpx_inval_way_s3 = wmt_compare_match_way_s3;
        end
        5'd2:
        begin
            cpx_req_val_s3 = 1'b1;
            cpx_type_s3 = 4'b0000;
            cpx_data_source_s3 = 3'd0;
        end
        5'd3:
        begin
            cpx_req_val_s3 = tagcheck_state_mes_s3;
            cpx_type_s3 = 4'b0000;
            cpx_data_source_s3 = 3'd0;
        end
        5'd4:
        begin
            cpx_req_val_s3 = tagcheck_state_mes_s3;
            cpx_type_s3 = 4'b0000;
            cpx_data_source_s3 = 3'd1;
        end
        5'd5:
        begin
            cpx_req_val_s3 = 1'b1;
            cpx_type_s3 = 4'b0000;
            cpx_data_source_s3 = 3'd2;
        end
        5'd6:
        begin
            cpx_req_val_s3 = 1'b1;
            cpx_type_s3 = 4'b0100;
        end
        5'd20:
        begin
            cpx_req_val_s3 = 1'b1;
            cpx_type_s3 = 4'b1110;
            cpx_data_source_s3 = 3'd5;
            cpx_atomic_bit_s3 = 1;
        end
        5'd11:
        begin
            
            
            
            
            
            cpx_req_val_s3 = 1'b1;
            cpx_invalidate_l1_s3 = wmt_compare_match_s3 && stbuf_compare_match_val_s3;
            cpx_type_s3 = 4'b0100;
            cpx_inval_way_s3 = wmt_compare_match_way_s3;
        end
        5'd7:
        begin
            cpx_req_val_s3 = tagcheck_state_me_s3;
            cpx_type_s3 = 4'b0100;
            cpx_invalidate_l1_s3 = wmt_compare_match_s3;
            cpx_inval_way_s3 = wmt_compare_match_way_s3;
        end
        5'd9:
        begin
            cpx_req_val_s3 = 1'b1;
            cpx_type_s3 = 4'b0001;
            cpx_data_source_s3 = 3'd2;
        end
        5'd10:
        begin
            cpx_req_val_s3 = 1'b1;
            cpx_type_s3 = 4'b1110;
            cpx_data_source_s3 = 3'd2;
            cpx_atomic_bit_s3 = 1;
        end
        5'd12:
        begin
            cpx_req_val_s3 = 1'b1;
            cpx_type_s3 = 4'b0111;
            
        end
        5'd13:
        begin
            cpx_req_val_s3 = 1'b1;
            cpx_type_s3 = 4'b0111;
            cpx_data_source_s3 = 3'd2;
            
        end
        5'd15:
        begin
            cpx_req_val_s3 = 1'b1;
            cpx_type_s3 = 4'b0000;
            cpx_data_source_s3 = 3'd3;
        end
        5'd16:
        begin
            
            cpx_req_val_s3 = 1'b1;
            cpx_type_s3 = 4'b0000;
            cpx_data_source_s3 = 3'd1;
        end
        5'd18:
        begin
            
            cpx_req_val_s3 = 1'b1;
            cpx_type_s3 = 4'b0000;
            cpx_data_source_s3 = 3'd4;
        end
    endcase
    l15_cpxencoder_returntype[3:0] = cpx_type_s3; 
    l15_cpxencoder_val = val_s3 && cpx_req_val_s3 && !cpxencoder_req_staled_s3;
    l15_cpxencoder_l2miss = 0;
    l15_cpxencoder_error[1:0] = 0;
    l15_cpxencoder_noncacheable = 0;
    l15_cpxencoder_threadid = 0;
    l15_cpxencoder_prefetch = 0;
    l15_cpxencoder_f4b = 0;
    l15_cpxencoder_atomic = 0;
    l15_cpxencoder_inval_icache_all_way = 0;
    l15_cpxencoder_inval_dcache_all_way = 0;
    l15_cpxencoder_inval_address_15_4[15:4] = 0;
    l15_cpxencoder_cross_invalidate = 0;
    l15_cpxencoder_cross_invalidate_way[1:0] = 0;
    l15_cpxencoder_inval_dcache_inval = 0;
    l15_cpxencoder_inval_icache_inval = 0;
    l15_cpxencoder_inval_way[1:0] = 0;
    l15_cpxencoder_blockinitstore = 0;
    if (cpx_operation_s3 != 5'd13)
    begin
        l15_cpxencoder_l2miss = l2_miss_s3;
        l15_cpxencoder_error[1:0] = 2'b00; 
        l15_cpxencoder_noncacheable = non_cacheable_s3;
        l15_cpxencoder_threadid = threadid_s3;
        l15_cpxencoder_prefetch = prefetch_s3;
        l15_cpxencoder_f4b = f4b_s3; 
        l15_cpxencoder_atomic = cpx_atomic_bit_s3;
        l15_cpxencoder_inval_icache_all_way = cpx_icache_inval_s3;
        
        l15_cpxencoder_inval_address_15_4[15:4] = address_s3[15:4];
        l15_cpxencoder_cross_invalidate = 0; 
        l15_cpxencoder_cross_invalidate_way[1:0] = 2'b0;
        l15_cpxencoder_inval_dcache_inval = cpx_invalidate_l1_s3; 
        
        l15_cpxencoder_inval_icache_inval = 0; 
        l15_cpxencoder_inval_way[1:0] = cpx_inval_way_s3[1:0];
        l15_cpxencoder_blockinitstore = blockstore_s3 || blockstoreinit_s3;
    end
    l15_cpxencoder_data_0[63:0] = 0;
    l15_cpxencoder_data_1[63:0] = 0;
    l15_cpxencoder_data_2[63:0] = 0;
    l15_cpxencoder_data_3[63:0] = 0;
    case (cpx_data_source_s3)
        3'd5:
        begin
            l15_cpxencoder_data_0[63:0] = ((size_s3 == 3'b011) ?
                {7'b0,(~tagcheck_lrsc_flag_s3),24'b0, 7'b0,(~tagcheck_lrsc_flag_s3),24'b0} :
                {7'b0,(~tagcheck_lrsc_flag_s3),56'b0});
            l15_cpxencoder_data_1[63:0] = ((size_s3 == 3'b011) ?
                {7'b0,(~tagcheck_lrsc_flag_s3),24'b0, 7'b0,(~tagcheck_lrsc_flag_s3),24'b0} :
                {7'b0,(~tagcheck_lrsc_flag_s3),56'b0}); 
        end
        3'd1:
        begin
            l15_cpxencoder_data_0[63:0] = dcache_l15_dout_s3[127:64];
            l15_cpxencoder_data_1[63:0] = dcache_l15_dout_s3[63:0];
        end
        3'd2:
        begin
            l15_cpxencoder_data_0[63:0] = noc2decoder_l15_data_0[63:0];
            l15_cpxencoder_data_1[63:0] = noc2decoder_l15_data_1[63:0];
            l15_cpxencoder_data_2[63:0] = noc2decoder_l15_data_2[63:0];
            l15_cpxencoder_data_3[63:0] = noc2decoder_l15_data_3[63:0];
        end
        3'd3:
        begin
            l15_cpxencoder_data_0[63:0] = config_l15_read_res_data_s3[63:0];
        end
        3'd4:
        begin
            l15_cpxencoder_data_0[63:0] = csm_l15_res_data_s3[63:0];
            l15_cpxencoder_data_1[63:0] = csm_l15_res_data_s3[63:0];
        end
    endcase
end
reg [(14+8+8)-1:0] expanded_hmt_homeid_s3;
always @ *
begin
    expanded_hmt_homeid_s3 = 0;
    
    expanded_hmt_homeid_s3[((14+8+8)-1):(8+8)] = hmt_l15_dout_s3[14 + 8 + 8 - 1 -:  14];
    expanded_hmt_homeid_s3[8+8-1:8] = hmt_l15_dout_s3[8 - 1 -: 8];
    expanded_hmt_homeid_s3[8-1:0] = hmt_l15_dout_s3[8 + 8 - 1 -: 8];
end
reg noc1_req_val_s3;
reg [5-1:0] noc1_type_s3;
reg [2-1:0] noc1_data_source_s3;
reg noc1_homeid_not_required_s3;
reg [2-1:0] noc1_homeid_source_s3;
always @ *
begin
    noc1_req_val_s3 = 0;
    noc1_type_s3 = 0;
    noc1_data_source_s3 = 0;
    noc1_homeid_not_required_s3 = 0;
    creditman_noc1_mispredicted_s3 = 0;
    creditman_noc1_reserve_s3 = 0;
    l15_noc1buffer_req_address = 0;
    noc1_homeid_source_s3 = 0;
    case (noc1_operation_s3)
        5'd8:
        begin
            noc1_req_val_s3 = val_s3 && lru_state_m_s3;
            noc1_type_s3 = 5'd1;
            l15_noc1buffer_req_address = lru_way_address_s3;
            creditman_noc1_mispredicted_s3 = noc1_req_val_s3 ? 0 : val_s3;
            noc1_homeid_source_s3 = 2'd3;
        end
        5'd12:
        begin
            noc1_req_val_s3 = val_s3 && flush_state_m_s3;
            noc1_type_s3 = 5'd1;
            l15_noc1buffer_req_address = flush_way_address_s3;
            creditman_noc1_mispredicted_s3 = noc1_req_val_s3 ? 0 : val_s3;
            noc1_homeid_source_s3 = 2'd3;
        end
        5'd9:
        begin
            noc1_req_val_s3 = val_s3 && tagcheck_state_m_s3;
            noc1_type_s3 = 5'd1;
            l15_noc1buffer_req_address = address_s3;
            creditman_noc1_mispredicted_s3 = noc1_req_val_s3 ? 0 : val_s3;
            noc1_homeid_source_s3 = 2'd3;
        end
        5'd1:
        begin
            noc1_req_val_s3 = val_s3;
            noc1_type_s3 = 5'd2;
            l15_noc1buffer_req_address = address_s3;
            noc1_homeid_source_s3 = 2'd1;
            
        end
        5'd2:
        begin
            noc1_req_val_s3 = val_s3 && !tagcheck_state_mes_s3;
            noc1_type_s3 = 5'd2;
            l15_noc1buffer_req_address = address_s3;
            noc1_homeid_source_s3 = 2'd1;
            creditman_noc1_mispredicted_s3 = noc1_req_val_s3 ? 1'b0 : val_s3;
            creditman_noc1_reserve_s3 = noc1_req_val_s3 ? 1'b1 : 1'b0;
        end
        5'd3:
        begin
            noc1_req_val_s3 = val_s3;
            noc1_type_s3 = 5'd3;
            l15_noc1buffer_req_address = address_s3;
            noc1_homeid_source_s3 = 2'd1;
        end
        5'd5:
        begin
            noc1_req_val_s3 = val_s3;
            noc1_type_s3 = 5'd4;
            noc1_data_source_s3 = 2'd1;
            l15_noc1buffer_req_address = address_s3;
            noc1_homeid_source_s3 = 2'd1;
        end
        5'd4:
        begin
            noc1_req_val_s3 = val_s3 && ((tagcheck_state_s3 == 2'd1) || (tagcheck_state_s3 == 2'd0));
            noc1_type_s3 = (tagcheck_state_s3 == 2'd1) ? 5'd5 :
                                                                        5'd6;
            noc1_data_source_s3 = 2'd1;
            l15_noc1buffer_req_address = address_s3;
            noc1_homeid_source_s3 = 2'd1;
            creditman_noc1_mispredicted_s3 = noc1_req_val_s3 ? 1'b0 : val_s3;
            creditman_noc1_reserve_s3 = noc1_req_val_s3 ? 1'b1 : 1'b0;
        end
        5'd21:
        begin
            noc1_req_val_s3 = val_s3;
            noc1_type_s3 = 5'd18;
            
            l15_noc1buffer_req_address = address_s3;
            noc1_homeid_source_s3 = 2'd1;
            creditman_noc1_reserve_s3 = val_s3;
        end
        5'd6:
        begin
            noc1_req_val_s3 = val_s3;
            noc1_type_s3 = 5'd7;
            noc1_data_source_s3 = 2'd2;
            l15_noc1buffer_req_address = address_s3;
            noc1_homeid_source_s3 = 2'd1;
        end
        5'd7:
        begin
            noc1_req_val_s3 = val_s3;
            noc1_type_s3 = 5'd8;
            noc1_data_source_s3 = 2'd1;
            l15_noc1buffer_req_address = address_s3;
            noc1_homeid_source_s3 = 2'd1;
        end
        5'd13:
        begin
            noc1_req_val_s3 = val_s3;
            noc1_type_s3 = 5'd10;
            noc1_data_source_s3 = 2'd1;
            l15_noc1buffer_req_address = address_s3;
            noc1_homeid_source_s3 = 2'd1;
        end
        5'd14:
        begin
            noc1_req_val_s3 = val_s3;
            noc1_type_s3 = 5'd11;
            noc1_data_source_s3 = 2'd1;
            l15_noc1buffer_req_address = address_s3;
            noc1_homeid_source_s3 = 2'd1;
        end
        5'd15:
        begin
            noc1_req_val_s3 = val_s3;
            noc1_type_s3 = 5'd12;
            noc1_data_source_s3 = 2'd1;
            l15_noc1buffer_req_address = address_s3;
            noc1_homeid_source_s3 = 2'd1;
        end
        5'd16:
        begin
            noc1_req_val_s3 = val_s3;
            noc1_type_s3 = 5'd13;
            noc1_data_source_s3 = 2'd1;
            l15_noc1buffer_req_address = address_s3;
            noc1_homeid_source_s3 = 2'd1;
        end
        5'd17:
        begin
            noc1_req_val_s3 = val_s3;
            noc1_type_s3 = 5'd14;
            noc1_data_source_s3 = 2'd1;
            l15_noc1buffer_req_address = address_s3;
            noc1_homeid_source_s3 = 2'd1;
        end
        5'd18:
        begin
            noc1_req_val_s3 = val_s3;
            noc1_type_s3 = 5'd15;
            noc1_data_source_s3 = 2'd1;
            l15_noc1buffer_req_address = address_s3;
            noc1_homeid_source_s3 = 2'd1;
        end
        5'd19:
        begin
            noc1_req_val_s3 = val_s3;
            noc1_type_s3 = 5'd16;
            noc1_data_source_s3 = 2'd1;
            l15_noc1buffer_req_address = address_s3;
            noc1_homeid_source_s3 = 2'd1;
        end
        5'd20:
        begin
            noc1_req_val_s3 = val_s3;
            noc1_type_s3 = 5'd17;
            noc1_data_source_s3 = 2'd1;
            l15_noc1buffer_req_address = address_s3;
            noc1_homeid_source_s3 = 2'd1;
        end
        5'd10:
        begin
            noc1_req_val_s3 = val_s3;
            noc1_type_s3 = 5'd9;
            noc1_data_source_s3 = 2'd1;
            noc1_homeid_not_required_s3 = 1'b1;
        end
    endcase
    l15_noc1buffer_req_val = noc1_req_val_s3 && !noc1encoder_req_staled_s3;
    l15_noc1buffer_req_type = noc1_type_s3;
    l15_noc1buffer_req_threadid = threadid_s3;
    l15_noc1buffer_req_mshrid = mshrid_s3;
    l15_noc1buffer_req_non_cacheable = non_cacheable_s3;
    l15_noc1buffer_req_size = size_s3;
    l15_noc1buffer_req_prefetch = prefetch_s3;
    
    
    l15_noc1buffer_req_data_0[63:0] = 0;
    l15_noc1buffer_req_data_1[63:0] = 0;
    case (noc1_data_source_s3)
        2'd1:
        begin
            l15_noc1buffer_req_data_0[63:0] = pcxdecoder_l15_data[63:0];
            
        end
        2'd2:
        begin
            l15_noc1buffer_req_data_0[63:0] = pcxdecoder_l15_data[63:0];
            l15_noc1buffer_req_data_1[63:0] = pcxdecoder_l15_data_next_entry[63:0];
        end
    endcase
    
    l15_noc1buffer_req_csm_ticket = csm_ticket_s3;
    l15_noc1buffer_req_homeid = 0;
    l15_noc1buffer_req_homeid_val = 0;
    case (noc1_homeid_source_s3)
        2'd1:
        begin
            l15_noc1buffer_req_homeid = csm_l15_res_data_s3;
            l15_noc1buffer_req_homeid_val = csm_l15_res_val_s3;
        end
        2'd3:
        begin
            l15_noc1buffer_req_homeid = expanded_hmt_homeid_s3;
            l15_noc1buffer_req_homeid_val = 1'b1;
        end
    endcase
    l15_noc1buffer_req_homeid_val = l15_noc1buffer_req_homeid_val || noc1_homeid_not_required_s3;
    l15_noc1buffer_req_csm_data = csm_pcx_data_s3; 
end
reg noc3_req_val_s3;
reg [3-1:0] noc3_type_s3;
reg noc3_with_data_s3;
reg [39:0] noc3_address_s3;
reg [2-1:0] noc3_homeid_source_s3;
always @ *
begin
    noc3_req_val_s3 = 0;
    noc3_type_s3 = 0;
    noc3_with_data_s3 = 0;
    noc3_address_s3 = 0;
    noc3_homeid_source_s3 = 0;
    case (noc3_operations_s3)
        4'd5:
        begin
            noc3_req_val_s3 = val_s3 && tagcheck_state_m_s3;
            noc3_type_s3 = 3'd1;
            noc3_with_data_s3 = 1;
            noc3_address_s3 = address_s3;
            noc3_homeid_source_s3 = 2'd3;
        end
        4'd6:
        begin
            noc3_req_val_s3 = val_s3 && lru_state_m_s3;
            noc3_type_s3 = 3'd1;
            noc3_with_data_s3 = 1;
            noc3_address_s3 = lru_way_address_s3;
            noc3_homeid_source_s3 = 2'd3;
        end
        4'd8:
        begin
            noc3_req_val_s3 = val_s3 && flush_state_m_s3;
            noc3_type_s3 = 3'd1;
            noc3_with_data_s3 = 1;
            noc3_address_s3 = flush_way_address_s3;
            noc3_homeid_source_s3 = 2'd3;
        end
        4'd1:
        begin
            noc3_req_val_s3 = val_s3;
            noc3_type_s3 = 3'd2;
            noc3_with_data_s3 = tagcheck_state_m_s3;
            noc3_address_s3 = address_s3;
            noc3_homeid_source_s3 = 2'd2;
        end
        4'd2:
        begin
            noc3_req_val_s3 = val_s3 && (tagcheck_state_m_s3);
            noc3_type_s3 = 3'd2;
            noc3_with_data_s3 = 1;
            noc3_address_s3 = address_s3;
            noc3_homeid_source_s3 = 2'd2;
        end
        4'd3:
        begin
            noc3_req_val_s3 = val_s3;
            noc3_type_s3 = 3'd3;
            noc3_with_data_s3 = tagcheck_state_m_s3;
            noc3_address_s3 = address_s3;
            noc3_homeid_source_s3 = 2'd2;
        end
        4'd4:
        begin
            noc3_req_val_s3 = val_s3 && (tagcheck_state_m_s3);
            noc3_type_s3 = 3'd3;
            noc3_with_data_s3 = 1;
            noc3_address_s3 = address_s3;
            noc3_homeid_source_s3 = 2'd2;
        end
        4'd7:
        begin
            noc3_req_val_s3 = val_s3;
            noc3_type_s3 = 3'd4;
            noc3_address_s3 = address_s3;
            noc3_homeid_source_s3 = 2'd2;
        end
    endcase
    l15_noc3encoder_req_val = noc3_req_val_s3 && !noc3encoder_req_staled_s3;
    l15_noc3encoder_req_type = noc3_type_s3;
    l15_noc3encoder_req_data_0 = dcache_l15_dout_s3[127:64];
    l15_noc3encoder_req_data_1 = dcache_l15_dout_s3[63:0];
    l15_noc3encoder_req_mshrid = mshrid_s3;
    l15_noc3encoder_req_sequenceid = cache_index_s3[1:0];
    l15_noc3encoder_req_threadid = threadid_s3[0:0];
    l15_noc3encoder_req_address[39:0] = noc3_address_s3[39:0];
    l15_noc3encoder_req_with_data = noc3_with_data_s3;
    l15_noc3encoder_req_was_inval = predecode_noc2_inval_s3;
    l15_noc3encoder_req_fwdack_vector = predecode_fwd_subcacheline_vector_s3;
    l15_noc3encoder_req_homeid = 0;
    
    
    
    case (noc3_homeid_source_s3)
        2'd2:
            l15_noc3encoder_req_homeid = noc2_src_homeid_s3[(14+8+8)-1:0];
        2'd3:
            
            
                
                l15_noc3encoder_req_homeid = expanded_hmt_homeid_s3;
            
    endcase
end
endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
module l15_priority_encoder_1(
    input wire [1:0] data_in,
    output wire [0:0] data_out,
    output wire [1:0] data_out_mask,
    output wire nonzero_out
);
assign data_out = data_in[0] ? 1'b0 : 1'b1;
assign data_out_mask = data_in[0] ? 2'b10 : 2'b01;
assign nonzero_out = | (data_in[1:0]);
endmodule
module l15_priority_encoder_2(
    input wire [3:0] data_in,
    output wire [1:0] data_out,
    output wire [3:0] data_out_mask,
    output wire nonzero_out
);
wire [0:0] data_low;
wire [0:0] data_high;
wire [1:0] data_low_mask;
wire [1:0] data_high_mask;
wire nonzero_low;
wire nonzero_high;
l15_priority_encoder_1 encoder_high_1 (.data_in(data_in[3:2]), .data_out(data_high), .data_out_mask(data_high_mask), .nonzero_out(nonzero_high));
l15_priority_encoder_1 encoder_low_1(.data_in(data_in[1:0]), .data_out(data_low), .data_out_mask(data_low_mask), .nonzero_out(nonzero_low));
assign data_out = nonzero_low ? {1'b0, data_low} : {1'b1, data_high};
assign data_out_mask = nonzero_low ? {{2{1'b1}}, data_low_mask} : {data_high_mask,{2{1'b1}}};
assign nonzero_out = nonzero_low | nonzero_high;
endmodule
module l15_priority_encoder_3(
    input wire [7:0] data_in,
    output wire [2:0] data_out,
    output wire [7:0] data_out_mask,
    output wire nonzero_out
);
wire [1:0] data_low;
wire [1:0] data_high;
wire [3:0] data_low_mask;
wire [3:0] data_high_mask;
wire nonzero_low;
wire nonzero_high;
l15_priority_encoder_2 encoder_high_2 (.data_in(data_in[7:4]), .data_out(data_high), .data_out_mask(data_high_mask), .nonzero_out(nonzero_high));
l15_priority_encoder_2 encoder_low_2(.data_in(data_in[3:0]), .data_out(data_low), .data_out_mask(data_low_mask), .nonzero_out(nonzero_low));
assign data_out = nonzero_low ? {1'b0, data_low} : {1'b1, data_high};
assign data_out_mask = nonzero_low ? {{4{1'b1}}, data_low_mask} : {data_high_mask,{4{1'b1}}};
assign nonzero_out = nonzero_low | nonzero_high;
endmodule
module l15_priority_encoder_4(
    input wire [15:0] data_in,
    output wire [3:0] data_out,
    output wire [15:0] data_out_mask,
    output wire nonzero_out
);
wire [2:0] data_low;
wire [2:0] data_high;
wire [7:0] data_low_mask;
wire [7:0] data_high_mask;
wire nonzero_low;
wire nonzero_high;
l15_priority_encoder_3 encoder_high_3 (.data_in(data_in[15:8]), .data_out(data_high), .data_out_mask(data_high_mask), .nonzero_out(nonzero_high));
l15_priority_encoder_3 encoder_low_3(.data_in(data_in[7:0]), .data_out(data_low), .data_out_mask(data_low_mask), .nonzero_out(nonzero_low));
assign data_out = nonzero_low ? {1'b0, data_low} : {1'b1, data_high};
assign data_out_mask = nonzero_low ? {{8{1'b1}}, data_low_mask} : {data_high_mask,{8{1'b1}}};
assign nonzero_out = nonzero_low | nonzero_high;
endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
 
module noc1buffer(
   input wire clk,
   input wire rst_n,
   input wire [63:0] l15_noc1buffer_req_data_0,
   input wire [63:0] l15_noc1buffer_req_data_1,
   input wire l15_noc1buffer_req_val,
   input wire [5-1:0] l15_noc1buffer_req_type,
   input wire [2-1:0] l15_noc1buffer_req_mshrid,
   input wire [0:0] l15_noc1buffer_req_threadid,
   input wire [39:0] l15_noc1buffer_req_address,
   input wire l15_noc1buffer_req_non_cacheable,
   input wire [3-1:0] l15_noc1buffer_req_size,
   input wire l15_noc1buffer_req_prefetch,
   
   
   input wire [3-1:0] l15_noc1buffer_req_csm_ticket,
   input wire [(14+8+8)-1:0] l15_noc1buffer_req_homeid,
   input wire l15_noc1buffer_req_homeid_val,
   input wire [33-1:0] l15_noc1buffer_req_csm_data,
   input wire noc1encoder_noc1buffer_req_ack,
   
   input wire [(14+8+8)-1:0] csm_l15_read_res_data,
   input wire csm_l15_read_res_val,
   output reg [63:0] noc1buffer_noc1encoder_req_data_0,
   output reg [63:0] noc1buffer_noc1encoder_req_data_1,
   output reg noc1buffer_noc1encoder_req_val,
   output reg [5-1:0] noc1buffer_noc1encoder_req_type,
   output reg [2-1:0] noc1buffer_noc1encoder_req_mshrid,
   output reg [0:0] noc1buffer_noc1encoder_req_threadid,
   output reg [39:0] noc1buffer_noc1encoder_req_address,
   output reg noc1buffer_noc1encoder_req_non_cacheable,
   output reg [3-1:0] noc1buffer_noc1encoder_req_size,
   output reg noc1buffer_noc1encoder_req_prefetch,
   
   
   output reg [(14+8+8)-1:0] noc1buffer_noc1encoder_req_homeid,
   output reg [10-1:0] noc1buffer_noc1encoder_req_csm_sdid,
   output reg [6-1:0] noc1buffer_noc1encoder_req_csm_lsid,
   
   output reg [3-1:0] l15_csm_read_ticket,
   output reg [3-1:0] l15_csm_clear_ticket,
   output reg l15_csm_clear_ticket_val,
   
   output reg noc1buffer_mshr_homeid_write_val_s4,
   output reg [2-1:0] noc1buffer_mshr_homeid_write_mshrid_s4,
   output reg [0:0] noc1buffer_mshr_homeid_write_threadid_s4,
   output reg [(14+8+8)-1:0] noc1buffer_mshr_homeid_write_data_s4,
   
   output reg noc1buffer_l15_req_sent,
   output reg [2-1:0] noc1buffer_l15_req_data_sent
);
reg [0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + (14+8+8) - 1 + 1 + 1 - 1 + 1 + 10 - 1 + 1 + 6 - 1 + 1-1:0] command_buffer [0:8-1];
reg [63:0] data_buffer [0:2-1];
reg [0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + (14+8+8) - 1 + 1 + 1 - 1 + 1 + 10 - 1 + 1 + 6 - 1 + 1-1:0] command_buffer_next [0:8-1];
reg [63:0] data_buffer_next [0:2-1];
reg command_buffer_val [0:8-1];
reg command_buffer_val_next [0:8-1];
reg [3-1:0] command_wrindex;
reg [3-1:0] command_wrindex_next;
reg [3-1:0] command_rdindex;
reg [3-1:0] command_rdindex_next;
reg [3-1:0] command_rdindex_plus1;
reg [1-1:0] data_wrindex;
reg [1-1:0] data_wrindex_next;
reg [1-1:0] data_wrindex_plus_1;
reg [1-1:0] data_wrindex_plus_2;
reg [1-1:0] data_rdindex;
reg [1-1:0] data_rdindex_plus1;
always @ (posedge clk)
begin
   if (!rst_n)
   begin
      command_buffer[0] <= 0;
command_buffer_val[0] <= 0;
command_buffer[1] <= 0;
command_buffer_val[1] <= 0;
command_buffer[2] <= 0;
command_buffer_val[2] <= 0;
command_buffer[3] <= 0;
command_buffer_val[3] <= 0;
command_buffer[4] <= 0;
command_buffer_val[4] <= 0;
command_buffer[5] <= 0;
command_buffer_val[5] <= 0;
command_buffer[6] <= 0;
command_buffer_val[6] <= 0;
command_buffer[7] <= 0;
command_buffer_val[7] <= 0;
data_buffer[0] <= 0;
data_buffer[1] <= 0;
      data_wrindex <= 0;
      command_wrindex <= 0;
      command_rdindex <= 0;
   end
   else
   begin
      
      
      
      
      
      
      
      
      
      command_buffer[0] <= command_buffer_next[0];
command_buffer_val[0] <= command_buffer_val_next[0];
command_buffer[1] <= command_buffer_next[1];
command_buffer_val[1] <= command_buffer_val_next[1];
command_buffer[2] <= command_buffer_next[2];
command_buffer_val[2] <= command_buffer_val_next[2];
command_buffer[3] <= command_buffer_next[3];
command_buffer_val[3] <= command_buffer_val_next[3];
command_buffer[4] <= command_buffer_next[4];
command_buffer_val[4] <= command_buffer_val_next[4];
command_buffer[5] <= command_buffer_next[5];
command_buffer_val[5] <= command_buffer_val_next[5];
command_buffer[6] <= command_buffer_next[6];
command_buffer_val[6] <= command_buffer_val_next[6];
command_buffer[7] <= command_buffer_next[7];
command_buffer_val[7] <= command_buffer_val_next[7];
data_buffer[0] <= data_buffer_next[0];
data_buffer[1] <= data_buffer_next[1];
      data_wrindex <= data_wrindex_next;
      command_wrindex <= command_wrindex_next;
      command_rdindex <= command_rdindex_next;
   end
end
always @ *
begin
   command_buffer_next[0] = command_buffer[0];
command_buffer_next[1] = command_buffer[1];
command_buffer_next[2] = command_buffer[2];
command_buffer_next[3] = command_buffer[3];
command_buffer_next[4] = command_buffer[4];
command_buffer_next[5] = command_buffer[5];
command_buffer_next[6] = command_buffer[6];
command_buffer_next[7] = command_buffer[7];
data_buffer_next[0] = data_buffer[0];
data_buffer_next[1] = data_buffer[1];
   command_wrindex_next = command_wrindex;
   data_wrindex_next = data_wrindex;
   data_wrindex_plus_1 = data_wrindex + 1;
   data_wrindex_plus_2 = data_wrindex + 2;
   if (l15_noc1buffer_req_val)
   begin
      command_buffer_next[command_wrindex][0 + 5 - 1:0] = l15_noc1buffer_req_type;
      command_buffer_next[command_wrindex][0 + 5 - 1 + 1 + 2 - 1:0 + 5 - 1 + 1] = l15_noc1buffer_req_mshrid;
      command_buffer_next[command_wrindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1:0 + 5 - 1 + 1 + 2 - 1 + 1] = l15_noc1buffer_req_threadid;
      command_buffer_next[command_wrindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1:0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1] = l15_noc1buffer_req_address;
      command_buffer_next[command_wrindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1:0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1] = l15_noc1buffer_req_non_cacheable;
      command_buffer_next[command_wrindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1:0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1] = l15_noc1buffer_req_size;
      command_buffer_next[command_wrindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1:0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1] = l15_noc1buffer_req_prefetch;
      
      
      command_buffer_next[command_wrindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1:0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1] = data_wrindex;
      command_buffer_next[command_wrindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1 + 3 - 1:0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1] = l15_noc1buffer_req_csm_ticket;
      command_buffer_next[command_wrindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + (14+8+8) - 1:0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1] = l15_noc1buffer_req_homeid;
      command_buffer_next[command_wrindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + (14+8+8) - 1 + 1 + 1 - 1:0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + (14+8+8) - 1 + 1] = l15_noc1buffer_req_homeid_val;
      command_buffer_next[command_wrindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + (14+8+8) - 1 + 1 + 1 - 1 + 1 + 10 - 1:0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + (14+8+8) - 1 + 1 + 1 - 1 + 1] = l15_noc1buffer_req_csm_data[15:6];
      command_buffer_next[command_wrindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + (14+8+8) - 1 + 1 + 1 - 1 + 1 + 10 - 1 + 1 + 6 - 1:0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + (14+8+8) - 1 + 1 + 1 - 1 + 1 + 10 - 1 + 1] = l15_noc1buffer_req_csm_data[5:0];
      command_wrindex_next = command_wrindex + 1;
      if (l15_noc1buffer_req_type == 5'd7)
      begin
         data_buffer_next[data_wrindex] = l15_noc1buffer_req_data_0;
         data_buffer_next[data_wrindex_plus_1] = l15_noc1buffer_req_data_1;
         data_wrindex_next = data_wrindex_plus_2;
      end
      else if (l15_noc1buffer_req_type == 5'd8 ||
               l15_noc1buffer_req_type == 5'd10 ||
               l15_noc1buffer_req_type == 5'd11 ||
               l15_noc1buffer_req_type == 5'd12 ||
               l15_noc1buffer_req_type == 5'd13 ||
               l15_noc1buffer_req_type == 5'd14 ||
               l15_noc1buffer_req_type == 5'd15 ||
               l15_noc1buffer_req_type == 5'd16 ||
               l15_noc1buffer_req_type == 5'd17 ||
               l15_noc1buffer_req_type == 5'd9 ||
               l15_noc1buffer_req_type == 5'd4)
      begin
         data_buffer_next[data_wrindex] = l15_noc1buffer_req_data_0;
         data_wrindex_next = data_wrindex_plus_1;
      end
   end
end
reg [(14+8+8)-1:0] homeid;
reg homeid_val;
always @ *
begin
   
                                                
   noc1buffer_noc1encoder_req_type = command_buffer[command_rdindex][0 + 5 - 1:0];
   noc1buffer_noc1encoder_req_mshrid = command_buffer[command_rdindex][0 + 5 - 1 + 1 + 2 - 1:0 + 5 - 1 + 1];
   noc1buffer_noc1encoder_req_threadid = command_buffer[command_rdindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1:0 + 5 - 1 + 1 + 2 - 1 + 1];
   noc1buffer_noc1encoder_req_address = command_buffer[command_rdindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1:0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1];
   noc1buffer_noc1encoder_req_non_cacheable = command_buffer[command_rdindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1:0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1];
   noc1buffer_noc1encoder_req_size = command_buffer[command_rdindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1:0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1];
   noc1buffer_noc1encoder_req_prefetch = command_buffer[command_rdindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1:0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1];
   
   
   noc1buffer_noc1encoder_req_csm_sdid = command_buffer[command_rdindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + (14+8+8) - 1 + 1 + 1 - 1 + 1 + 10 - 1:0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + (14+8+8) - 1 + 1 + 1 - 1 + 1];
   noc1buffer_noc1encoder_req_csm_lsid = command_buffer[command_rdindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + (14+8+8) - 1 + 1 + 1 - 1 + 1 + 10 - 1 + 1 + 6 - 1:0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + (14+8+8) - 1 + 1 + 1 - 1 + 1 + 10 - 1 + 1];
   data_rdindex = command_buffer[command_rdindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1:0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1];
   data_rdindex_plus1 = data_rdindex + 1;
   noc1buffer_noc1encoder_req_data_0 = data_buffer[data_rdindex];
   noc1buffer_noc1encoder_req_data_1 = data_buffer[data_rdindex_plus1];
   noc1buffer_noc1encoder_req_homeid = homeid;
   noc1buffer_noc1encoder_req_val = command_buffer_val[command_rdindex] && homeid_val;
end
reg [(14+8+8)-1:0] cached_homeid;
reg cached_homeid_val;
reg [(14+8+8)-1:0] fetch_homeid;
reg fetch_homeid_val;
   
   
   
always @ *
begin
   cached_homeid_val = command_buffer[command_rdindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + (14+8+8) - 1 + 1 + 1 - 1:0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + (14+8+8) - 1 + 1];
   cached_homeid = command_buffer[command_rdindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + (14+8+8) - 1:0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1];
   fetch_homeid_val = csm_l15_read_res_val;
   fetch_homeid = csm_l15_read_res_data;
   homeid_val = cached_homeid_val | fetch_homeid_val;
   homeid = cached_homeid_val ? cached_homeid : fetch_homeid;
   
   l15_csm_read_ticket = command_buffer[command_rdindex][0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1 + 3 - 1:0 + 5 - 1 + 1 + 2 - 1 + 1 + 1 - 1 + 1 + 40 - 1 + 1 + 1 - 1 + 1 + 3 - 1 + 1 + 1 - 1 + 1 + 1 - 1 + 1]; 
   l15_csm_clear_ticket = l15_csm_read_ticket;
   l15_csm_clear_ticket_val = noc1encoder_noc1buffer_req_ack; 
   
   noc1buffer_mshr_homeid_write_val_s4 = (noc1buffer_noc1encoder_req_mshrid == 2'd2 || noc1buffer_noc1encoder_req_mshrid == 2'd3) &&
                                    noc1encoder_noc1buffer_req_ack;
   noc1buffer_mshr_homeid_write_mshrid_s4 = noc1buffer_noc1encoder_req_mshrid;
   noc1buffer_mshr_homeid_write_threadid_s4 = noc1buffer_noc1encoder_req_threadid;
   noc1buffer_mshr_homeid_write_data_s4 = homeid;
end
always @ *
begin
   
   if (l15_noc1buffer_req_val && (command_wrindex == 0))
      command_buffer_val_next[0] = 1'b1;
   else if (noc1encoder_noc1buffer_req_ack && (command_rdindex == 0))
      command_buffer_val_next[0] = 1'b0;
   else
      command_buffer_val_next[0] = command_buffer_val[0];
   
   if (l15_noc1buffer_req_val && (command_wrindex == 1))
      command_buffer_val_next[1] = 1'b1;
   else if (noc1encoder_noc1buffer_req_ack && (command_rdindex == 1))
      command_buffer_val_next[1] = 1'b0;
   else
      command_buffer_val_next[1] = command_buffer_val[1];
   
   if (l15_noc1buffer_req_val && (command_wrindex == 2))
      command_buffer_val_next[2] = 1'b1;
   else if (noc1encoder_noc1buffer_req_ack && (command_rdindex == 2))
      command_buffer_val_next[2] = 1'b0;
   else
      command_buffer_val_next[2] = command_buffer_val[2];
   
   if (l15_noc1buffer_req_val && (command_wrindex == 3))
      command_buffer_val_next[3] = 1'b1;
   else if (noc1encoder_noc1buffer_req_ack && (command_rdindex == 3))
      command_buffer_val_next[3] = 1'b0;
   else
      command_buffer_val_next[3] = command_buffer_val[3];
   
   if (l15_noc1buffer_req_val && (command_wrindex == 4))
      command_buffer_val_next[4] = 1'b1;
   else if (noc1encoder_noc1buffer_req_ack && (command_rdindex == 4))
      command_buffer_val_next[4] = 1'b0;
   else
      command_buffer_val_next[4] = command_buffer_val[4];
   
   if (l15_noc1buffer_req_val && (command_wrindex == 5))
      command_buffer_val_next[5] = 1'b1;
   else if (noc1encoder_noc1buffer_req_ack && (command_rdindex == 5))
      command_buffer_val_next[5] = 1'b0;
   else
      command_buffer_val_next[5] = command_buffer_val[5];
   
   if (l15_noc1buffer_req_val && (command_wrindex == 6))
      command_buffer_val_next[6] = 1'b1;
   else if (noc1encoder_noc1buffer_req_ack && (command_rdindex == 6))
      command_buffer_val_next[6] = 1'b0;
   else
      command_buffer_val_next[6] = command_buffer_val[6];
   
   if (l15_noc1buffer_req_val && (command_wrindex == 7))
      command_buffer_val_next[7] = 1'b1;
   else if (noc1encoder_noc1buffer_req_ack && (command_rdindex == 7))
      command_buffer_val_next[7] = 1'b0;
   else
      command_buffer_val_next[7] = command_buffer_val[7];
   
end
always @ *
begin
   noc1buffer_l15_req_data_sent = 0;
   noc1buffer_l15_req_sent = noc1encoder_noc1buffer_req_ack;
   command_rdindex_plus1 = command_rdindex + 1;
   command_rdindex_next = command_rdindex;
   if (noc1encoder_noc1buffer_req_ack == 1'b1)
   begin
      command_rdindex_next = command_rdindex_plus1;
      case (noc1buffer_noc1encoder_req_type)
         5'd4,
         5'd8,
         5'd10,
         5'd11,
         5'd12,
         5'd13,
         5'd14,
         5'd15,
         5'd16,
         5'd17,
         5'd9:
         begin
            noc1buffer_l15_req_data_sent = 2'd1;
         end
         5'd7:
         begin
            noc1buffer_l15_req_data_sent = 2'd2;
         end
      endcase
   end
end
endmodule
module rf_l15_lrsc_flag(
   input wire clk,
   input wire rst_n,
   input wire read_valid,
   input wire [((9-2))-1:0] read_index,
   input wire write_valid,
   input wire [((9-2))-1:0] write_index,
   input wire [3:0] write_mask,
   input wire [3:0] write_data,
   output wire [3:0] read_data
   );
reg [((9-2))-1:0] read_index_f;
reg [((9-2))-1:0] write_index_f;
reg [3:0] write_data_f;
reg [3:0] write_mask_f;
reg write_valid_f;
reg [3:0] regfile [0:(512/4)-1];
always @ (posedge clk)
begin
   if (!rst_n)
   begin
      read_index_f <= 0;
   end
   else
   if (read_valid)
      read_index_f <= read_index;
   else
      read_index_f <= read_index_f;
end
assign read_data = regfile[read_index_f];
always @ (posedge clk)
begin
   write_valid_f <= write_valid;
   if (write_valid)
   begin
      write_data_f <= write_data;
      write_index_f <= write_index;
      write_mask_f <= write_mask;
   end
end
always @ (posedge clk)
begin
   if (!rst_n)
   begin
      regfile[0] <= 4'b0;
regfile[1] <= 4'b0;
regfile[2] <= 4'b0;
regfile[3] <= 4'b0;
regfile[4] <= 4'b0;
regfile[5] <= 4'b0;
regfile[6] <= 4'b0;
regfile[7] <= 4'b0;
regfile[8] <= 4'b0;
regfile[9] <= 4'b0;
regfile[10] <= 4'b0;
regfile[11] <= 4'b0;
regfile[12] <= 4'b0;
regfile[13] <= 4'b0;
regfile[14] <= 4'b0;
regfile[15] <= 4'b0;
regfile[16] <= 4'b0;
regfile[17] <= 4'b0;
regfile[18] <= 4'b0;
regfile[19] <= 4'b0;
regfile[20] <= 4'b0;
regfile[21] <= 4'b0;
regfile[22] <= 4'b0;
regfile[23] <= 4'b0;
regfile[24] <= 4'b0;
regfile[25] <= 4'b0;
regfile[26] <= 4'b0;
regfile[27] <= 4'b0;
regfile[28] <= 4'b0;
regfile[29] <= 4'b0;
regfile[30] <= 4'b0;
regfile[31] <= 4'b0;
regfile[32] <= 4'b0;
regfile[33] <= 4'b0;
regfile[34] <= 4'b0;
regfile[35] <= 4'b0;
regfile[36] <= 4'b0;
regfile[37] <= 4'b0;
regfile[38] <= 4'b0;
regfile[39] <= 4'b0;
regfile[40] <= 4'b0;
regfile[41] <= 4'b0;
regfile[42] <= 4'b0;
regfile[43] <= 4'b0;
regfile[44] <= 4'b0;
regfile[45] <= 4'b0;
regfile[46] <= 4'b0;
regfile[47] <= 4'b0;
regfile[48] <= 4'b0;
regfile[49] <= 4'b0;
regfile[50] <= 4'b0;
regfile[51] <= 4'b0;
regfile[52] <= 4'b0;
regfile[53] <= 4'b0;
regfile[54] <= 4'b0;
regfile[55] <= 4'b0;
regfile[56] <= 4'b0;
regfile[57] <= 4'b0;
regfile[58] <= 4'b0;
regfile[59] <= 4'b0;
regfile[60] <= 4'b0;
regfile[61] <= 4'b0;
regfile[62] <= 4'b0;
regfile[63] <= 4'b0;
regfile[64] <= 4'b0;
regfile[65] <= 4'b0;
regfile[66] <= 4'b0;
regfile[67] <= 4'b0;
regfile[68] <= 4'b0;
regfile[69] <= 4'b0;
regfile[70] <= 4'b0;
regfile[71] <= 4'b0;
regfile[72] <= 4'b0;
regfile[73] <= 4'b0;
regfile[74] <= 4'b0;
regfile[75] <= 4'b0;
regfile[76] <= 4'b0;
regfile[77] <= 4'b0;
regfile[78] <= 4'b0;
regfile[79] <= 4'b0;
regfile[80] <= 4'b0;
regfile[81] <= 4'b0;
regfile[82] <= 4'b0;
regfile[83] <= 4'b0;
regfile[84] <= 4'b0;
regfile[85] <= 4'b0;
regfile[86] <= 4'b0;
regfile[87] <= 4'b0;
regfile[88] <= 4'b0;
regfile[89] <= 4'b0;
regfile[90] <= 4'b0;
regfile[91] <= 4'b0;
regfile[92] <= 4'b0;
regfile[93] <= 4'b0;
regfile[94] <= 4'b0;
regfile[95] <= 4'b0;
regfile[96] <= 4'b0;
regfile[97] <= 4'b0;
regfile[98] <= 4'b0;
regfile[99] <= 4'b0;
regfile[100] <= 4'b0;
regfile[101] <= 4'b0;
regfile[102] <= 4'b0;
regfile[103] <= 4'b0;
regfile[104] <= 4'b0;
regfile[105] <= 4'b0;
regfile[106] <= 4'b0;
regfile[107] <= 4'b0;
regfile[108] <= 4'b0;
regfile[109] <= 4'b0;
regfile[110] <= 4'b0;
regfile[111] <= 4'b0;
regfile[112] <= 4'b0;
regfile[113] <= 4'b0;
regfile[114] <= 4'b0;
regfile[115] <= 4'b0;
regfile[116] <= 4'b0;
regfile[117] <= 4'b0;
regfile[118] <= 4'b0;
regfile[119] <= 4'b0;
regfile[120] <= 4'b0;
regfile[121] <= 4'b0;
regfile[122] <= 4'b0;
regfile[123] <= 4'b0;
regfile[124] <= 4'b0;
regfile[125] <= 4'b0;
regfile[126] <= 4'b0;
regfile[127] <= 4'b0;
      
   end
   else
   if (write_valid_f)
   begin
      
      regfile[write_index_f] <= (write_data_f & write_mask_f) | (regfile[write_index_f] & ~write_mask_f);
   end
end
endmodule
module rf_l15_lruarray(
   input wire clk,
   input wire rst_n,
   input wire read_valid,
   input wire [((9-2))-1:0] read_index,
   input wire write_valid,
   input wire [((9-2))-1:0] write_index,
   input wire [5:0] write_mask,
   input wire [5:0] write_data,
   output wire [5:0] read_data
   );
reg [((9-2))-1:0] read_index_f;
reg [5:0] regfile [0:(512/4)-1];
always @ (posedge clk)
begin
   if (!rst_n)
   begin
      read_index_f <= 0;
   end
   else
   if (read_valid)
      read_index_f <= read_index;
   else
      read_index_f <= read_index_f;
end
assign read_data = regfile[read_index_f];
always @ (posedge clk)
begin
   if (!rst_n)
   begin
      regfile[0] <= 6'b0;
regfile[1] <= 6'b0;
regfile[2] <= 6'b0;
regfile[3] <= 6'b0;
regfile[4] <= 6'b0;
regfile[5] <= 6'b0;
regfile[6] <= 6'b0;
regfile[7] <= 6'b0;
regfile[8] <= 6'b0;
regfile[9] <= 6'b0;
regfile[10] <= 6'b0;
regfile[11] <= 6'b0;
regfile[12] <= 6'b0;
regfile[13] <= 6'b0;
regfile[14] <= 6'b0;
regfile[15] <= 6'b0;
regfile[16] <= 6'b0;
regfile[17] <= 6'b0;
regfile[18] <= 6'b0;
regfile[19] <= 6'b0;
regfile[20] <= 6'b0;
regfile[21] <= 6'b0;
regfile[22] <= 6'b0;
regfile[23] <= 6'b0;
regfile[24] <= 6'b0;
regfile[25] <= 6'b0;
regfile[26] <= 6'b0;
regfile[27] <= 6'b0;
regfile[28] <= 6'b0;
regfile[29] <= 6'b0;
regfile[30] <= 6'b0;
regfile[31] <= 6'b0;
regfile[32] <= 6'b0;
regfile[33] <= 6'b0;
regfile[34] <= 6'b0;
regfile[35] <= 6'b0;
regfile[36] <= 6'b0;
regfile[37] <= 6'b0;
regfile[38] <= 6'b0;
regfile[39] <= 6'b0;
regfile[40] <= 6'b0;
regfile[41] <= 6'b0;
regfile[42] <= 6'b0;
regfile[43] <= 6'b0;
regfile[44] <= 6'b0;
regfile[45] <= 6'b0;
regfile[46] <= 6'b0;
regfile[47] <= 6'b0;
regfile[48] <= 6'b0;
regfile[49] <= 6'b0;
regfile[50] <= 6'b0;
regfile[51] <= 6'b0;
regfile[52] <= 6'b0;
regfile[53] <= 6'b0;
regfile[54] <= 6'b0;
regfile[55] <= 6'b0;
regfile[56] <= 6'b0;
regfile[57] <= 6'b0;
regfile[58] <= 6'b0;
regfile[59] <= 6'b0;
regfile[60] <= 6'b0;
regfile[61] <= 6'b0;
regfile[62] <= 6'b0;
regfile[63] <= 6'b0;
regfile[64] <= 6'b0;
regfile[65] <= 6'b0;
regfile[66] <= 6'b0;
regfile[67] <= 6'b0;
regfile[68] <= 6'b0;
regfile[69] <= 6'b0;
regfile[70] <= 6'b0;
regfile[71] <= 6'b0;
regfile[72] <= 6'b0;
regfile[73] <= 6'b0;
regfile[74] <= 6'b0;
regfile[75] <= 6'b0;
regfile[76] <= 6'b0;
regfile[77] <= 6'b0;
regfile[78] <= 6'b0;
regfile[79] <= 6'b0;
regfile[80] <= 6'b0;
regfile[81] <= 6'b0;
regfile[82] <= 6'b0;
regfile[83] <= 6'b0;
regfile[84] <= 6'b0;
regfile[85] <= 6'b0;
regfile[86] <= 6'b0;
regfile[87] <= 6'b0;
regfile[88] <= 6'b0;
regfile[89] <= 6'b0;
regfile[90] <= 6'b0;
regfile[91] <= 6'b0;
regfile[92] <= 6'b0;
regfile[93] <= 6'b0;
regfile[94] <= 6'b0;
regfile[95] <= 6'b0;
regfile[96] <= 6'b0;
regfile[97] <= 6'b0;
regfile[98] <= 6'b0;
regfile[99] <= 6'b0;
regfile[100] <= 6'b0;
regfile[101] <= 6'b0;
regfile[102] <= 6'b0;
regfile[103] <= 6'b0;
regfile[104] <= 6'b0;
regfile[105] <= 6'b0;
regfile[106] <= 6'b0;
regfile[107] <= 6'b0;
regfile[108] <= 6'b0;
regfile[109] <= 6'b0;
regfile[110] <= 6'b0;
regfile[111] <= 6'b0;
regfile[112] <= 6'b0;
regfile[113] <= 6'b0;
regfile[114] <= 6'b0;
regfile[115] <= 6'b0;
regfile[116] <= 6'b0;
regfile[117] <= 6'b0;
regfile[118] <= 6'b0;
regfile[119] <= 6'b0;
regfile[120] <= 6'b0;
regfile[121] <= 6'b0;
regfile[122] <= 6'b0;
regfile[123] <= 6'b0;
regfile[124] <= 6'b0;
regfile[125] <= 6'b0;
regfile[126] <= 6'b0;
regfile[127] <= 6'b0;
      
   end
   else
   if (write_valid)
   begin
      regfile[write_index] <= (write_data & write_mask) | (regfile[write_index] & ~write_mask);
   end
end
endmodule
module rf_l15_mesi(
   input wire clk,
   input wire rst_n,
   input wire read_valid,
   input wire [((9-2))-1:0] read_index,
   input wire write_valid,
   input wire [((9-2))-1:0] write_index,
   input wire [7:0] write_mask,
   input wire [7:0] write_data,
   output wire [7:0] read_data
   );
reg [((9-2))-1:0] read_index_f;
reg [((9-2))-1:0] write_index_f;
reg [7:0] write_data_f;
reg [7:0] write_mask_f;
reg write_valid_f;
reg [7:0] regfile [0:(512/4)-1];
always @ (posedge clk)
begin
   if (!rst_n)
   begin
      read_index_f <= 0;
   end
   else
   if (read_valid)
      read_index_f <= read_index;
   else
      read_index_f <= read_index_f;
end
assign read_data = regfile[read_index_f];
always @ (posedge clk)
begin
   write_valid_f <= write_valid;
   if (write_valid)
   begin
      write_data_f <= write_data;
      write_index_f <= write_index;
      write_mask_f <= write_mask;
   end
end
always @ (posedge clk)
begin
   if (!rst_n)
   begin
      regfile[0] <= 8'b0;
regfile[1] <= 8'b0;
regfile[2] <= 8'b0;
regfile[3] <= 8'b0;
regfile[4] <= 8'b0;
regfile[5] <= 8'b0;
regfile[6] <= 8'b0;
regfile[7] <= 8'b0;
regfile[8] <= 8'b0;
regfile[9] <= 8'b0;
regfile[10] <= 8'b0;
regfile[11] <= 8'b0;
regfile[12] <= 8'b0;
regfile[13] <= 8'b0;
regfile[14] <= 8'b0;
regfile[15] <= 8'b0;
regfile[16] <= 8'b0;
regfile[17] <= 8'b0;
regfile[18] <= 8'b0;
regfile[19] <= 8'b0;
regfile[20] <= 8'b0;
regfile[21] <= 8'b0;
regfile[22] <= 8'b0;
regfile[23] <= 8'b0;
regfile[24] <= 8'b0;
regfile[25] <= 8'b0;
regfile[26] <= 8'b0;
regfile[27] <= 8'b0;
regfile[28] <= 8'b0;
regfile[29] <= 8'b0;
regfile[30] <= 8'b0;
regfile[31] <= 8'b0;
regfile[32] <= 8'b0;
regfile[33] <= 8'b0;
regfile[34] <= 8'b0;
regfile[35] <= 8'b0;
regfile[36] <= 8'b0;
regfile[37] <= 8'b0;
regfile[38] <= 8'b0;
regfile[39] <= 8'b0;
regfile[40] <= 8'b0;
regfile[41] <= 8'b0;
regfile[42] <= 8'b0;
regfile[43] <= 8'b0;
regfile[44] <= 8'b0;
regfile[45] <= 8'b0;
regfile[46] <= 8'b0;
regfile[47] <= 8'b0;
regfile[48] <= 8'b0;
regfile[49] <= 8'b0;
regfile[50] <= 8'b0;
regfile[51] <= 8'b0;
regfile[52] <= 8'b0;
regfile[53] <= 8'b0;
regfile[54] <= 8'b0;
regfile[55] <= 8'b0;
regfile[56] <= 8'b0;
regfile[57] <= 8'b0;
regfile[58] <= 8'b0;
regfile[59] <= 8'b0;
regfile[60] <= 8'b0;
regfile[61] <= 8'b0;
regfile[62] <= 8'b0;
regfile[63] <= 8'b0;
regfile[64] <= 8'b0;
regfile[65] <= 8'b0;
regfile[66] <= 8'b0;
regfile[67] <= 8'b0;
regfile[68] <= 8'b0;
regfile[69] <= 8'b0;
regfile[70] <= 8'b0;
regfile[71] <= 8'b0;
regfile[72] <= 8'b0;
regfile[73] <= 8'b0;
regfile[74] <= 8'b0;
regfile[75] <= 8'b0;
regfile[76] <= 8'b0;
regfile[77] <= 8'b0;
regfile[78] <= 8'b0;
regfile[79] <= 8'b0;
regfile[80] <= 8'b0;
regfile[81] <= 8'b0;
regfile[82] <= 8'b0;
regfile[83] <= 8'b0;
regfile[84] <= 8'b0;
regfile[85] <= 8'b0;
regfile[86] <= 8'b0;
regfile[87] <= 8'b0;
regfile[88] <= 8'b0;
regfile[89] <= 8'b0;
regfile[90] <= 8'b0;
regfile[91] <= 8'b0;
regfile[92] <= 8'b0;
regfile[93] <= 8'b0;
regfile[94] <= 8'b0;
regfile[95] <= 8'b0;
regfile[96] <= 8'b0;
regfile[97] <= 8'b0;
regfile[98] <= 8'b0;
regfile[99] <= 8'b0;
regfile[100] <= 8'b0;
regfile[101] <= 8'b0;
regfile[102] <= 8'b0;
regfile[103] <= 8'b0;
regfile[104] <= 8'b0;
regfile[105] <= 8'b0;
regfile[106] <= 8'b0;
regfile[107] <= 8'b0;
regfile[108] <= 8'b0;
regfile[109] <= 8'b0;
regfile[110] <= 8'b0;
regfile[111] <= 8'b0;
regfile[112] <= 8'b0;
regfile[113] <= 8'b0;
regfile[114] <= 8'b0;
regfile[115] <= 8'b0;
regfile[116] <= 8'b0;
regfile[117] <= 8'b0;
regfile[118] <= 8'b0;
regfile[119] <= 8'b0;
regfile[120] <= 8'b0;
regfile[121] <= 8'b0;
regfile[122] <= 8'b0;
regfile[123] <= 8'b0;
regfile[124] <= 8'b0;
regfile[125] <= 8'b0;
regfile[126] <= 8'b0;
regfile[127] <= 8'b0;
      
   end
   else
   if (write_valid_f)
   begin
      
      regfile[write_index_f] <= (write_data_f & write_mask_f) | (regfile[write_index_f] & ~write_mask_f);
   end
end
endmodule
module rf_l15_wmt(
   input wire clk,
   input wire rst_n,
   input wire read_valid,
   input wire [6:0] read_index,
   input wire write_valid,
   input wire [6:0] write_index,
   input wire [4*((2+0)+1)-1:0] write_mask,
   input wire [4*((2+0)+1)-1:0] write_data,
   output wire [4*((2+0)+1)-1:0] read_data
   );
reg [4*((2+0)+1)-1:0] data_out_f;
reg [6:0] write_index_f;
reg [4*((2+0)+1)-1:0] write_data_f;
reg [4*((2+0)+1)-1:0] write_mask_f;
reg write_valid_f;
reg [4*((2+0)+1)-1:0] regfile [0:(512/4)-1];
always @ (posedge clk)
begin
   if (read_valid)
      data_out_f <= regfile[read_index];
end
assign read_data = data_out_f;
always @ (posedge clk)
begin
   write_valid_f <= write_valid;
   if (write_valid)
   begin
      write_data_f <= write_data;
      write_index_f <= write_index;
      write_mask_f <= write_mask;
   end
end
always @ (posedge clk)
begin
   if (!rst_n)
   begin
      regfile[0][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[0][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[0][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[0][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[1][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[1][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[1][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[1][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[2][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[2][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[2][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[2][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[3][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[3][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[3][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[3][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[4][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[4][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[4][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[4][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[5][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[5][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[5][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[5][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[6][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[6][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[6][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[6][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[7][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[7][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[7][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[7][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[8][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[8][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[8][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[8][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[9][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[9][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[9][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[9][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[10][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[10][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[10][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[10][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[11][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[11][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[11][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[11][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[12][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[12][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[12][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[12][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[13][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[13][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[13][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[13][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[14][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[14][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[14][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[14][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[15][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[15][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[15][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[15][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[16][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[16][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[16][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[16][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[17][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[17][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[17][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[17][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[18][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[18][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[18][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[18][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[19][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[19][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[19][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[19][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[20][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[20][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[20][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[20][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[21][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[21][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[21][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[21][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[22][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[22][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[22][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[22][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[23][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[23][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[23][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[23][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[24][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[24][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[24][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[24][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[25][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[25][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[25][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[25][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[26][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[26][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[26][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[26][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[27][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[27][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[27][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[27][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[28][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[28][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[28][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[28][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[29][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[29][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[29][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[29][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[30][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[30][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[30][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[30][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[31][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[31][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[31][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[31][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[32][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[32][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[32][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[32][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[33][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[33][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[33][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[33][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[34][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[34][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[34][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[34][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[35][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[35][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[35][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[35][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[36][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[36][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[36][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[36][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[37][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[37][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[37][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[37][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[38][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[38][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[38][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[38][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[39][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[39][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[39][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[39][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[40][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[40][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[40][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[40][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[41][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[41][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[41][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[41][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[42][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[42][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[42][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[42][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[43][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[43][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[43][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[43][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[44][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[44][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[44][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[44][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[45][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[45][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[45][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[45][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[46][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[46][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[46][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[46][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[47][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[47][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[47][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[47][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[48][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[48][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[48][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[48][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[49][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[49][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[49][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[49][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[50][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[50][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[50][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[50][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[51][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[51][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[51][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[51][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[52][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[52][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[52][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[52][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[53][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[53][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[53][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[53][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[54][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[54][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[54][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[54][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[55][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[55][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[55][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[55][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[56][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[56][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[56][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[56][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[57][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[57][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[57][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[57][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[58][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[58][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[58][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[58][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[59][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[59][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[59][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[59][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[60][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[60][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[60][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[60][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[61][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[61][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[61][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[61][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[62][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[62][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[62][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[62][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[63][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[63][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[63][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[63][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[64][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[64][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[64][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[64][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[65][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[65][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[65][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[65][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[66][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[66][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[66][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[66][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[67][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[67][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[67][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[67][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[68][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[68][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[68][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[68][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[69][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[69][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[69][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[69][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[70][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[70][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[70][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[70][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[71][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[71][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[71][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[71][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[72][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[72][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[72][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[72][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[73][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[73][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[73][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[73][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[74][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[74][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[74][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[74][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[75][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[75][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[75][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[75][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[76][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[76][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[76][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[76][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[77][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[77][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[77][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[77][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[78][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[78][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[78][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[78][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[79][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[79][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[79][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[79][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[80][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[80][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[80][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[80][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[81][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[81][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[81][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[81][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[82][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[82][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[82][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[82][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[83][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[83][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[83][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[83][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[84][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[84][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[84][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[84][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[85][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[85][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[85][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[85][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[86][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[86][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[86][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[86][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[87][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[87][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[87][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[87][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[88][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[88][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[88][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[88][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[89][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[89][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[89][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[89][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[90][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[90][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[90][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[90][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[91][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[91][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[91][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[91][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[92][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[92][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[92][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[92][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[93][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[93][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[93][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[93][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[94][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[94][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[94][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[94][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[95][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[95][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[95][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[95][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[96][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[96][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[96][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[96][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[97][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[97][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[97][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[97][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[98][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[98][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[98][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[98][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[99][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[99][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[99][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[99][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[100][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[100][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[100][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[100][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[101][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[101][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[101][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[101][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[102][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[102][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[102][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[102][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[103][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[103][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[103][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[103][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[104][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[104][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[104][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[104][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[105][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[105][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[105][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[105][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[106][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[106][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[106][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[106][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[107][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[107][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[107][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[107][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[108][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[108][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[108][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[108][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[109][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[109][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[109][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[109][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[110][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[110][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[110][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[110][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[111][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[111][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[111][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[111][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[112][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[112][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[112][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[112][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[113][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[113][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[113][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[113][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[114][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[114][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[114][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[114][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[115][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[115][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[115][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[115][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[116][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[116][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[116][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[116][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[117][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[117][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[117][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[117][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[118][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[118][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[118][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[118][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[119][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[119][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[119][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[119][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[120][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[120][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[120][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[120][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[121][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[121][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[121][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[121][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[122][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[122][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[122][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[122][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[123][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[123][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[123][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[123][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[124][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[124][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[124][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[124][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[125][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[125][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[125][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[125][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[126][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[126][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[126][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[126][(3+1)*((2+0)+1)-1] <= 1'b0;
regfile[127][(0+1)*((2+0)+1)-1] <= 1'b0;
regfile[127][(1+1)*((2+0)+1)-1] <= 1'b0;
regfile[127][(2+1)*((2+0)+1)-1] <= 1'b0;
regfile[127][(3+1)*((2+0)+1)-1] <= 1'b0;
   end
   else
   if (write_valid_f)
   begin
      
      regfile[write_index_f] <= (write_data_f & write_mask_f) | (regfile[write_index_f] & ~write_mask_f);
   end
end
endmodule
      
 
module l2(
    input wire clk,
    input wire rst_n,
    input wire [14-1:0] chipid,
    input wire [8-1:0] coreid_x,
    input wire [8-1:0] coreid_y,
    input wire noc1_valid_in,
    input wire [64-1:0] noc1_data_in,
    output wire noc1_ready_in,
    input wire noc3_valid_in,
    input wire [64-1:0] noc3_data_in,
    output wire noc3_ready_in,
    output wire noc2_valid_out,
    output wire [64-1:0] noc2_data_out,
    input wire noc2_ready_out,
    
    output wire [4-1:0] srams_rtap_data,
    input wire  [4-1:0] rtap_srams_bist_command,
    input wire  [4-1:0] rtap_srams_bist_data
);
wire [4-1:0] data_rtap_data;
wire [4-1:0] dir_rtap_data;
wire [4-1:0] tag_rtap_data;
wire [4-1:0] state_rtap_data;
assign srams_rtap_data = data_rtap_data
                            | dir_rtap_data
                            | tag_rtap_data
                            | state_rtap_data;
localparam y = 1'b1;
localparam n = 1'b0;
wire mshr_cam_en_p1;
wire mshr_wr_state_en_p1;
wire mshr_wr_data_en_p1;
wire mshr_pending_ready_p1;
wire [2-1:0] mshr_state_in_p1;
wire [120+2-1:0] mshr_data_in_p1;
wire [120+2-1:0] mshr_data_mask_in_p1;
wire [3-1:0] mshr_inv_counter_rd_index_in_p1;
wire [3-1:0] mshr_wr_index_in_p1;
wire [8-1:0] mshr_addr_in_p1;
wire mshr_rd_en_p2;
wire mshr_wr_state_en_p2;
wire mshr_wr_data_en_p2;
wire mshr_inc_counter_en_p2;
wire [2-1:0] mshr_state_in_p2;
wire [120+2-1:0] mshr_data_in_p2;
wire [120+2-1:0] mshr_data_mask_in_p2;
wire [3-1:0] mshr_rd_index_in_p2;
wire [3-1:0] mshr_wr_index_in_p2;
wire mshr_hit;
wire [3-1:0] mshr_hit_index;
wire [2-1:0] rd_mshr_state_out;
wire [120+2-1:0] rd_mshr_data_out;
wire [120+2-1:0] cam_mshr_data_out;
wire [120+2-1:0] pending_mshr_data_out;
wire [6-1:0] mshr_inv_counter_out;
wire [3:0] mshr_empty_slots;
wire mshr_pending;
wire [3-1:0] mshr_pending_index;
wire [3-1:0] mshr_empty_index;
wire state_rd_en_p1;
wire state_wr_en_p1;
wire [8-1:0] state_rd_addr_p1;
wire [8-1:0] state_wr_addr_p1;
wire [15*4+2+4-1:0] state_data_in_p1;
wire [15*4+2+4-1:0] state_data_mask_in_p1;
wire state_rd_en_p2;
wire state_wr_en_p2;
wire [8-1:0] state_rd_addr_p2;
wire [8-1:0] state_wr_addr_p2;
wire [15*4+2+4-1:0] state_data_in_p2;
wire [15*4+2+4-1:0] state_data_mask_in_p2;
wire [15*4+2+4-1:0] state_data_out;
wire tag_clk_en_p1;
wire tag_rdw_en_p1;
wire [8-1:0] tag_addr_p1;
wire [104-1:0] tag_data_in_p1;
wire [104-1:0] tag_data_mask_in_p1;
wire tag_clk_en_p2;
wire tag_rdw_en_p2;
wire [8-1:0] tag_addr_p2;
wire [104-1:0] tag_data_in_p2;
wire [104-1:0] tag_data_mask_in_p2;
wire [104-1:0] tag_data_out;
wire dir_clk_en_p1;
wire dir_rdw_en_p1;
wire [8+2-1:0] dir_addr_p1;
wire [64-1:0] dir_data_in_p1;
wire [64-1:0] dir_data_mask_in_p1;
wire dir_clk_en_p2;
wire dir_rdw_en_p2;
wire [8+2-1:0] dir_addr_p2;
wire [64-1:0] dir_data_in_p2;
wire [64-1:0] dir_data_mask_in_p2;
wire [64-1:0] dir_data_out;
wire data_clk_en_p1;
wire data_rdw_en_p1;
wire [8+2+2-1:0] data_addr_p1;
wire [144-1:0] data_data_in_p1;
wire [144-1:0] data_data_mask_in_p1;
wire data_clk_en_p2;
wire data_rdw_en_p2;
wire [8+2+2-1:0] data_addr_p2;
wire [144-1:0] data_data_in_p2;
wire [144-1:0] data_data_mask_in_p2;
wire [144-1:0] data_data_out;
wire smc_rd_en;
wire smc_rd_diag_en;
wire smc_wr_diag_en;
wire smc_flush_en;
wire [2-1:0] smc_addr_op;
wire [16-1:0] smc_rd_addr_in;
wire smc_wr_en_p1;
wire [16-1:0] smc_wr_addr_in_p1;
wire [128-1:0] smc_data_in_p1;
wire smc_wr_en_p2;
wire [16-1:0] smc_wr_addr_in_p2;
wire [128-1:0] smc_data_in_p2;
wire [2-1:0] broadcast_counter_op_p1;
wire broadcast_counter_op_val_p1;
wire [2-1:0] broadcast_counter_op_p2;
wire broadcast_counter_op_val_p2;
wire smc_hit;
wire [30-1:0] smc_data_out;
wire [4-1:0] smc_valid_out;
wire [14-1:0] smc_tag_out;
wire broadcast_counter_zero1;
wire broadcast_counter_max1;
wire broadcast_counter_avail1;
wire [14-1:0] broadcast_chipid_out1;
wire [8-1:0] broadcast_x_out1;
wire [8-1:0] broadcast_y_out1;
wire broadcast_counter_zero2;
wire broadcast_counter_max2;
wire broadcast_counter_avail2;
wire [14-1:0] broadcast_chipid_out2;
wire [8-1:0] broadcast_x_out2;
wire [8-1:0] broadcast_y_out2;
wire reg_rd_en;
wire reg_wr_en;
wire [8-1:0] reg_rd_addr_type;
wire [8-1:0] reg_wr_addr_type;
wire [64-1:0] reg_data_out;
wire [64-1:0] reg_data_in;
wire l2_access_valid;
wire l2_miss_valid;
wire data_ecc_corr_error;
wire data_ecc_uncorr_error;
wire [8+2+2-1:0] data_ecc_addr;
wire [40-1:0] error_addr;
wire [34-1:0] my_nodeid;
wire [14+8+8-1:0] core_max;
wire csm_en;
wire [22-1:0] smt_base_addr;
wire pipe2_valid_S1;
wire pipe2_valid_S2;
wire pipe2_valid_S3;
wire [8-1:0] pipe2_msg_type_S1;
wire [8-1:0] pipe2_msg_type_S2;
wire [8-1:0] pipe2_msg_type_S3;
wire [40-1:0] pipe2_addr_S1;
wire [40-1:0] pipe2_addr_S2;
wire [40-1:0] pipe2_addr_S3;
wire active_S1;
wire active_S2;
wire active_S3;
l2_config_regs config_regs(
    .clk                    (clk),
    .rst_n                  (rst_n),
    .chipid                 (chipid),
    .coreid_x               (coreid_x),
    .coreid_y               (coreid_y),
    .l2_access_valid        (l2_access_valid),
    .l2_miss_valid          (l2_miss_valid),
    .data_ecc_corr_error    (data_ecc_corr_error),
    .data_ecc_uncorr_error  (data_ecc_uncorr_error),
    .data_ecc_addr          (data_ecc_addr),
    .error_addr             (error_addr),
    .reg_rd_en              (reg_rd_en),
    .reg_wr_en              (reg_wr_en),
    .reg_rd_addr_type       (reg_rd_addr_type),
    .reg_wr_addr_type       (reg_wr_addr_type),
    .reg_data_in            (reg_data_in),
    .reg_data_out           (reg_data_out),
    .my_nodeid              (my_nodeid),
    .core_max               (core_max),
    
    .csm_en                 (csm_en),
    
    
    .smt_base_addr          (smt_base_addr)
);
l2_mshr_wrap mshr_wrap(
    .clk                    (clk),
    .rst_n                  (rst_n),
    .pipe_wr_sel            (active_S3),
    .cam_en1                (mshr_cam_en_p1),
    .wr_state_en1           (mshr_wr_state_en_p1),
    .wr_data_en1            (mshr_wr_data_en_p1),
    .pending_ready1         (mshr_pending_ready_p1),
    .state_in1              (mshr_state_in_p1),
    .data_in1               (mshr_data_in_p1),
    .data_mask_in1          (mshr_data_mask_in_p1),
    .inv_counter_rd_index_in1(mshr_inv_counter_rd_index_in_p1),
    .wr_index_in1           (mshr_wr_index_in_p1),
    .addr_in1               (mshr_addr_in_p1),
    .wr_state_en2           (mshr_wr_state_en_p2),
    .wr_data_en2            (mshr_wr_data_en_p2),
 
    .inc_counter_en2        (mshr_inc_counter_en_p2),
    .state_in2              (mshr_state_in_p2),
    .data_in2               (mshr_data_in_p2),
    .data_mask_in2          (mshr_data_mask_in_p2),
    .rd_index_in2           (mshr_rd_index_in_p2),
    .wr_index_in2           (mshr_wr_index_in_p2),
    .hit                    (mshr_hit),
    .hit_index              (mshr_hit_index),
    .rd_state_out           (rd_mshr_state_out),
    .rd_data_out            (rd_mshr_data_out),
    
    .cam_data_out           (cam_mshr_data_out),
    .pending_data_out       (pending_mshr_data_out),
    .inv_counter_out        (mshr_inv_counter_out), 
    .empty_slots            (mshr_empty_slots),
    .pending                (mshr_pending),
    .pending_index          (mshr_pending_index),
    .empty_index            (mshr_empty_index)
);
l2_state_wrap state_wrap(
    .clk                    (clk),
    .rst_n                  (rst_n),
    .pdout_en               (1'b0),
    .deepsleep              (1'b0),
    .pipe_rd_sel            (active_S1),
    .pipe_wr_sel            (active_S3),
    .rd_en1                 (state_rd_en_p1),
    .wr_en1                 (state_wr_en_p1),
    .rd_addr1               (state_rd_addr_p1),
    .wr_addr1               (state_wr_addr_p1),
    .data_in1               (state_data_in_p1),
    .data_mask_in1          (state_data_mask_in_p1),
    .rd_en2                 (state_rd_en_p2),
    .wr_en2                 (state_wr_en_p2),
    .rd_addr2               (state_rd_addr_p2),
    .wr_addr2               (state_wr_addr_p2),
    .data_in2               (state_data_in_p2),
    .data_mask_in2          (state_data_mask_in_p2),
    .data_out               (state_data_out),
    .pdata_out              (),
    
    .srams_rtap_data (state_rtap_data),
    .rtap_srams_bist_command (rtap_srams_bist_command),
    .rtap_srams_bist_data (rtap_srams_bist_data)
);
l2_tag_wrap tag_wrap(
    .clk                    (clk),
    .rst_n                  (rst_n),
    .pdout_en               (1'b0),
    .deepsleep              (1'b0),
    .pipe_sel               (active_S1),
    .clk_en1                (tag_clk_en_p1),
    .rdw_en1                (tag_rdw_en_p1),
    .addr1                  (tag_addr_p1),
    .data_in1               (tag_data_in_p1),
    .data_mask_in1          (tag_data_mask_in_p1),
    .clk_en2                (tag_clk_en_p2),
    .rdw_en2                (tag_rdw_en_p2),
    .addr2                  (tag_addr_p2),
    .data_in2               (tag_data_in_p2),
    .data_mask_in2          (tag_data_mask_in_p2),
    .data_out               (tag_data_out),
    .pdata_out              (),
    
    .srams_rtap_data (tag_rtap_data),
    .rtap_srams_bist_command (rtap_srams_bist_command),
    .rtap_srams_bist_data (rtap_srams_bist_data)
);
l2_dir_wrap dir_wrap(
    .clk                    (clk),
    .rst_n                  (rst_n),
    .pdout_en               (1'b0),
    .deepsleep              (1'b0),
    .pipe_sel               (active_S2),
    .clk_en1                (dir_clk_en_p1),
    .rdw_en1                (dir_rdw_en_p1),
    .addr1                  (dir_addr_p1),
    .data_in1               (dir_data_in_p1),
    .data_mask_in1          (dir_data_mask_in_p1),
    .clk_en2                (dir_clk_en_p2),
    .rdw_en2                (dir_rdw_en_p2),
    .addr2                  (dir_addr_p2),
    .data_in2               (dir_data_in_p2),
    .data_mask_in2          (dir_data_mask_in_p2),
    .data_out               (dir_data_out),
    .pdata_out              (),
    
    .srams_rtap_data (dir_rtap_data),
    .rtap_srams_bist_command (rtap_srams_bist_command),
    .rtap_srams_bist_data (rtap_srams_bist_data)
);
l2_data_wrap data_wrap(
    .clk                    (clk),
    .rst_n                  (rst_n),
    .pdout_en               (1'b0),
    .deepsleep              (1'b0),
    .pipe_sel               (active_S2),
    .clk_en1                (data_clk_en_p1),
    .rdw_en1                (data_rdw_en_p1),
    .addr1                  (data_addr_p1),
    .data_in1               (data_data_in_p1),
    .data_mask_in1          (data_data_mask_in_p1),
    .clk_en2                (data_clk_en_p2),
    .rdw_en2                (data_rdw_en_p2),
    .addr2                  (data_addr_p2),
    .data_in2               (data_data_in_p2),
    .data_mask_in2          (data_data_mask_in_p2),
    .data_out               (data_data_out),
    .pdata_out              (),
    
    .srams_rtap_data (data_rtap_data),
    .rtap_srams_bist_command (rtap_srams_bist_command),
    .rtap_srams_bist_data (rtap_srams_bist_data)
);
l2_smc_wrap smc_wrap(
    .clk                    (clk),
    .rst_n                  (rst_n),
    .pipe_sel               (active_S2),
    .rd_en                  (smc_rd_en),
    .rd_diag_en             (smc_rd_diag_en),
    .flush_en               (smc_flush_en),
    .addr_op                (smc_addr_op),
    .rd_addr_in             (smc_rd_addr_in),
    .wr_en1                 (smc_wr_en_p1),
    .wr_addr_in1            (smc_wr_addr_in_p1),
    .data_in1               (smc_data_in_p1),
    .wr_diag_en1            (smc_wr_diag_en),
    .wr_en2                 (smc_wr_en_p2),
    .wr_addr_in2            (smc_wr_addr_in_p2),
    .data_in2               (smc_data_in_p2),
    .wr_diag_en2            (1'b0),
    .hit                    (smc_hit),
    .data_out               (smc_data_out),
    .valid_out              (smc_valid_out),
    .tag_out                (smc_tag_out)
);
l2_broadcast_counter_wrap l2_broadcast_counter_wrap(
    .clk                    (clk),
    .rst_n                  (rst_n),
    .chipid_max             (core_max[29:16]),
    .x_max                  (core_max[7:0]),
    .y_max                  (core_max[15:8]),
    .pipe_sel               (active_S2),
    .counter_op1            (broadcast_counter_op_p1),
    .counter_op_val1        (broadcast_counter_op_val_p1),
    .counter_op2            (broadcast_counter_op_p2),
    .counter_op_val2        (broadcast_counter_op_val_p2),
    .zero1                  (broadcast_counter_zero1),
    .max1                   (broadcast_counter_max1),
    .avail1                 (broadcast_counter_avail1),
    .chipid_out1            (broadcast_chipid_out1),
    .x_out1                 (broadcast_x_out1),
    .y_out1                 (broadcast_y_out1),
    .zero2                  (broadcast_counter_zero2),
    .max2                   (broadcast_counter_max2),
    .avail2                 (broadcast_counter_avail2),
    .chipid_out2            (broadcast_chipid_out2),
    .x_out2                 (broadcast_x_out2),
    .y_out2                 (broadcast_y_out2)
);
l2_pipe1 pipe1(
    .clk                    (clk),
    .rst_n                  (rst_n),
    .my_nodeid              (my_nodeid),
    
    .csm_en                 (csm_en),
    
    .smt_base_addr          (smt_base_addr),
    .noc_valid_in           (noc1_valid_in),
    .noc_data_in            (noc1_data_in),
    .noc_ready_in           (noc1_ready_in),
    .noc_valid_out          (noc2_valid_out),
    .noc_data_out           (noc2_data_out),
    .noc_ready_out          (noc2_ready_out),
    .pipe2_valid_S1         (pipe2_valid_S1),
    .pipe2_valid_S2         (pipe2_valid_S2),
    .pipe2_valid_S3         (pipe2_valid_S3),
    .pipe2_msg_type_S1      (pipe2_msg_type_S1),
    .pipe2_msg_type_S2      (pipe2_msg_type_S2),
    .pipe2_msg_type_S3      (pipe2_msg_type_S3),
    .pipe2_addr_S1          (pipe2_addr_S1),
    .pipe2_addr_S2          (pipe2_addr_S2),
    .pipe2_addr_S3          (pipe2_addr_S3),
    .global_stall_S1        (active_S1),
    .global_stall_S2        (active_S2),
    .global_stall_S4        (active_S3),
    .mshr_hit               (mshr_hit),
    .cam_mshr_data_out      (cam_mshr_data_out),
    .pending_mshr_data_out  (pending_mshr_data_out),
    .mshr_inv_counter_out   (mshr_inv_counter_out),
    .mshr_empty_slots       (mshr_empty_slots),
    .mshr_pending           (mshr_pending),
    .mshr_pending_index     (mshr_pending_index),
    .mshr_empty_index       (mshr_empty_index),
    
    .broadcast_counter_zero (broadcast_counter_zero1),
    .broadcast_counter_max  (broadcast_counter_max1),
    .broadcast_counter_avail(broadcast_counter_avail1),
    .broadcast_chipid_out   (broadcast_chipid_out1),
    .broadcast_x_out        (broadcast_x_out1),
    .broadcast_y_out        (broadcast_y_out1),
    
    .state_data_out         (state_data_out),
    .tag_data_out           (tag_data_out),
    .dir_data_out           (dir_data_out),
    .data_data_out          (data_data_out),
    .l2_access_valid        (l2_access_valid),
    .l2_miss_valid          (l2_miss_valid),
    .data_ecc_corr_error    (data_ecc_corr_error),
    .data_ecc_uncorr_error  (data_ecc_uncorr_error),
    .data_ecc_addr          (data_ecc_addr),
    .error_addr             (error_addr),
    .reg_rd_en              (reg_rd_en),
    .reg_wr_en              (reg_wr_en),
    .reg_rd_addr_type       (reg_rd_addr_type),
    .reg_wr_addr_type       (reg_wr_addr_type),
    .reg_data_out           (reg_data_out),
    .reg_data_in            (reg_data_in),
    .mshr_cam_en            (mshr_cam_en_p1),
    .mshr_wr_state_en       (mshr_wr_state_en_p1),
    .mshr_wr_data_en        (mshr_wr_data_en_p1),
    .mshr_pending_ready     (mshr_pending_ready_p1),
    .mshr_state_in          (mshr_state_in_p1),
    .mshr_data_in           (mshr_data_in_p1),
    .mshr_data_mask_in      (mshr_data_mask_in_p1),
    .mshr_inv_counter_rd_index_in(mshr_inv_counter_rd_index_in_p1),
    .mshr_wr_index_in       (mshr_wr_index_in_p1),
    .mshr_addr_in           (mshr_addr_in_p1),
    .state_rd_en            (state_rd_en_p1),
    .state_wr_en            (state_wr_en_p1),
    .state_rd_addr          (state_rd_addr_p1),
    .state_wr_addr          (state_wr_addr_p1),
    .state_data_in          (state_data_in_p1),
    .state_data_mask_in     (state_data_mask_in_p1),
    .tag_clk_en             (tag_clk_en_p1),
    .tag_rdw_en             (tag_rdw_en_p1),
    .tag_addr               (tag_addr_p1),
    .tag_data_in            (tag_data_in_p1),
    .tag_data_mask_in       (tag_data_mask_in_p1),
    .dir_clk_en             (dir_clk_en_p1),
    .dir_rdw_en             (dir_rdw_en_p1),
    .dir_addr               (dir_addr_p1),
    .dir_data_in            (dir_data_in_p1),
    .dir_data_mask_in       (dir_data_mask_in_p1),
    
    .broadcast_counter_op   (broadcast_counter_op_p1),
    .broadcast_counter_op_val(broadcast_counter_op_val_p1),
    .smc_rd_en              (smc_rd_en),
    .smc_rd_addr_in         (smc_rd_addr_in),
    .smc_rd_diag_en         (smc_rd_diag_en),
    .smc_flush_en           (smc_flush_en),
    .smc_addr_op            (smc_addr_op),
    .smc_wr_diag_en         (smc_wr_diag_en),
    .smc_wr_en              (smc_wr_en_p1),
    .smc_wr_addr_in         (smc_wr_addr_in_p1),
    .smc_data_in            (smc_data_in_p1),
    .smc_hit                (smc_hit),
    .smc_data_out           (smc_data_out),
    .smc_valid_out          (smc_valid_out),
    .smc_tag_out            (smc_tag_out),
    
    .data_clk_en            (data_clk_en_p1),
    .data_rdw_en            (data_rdw_en_p1),
    .data_addr              (data_addr_p1),
    .data_data_in           (data_data_in_p1),
    .data_data_mask_in      (data_data_mask_in_p1)
);
l2_pipe2 pipe2(
    .clk                    (clk),
    .rst_n                  (rst_n),
    
    .csm_en                 (csm_en),
    
    .noc_valid_in           (noc3_valid_in),
    .noc_data_in            (noc3_data_in),
    .noc_ready_in           (noc3_ready_in),
    .mshr_state_out         (rd_mshr_state_out),
    .mshr_data_out          (rd_mshr_data_out),
    
    .broadcast_counter_zero (broadcast_counter_zero2),
    .broadcast_counter_max  (broadcast_counter_max2),
    .broadcast_chipid_out   (broadcast_chipid_out2),
    .broadcast_x_out        (broadcast_x_out2),
    .broadcast_y_out        (broadcast_y_out2),
    
    .state_data_out         (state_data_out),
    .tag_data_out           (tag_data_out),
    .dir_data_out           (dir_data_out),
    .mshr_rd_en             (mshr_rd_en_p2),
    .mshr_wr_state_en       (mshr_wr_state_en_p2),
    .mshr_wr_data_en        (mshr_wr_data_en_p2),
    .mshr_inc_counter_en    (mshr_inc_counter_en_p2),
    .mshr_state_in          (mshr_state_in_p2),
    .mshr_data_in           (mshr_data_in_p2),
    .mshr_data_mask_in      (mshr_data_mask_in_p2),
    .mshr_rd_index_in       (mshr_rd_index_in_p2),
    .mshr_wr_index_in       (mshr_wr_index_in_p2),
    .state_rd_en            (state_rd_en_p2),
    .state_wr_en            (state_wr_en_p2),
    .state_rd_addr          (state_rd_addr_p2),
    .state_wr_addr          (state_wr_addr_p2),
    .state_data_in          (state_data_in_p2),
    .state_data_mask_in     (state_data_mask_in_p2),
    .tag_clk_en             (tag_clk_en_p2),
    .tag_rdw_en             (tag_rdw_en_p2),
    .tag_addr               (tag_addr_p2),
    .tag_data_in            (tag_data_in_p2),
    .tag_data_mask_in       (tag_data_mask_in_p2),
    .dir_clk_en             (dir_clk_en_p2),
    .dir_rdw_en             (dir_rdw_en_p2),
    .dir_addr               (dir_addr_p2),
    .dir_data_in            (dir_data_in_p2),
    .dir_data_mask_in       (dir_data_mask_in_p2),
    .data_clk_en            (data_clk_en_p2),
    .data_rdw_en            (data_rdw_en_p2),
    .data_addr              (data_addr_p2),
    .data_data_in           (data_data_in_p2),
    .data_data_mask_in      (data_data_mask_in_p2),
    
    .broadcast_counter_op   (broadcast_counter_op_p2),
    .broadcast_counter_op_val(broadcast_counter_op_val_p2),
    .smc_wr_en              (smc_wr_en_p2),
    .smc_wr_addr_in         (smc_wr_addr_in_p2),
    .smc_data_in            (smc_data_in_p2),
    
    .valid_S1               (pipe2_valid_S1),
    .valid_S2               (pipe2_valid_S2),
    .valid_S3               (pipe2_valid_S3),
    .msg_type_S1            (pipe2_msg_type_S1),
    .msg_type_S2            (pipe2_msg_type_S2),
    .msg_type_S3            (pipe2_msg_type_S3),
    .addr_S1                (pipe2_addr_S1),
    .addr_S2                (pipe2_addr_S2),
    .addr_S3                (pipe2_addr_S3),
    .active_S1              (active_S1),
    .active_S2              (active_S2),
    .active_S3              (active_S3)
);
endmodule
      
 
module l2_amo_alu #(
  parameter SWAP_ENDIANESS = 1
) (
  input      [4-1:0] amo_alu_op,
  input      [40-1:0]      address,
  input      [3-1:0] data_size,
  input      [128-1:0]  memory_operand,
  input      [128-1:0]  cpu_operand,
  output reg [128-1:0]  amo_result
);
wire [63:0] amo_operand_a_mux, amo_operand_b_mux;
wire [63:0] amo_operand_a_swp, amo_operand_b_swp;
reg  [63:0] amo_operand_a, amo_operand_b;
reg  [63:0] amo_64b_tmp, amo_64b_result;
reg  [64:0] adder_operand_a, adder_operand_b;
wire [64:0] adder_sum;
wire [7-7:0] dword_offset;
assign dword_offset      = address[7-4:3];
assign amo_operand_a_mux = memory_operand[dword_offset*64 +: 64];
assign amo_operand_b_mux = cpu_operand[dword_offset*64 +: 64];
generate
  if (SWAP_ENDIANESS) begin : g_swap_in
    assign amo_operand_a_swp = {amo_operand_a_mux[ 0 +:8],
                                amo_operand_a_mux[ 8 +:8],
                                amo_operand_a_mux[16 +:8],
                                amo_operand_a_mux[24 +:8],
                                amo_operand_a_mux[32 +:8],
                                amo_operand_a_mux[40 +:8],
                                amo_operand_a_mux[48 +:8],
                                amo_operand_a_mux[56 +:8]};
    assign amo_operand_b_swp = {amo_operand_b_mux[ 0 +:8],
                                amo_operand_b_mux[ 8 +:8],
                                amo_operand_b_mux[16 +:8],
                                amo_operand_b_mux[24 +:8],
                                amo_operand_b_mux[32 +:8],
                                amo_operand_b_mux[40 +:8],
                                amo_operand_b_mux[48 +:8],
                                amo_operand_b_mux[56 +:8]};
  end else begin : g_swap_in
    assign amo_operand_a_swp = amo_operand_a_mux;
    assign amo_operand_b_swp = amo_operand_b_mux;
  end
endgenerate
always @* begin
  amo_operand_a = 64'h0;
  amo_operand_b = 64'h0;
  case (data_size)
    3'b001: begin
      amo_operand_a[56 +: 8]     = amo_operand_a_swp[address[2:0]*8 +: 8];
      amo_operand_b[56 +: 8]     = amo_operand_b_swp[address[2:0]*8 +: 8];
    end
    3'b010: begin
        amo_operand_a[48 +: 16]  = amo_operand_a_swp[address[2:1]*16 +: 16];
        amo_operand_b[48 +: 16]  = amo_operand_b_swp[address[2:1]*16 +: 16];
     end
    3'b011: begin
        amo_operand_a[32 +: 32]  = amo_operand_a_swp[address[2:2]*32 +: 32];
        amo_operand_b[32 +: 32]  = amo_operand_b_swp[address[2:2]*32 +: 32];
    end
    3'b100: begin
        amo_operand_a  = amo_operand_a_swp;
        amo_operand_b  = amo_operand_b_swp;
    end
    default: ;
  endcase 
end
assign adder_sum     = adder_operand_a + adder_operand_b;
always @*
begin
    adder_operand_a = $signed(amo_operand_a);
    adder_operand_b = $signed(amo_operand_b);
    amo_64b_tmp     = amo_operand_a;
    case (amo_alu_op)
        4'd0: ;
        4'd1: amo_64b_tmp = adder_sum[63:0];
        4'd2: amo_64b_tmp = amo_operand_a & amo_operand_b;
        4'd3:  amo_64b_tmp = amo_operand_a | amo_operand_b;
        4'd4: amo_64b_tmp = amo_operand_a ^ amo_operand_b;
        4'd5: begin
            adder_operand_b = -$signed(amo_operand_b);
            amo_64b_tmp = adder_sum[64] ? amo_operand_b : amo_operand_a;
        end
        4'd6: begin
            adder_operand_a = $unsigned(amo_operand_a);
            adder_operand_b = -$unsigned(amo_operand_b);
            amo_64b_tmp = adder_sum[64] ? amo_operand_b : amo_operand_a;
        end
        4'd7: begin
            adder_operand_b = -$signed(amo_operand_b);
            amo_64b_tmp = adder_sum[64] ? amo_operand_a : amo_operand_b;
        end
        4'd8: begin
            adder_operand_a = $unsigned(amo_operand_a);
            adder_operand_b = -$unsigned(amo_operand_b);
            amo_64b_tmp = adder_sum[64] ? amo_operand_a : amo_operand_b;
        end
        default: ;
    endcase
end
always @* begin
  
  amo_64b_result = amo_operand_a_swp;
  case (data_size)
    3'b001: begin
      amo_64b_result[address[2:0]*8 +: 8]     = amo_64b_tmp[56 +: 8];
    end
    3'b010: begin
        amo_64b_result[address[2:1]*16 +: 16]  = amo_64b_tmp[48 +: 16];
     end
    3'b011: begin
        amo_64b_result[address[2:2]*32 +: 32]  = amo_64b_tmp[32 +: 32];
    end
    3'b100: begin
        amo_64b_result  = amo_64b_tmp;
    end
    default: ;
  endcase 
  
  amo_result     = memory_operand;
  if (SWAP_ENDIANESS) begin
    amo_result[dword_offset*64 +: 64] = {amo_64b_result[ 0 +:8],
                                         amo_64b_result[ 8 +:8],
                                         amo_64b_result[16 +:8],
                                         amo_64b_result[24 +:8],
                                         amo_64b_result[32 +:8],
                                         amo_64b_result[40 +:8],
                                         amo_64b_result[48 +:8],
                                         amo_64b_result[56 +:8]};
  end else begin
    amo_result[dword_offset*64 +: 64] = amo_64b_result;
  end
end
endmodule
      
 
module l2_broadcast_counter(
    input wire clk,
    input wire rst_n,
    input wire [14-1:0] chipid_max,
    input wire [8-1:0] x_max,
    input wire [8-1:0] y_max,
    input wire [2-1:0] counter_op,
    input wire counter_op_val,
    
    output reg zero,
    output reg max,
    output reg [14-1:0] chipid_out,
    output reg [8-1:0] x_out,
    output reg [8-1:0] y_out
);
reg [14-1:0] chipid_f;
reg [14-1:0] chipid_next;
reg [8-1:0] x_f;
reg [8-1:0] x_next;
reg [8-1:0] y_f;
reg [8-1:0] y_next;
always @ *
begin
    if (!rst_n)
    begin
        chipid_next = 0;
        x_next = 0;
        y_next = 0;
    end
    else if (counter_op_val)
    begin
        if (counter_op == 2'd1)
        begin
            chipid_next = chipid_max;
            x_next = x_max;
            y_next = y_max;
        end
        else if (counter_op == 2'd0)
        begin
            chipid_next = 0;
            x_next = 0;
            y_next = 0;
        end
        else if (counter_op == 2'd2)
        begin
            if (x_f == x_max)
            begin
                if (y_f == y_max)
                begin
                    if(chipid_f == chipid_max)
                    begin
                        chipid_next = 0;
                        x_next = 0;
                        y_next = 0;
                    end
                    else        
                    begin
                        chipid_next = chipid_f + 1;
                        x_next = 0;
                        y_next = 0;
                    end
                end
                else
                begin
                    chipid_next = chipid_f;
                    x_next = 0;
                    y_next = y_f + 1;
                end
            end
            else
            begin
                chipid_next = chipid_f;
                x_next = x_f + 1;
                y_next = y_f;
            end
        end
        else
        begin
            chipid_next = chipid_f;
            x_next = x_f;
            y_next = y_f;
        end
    end
    else
    begin
        chipid_next = chipid_f;
        x_next = x_f;
        y_next = y_f;
    end
end
always @ (posedge clk)
begin
    chipid_f <= chipid_next;
    x_f <= x_next;
    y_f <= y_next;
end
always @ *
begin
    zero = (x_f == 0) && (y_f == 0) && (chipid_f == 0);
    max = (x_f == x_max) && (y_f == y_max) && (chipid_f == chipid_max);
end
always @ *
begin
    chipid_out = chipid_f;
    x_out = x_f;
    y_out = y_f;
end
endmodule
      
 
module l2_broadcast_counter_wrap(
    input wire clk,
    input wire rst_n,
    input wire [14-1:0] chipid_max,
    input wire [8-1:0] x_max,
    input wire [8-1:0] y_max,
    input wire pipe_sel,
    input wire [2-1:0] counter_op1,
    input wire counter_op_val1,
   
    input wire [2-1:0] counter_op2,
    input wire counter_op_val2,
 
    output wire zero1,
    output wire max1,
    output reg  avail1,
    output wire [14-1:0] chipid_out1,
    output wire [8-1:0] x_out1,
    output wire [8-1:0] y_out1,
    output wire zero2,
    output wire max2,
    output reg  avail2,
    output wire [14-1:0] chipid_out2,
    output wire [8-1:0] x_out2,
    output wire [8-1:0] y_out2
);
reg state_f;
reg state_next;
always @ *
begin
    if (!rst_n)
    begin
        state_next = 1'b0;
    end
    else
    begin
        if (counter_op_val1 && (counter_op1 == 2'd2))
        begin
            state_next = 1'b1;
        end
        else if (counter_op_val2 && (counter_op2 == 2'd0))
        begin
            state_next = 1'b0;
        end
        else
        begin
            state_next = state_f;
        end
    end
end
always @ (posedge clk)
begin
    state_f <= state_next;
end
always @ *
begin
    avail1 = (state_f == 1'b0);
    avail2 = (state_f == 1'b0);
end
l2_broadcast_counter l2_broadcast_counter1(
    .clk                (clk),
    .rst_n              (rst_n), 
    .chipid_max         (chipid_max),
    .x_max              (x_max),
    .y_max              (y_max),
    .counter_op         (counter_op1),
    .counter_op_val     (counter_op_val1),
    .zero               (zero1),
    .max                (max1),
    .chipid_out         (chipid_out1),
    .x_out              (x_out1),
    .y_out              (y_out1)
);
l2_broadcast_counter l2_broadcast_counter2(
    .clk                (clk),
    .rst_n              (rst_n), 
    .chipid_max         (chipid_max),
    .x_max              (x_max),
    .y_max              (y_max),
    .counter_op         (counter_op2),
    .counter_op_val     (counter_op_val2),
    .zero               (zero2),
    .max                (max2),
    .chipid_out         (chipid_out2),
    .x_out              (x_out2),
    .y_out              (y_out2)
);
endmodule
      
 
module l2_config_regs(
    input wire clk,
    input wire rst_n,
    input wire [14-1:0] chipid,
    input wire [8-1:0] coreid_x,
    input wire [8-1:0] coreid_y,
    input wire l2_access_valid,
    input wire l2_miss_valid,
    input wire data_ecc_corr_error,
    input wire data_ecc_uncorr_error,
    input wire [8+2+2-1:0] data_ecc_addr,
    input wire [40-1:0] error_addr,
    input wire reg_rd_en,
    input wire reg_wr_en,
    input wire [8-1:0] reg_rd_addr_type,
    input wire [8-1:0] reg_wr_addr_type,
    input wire [64-1:0] reg_data_in,
    output reg [64-1:0] reg_data_out,
    output reg [34-1:0] my_nodeid,
    output reg [14+8+8-1:0] core_max,
    output reg csm_en,
    output reg [22-1:0] smt_base_addr
);
reg [64-1:0] ctrl_reg_f;
reg [64-1:0] coreid_reg_f;
reg [64-1:0] l2_access_counter_reg_f;
reg [64-1:0] l2_miss_counter_reg_f;
reg [64-1:0] error_status_reg_f;
reg ctrl_reg_wr_en;
reg coreid_reg_wr_en;
reg l2_access_counter_reg_wr_en;
reg l2_miss_counter_reg_wr_en;
reg error_status_reg_wr_en;
reg error_status_en;
reg l2_access_counter_inc_en;
reg l2_miss_counter_inc_en;
always @ *
begin
    ctrl_reg_wr_en = reg_wr_en && (reg_wr_addr_type == 8'ha9); 
    coreid_reg_wr_en = reg_wr_en && (reg_wr_addr_type == 8'ha7); 
    l2_access_counter_reg_wr_en = reg_wr_en && (reg_wr_addr_type == 8'haa); 
    l2_miss_counter_reg_wr_en = reg_wr_en && (reg_wr_addr_type == 8'hab); 
    error_status_reg_wr_en = reg_wr_en && (reg_wr_addr_type == 8'ha8); 
    
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        ctrl_reg_f <= 0;
    end
    else if (ctrl_reg_wr_en)
    begin
        ctrl_reg_f <= reg_data_in; 
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        coreid_reg_f <= {{(64-34){1'b0}},chipid, coreid_x, coreid_y, 4'd0};
    end
    else if (coreid_reg_wr_en)
    begin
        coreid_reg_f <= reg_data_in; 
    end
end
reg l2_access_counter_inc_en_f;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        l2_access_counter_reg_f <= 0;
    end
    else if (l2_access_counter_reg_wr_en)
    begin
        l2_access_counter_reg_f <= reg_data_in; 
    end
    
    
    
    
    
    l2_access_counter_inc_en_f <= l2_access_counter_inc_en && l2_access_valid;
    if (l2_access_counter_inc_en_f) begin
        l2_access_counter_reg_f <= l2_access_counter_reg_f + 1;
    end
end
reg l2_miss_counter_inc_en_f;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        l2_miss_counter_reg_f <= 0;
    end
    else if (l2_miss_counter_reg_wr_en)
    begin
        l2_miss_counter_reg_f <= reg_data_in; 
    end
    
    
    
    
    
    l2_miss_counter_inc_en_f <= l2_miss_counter_inc_en && l2_miss_valid;
    if (l2_miss_counter_inc_en_f) begin
        l2_miss_counter_reg_f <= l2_miss_counter_reg_f + 1;
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        error_status_reg_f <= 0;
    end
    else if (error_status_reg_wr_en)
    begin
        error_status_reg_f <= reg_data_in; 
    end
    else if (error_status_en && data_ecc_corr_error)
    begin
        if (|error_status_reg_f[1:0])
        begin
            error_status_reg_f <= {error_status_reg_f[63:55], error_addr, data_ecc_addr, 1'b1, 1'b0, 1'b1};
        end
        else
        begin
            error_status_reg_f <= {error_status_reg_f[63:55], error_addr, data_ecc_addr, 1'b0, 1'b0, 1'b1};
        end
    end
    else if (error_status_en && data_ecc_uncorr_error)
    begin
        if (|error_status_reg_f[1:0])
        begin
            error_status_reg_f <= {error_status_reg_f[63:55], error_addr, data_ecc_addr, 1'b1, 1'b1, 1'b0};
        end
        else
        begin
            error_status_reg_f <= {error_status_reg_f[63:55], error_addr, data_ecc_addr, 1'b0, 1'b1, 1'b0};
        end
    end
end
always @ * 
begin
    if (reg_rd_en)
    begin
        if (reg_rd_addr_type == 8'ha9)
        begin
            reg_data_out = ctrl_reg_f;
        end
        else if (reg_rd_addr_type == 8'ha7)
        begin
            reg_data_out = coreid_reg_f;
        end
        else if (reg_rd_addr_type == 8'haa)
        begin
            reg_data_out = l2_access_counter_reg_f;
        end
        else if (reg_rd_addr_type == 8'hab)
        begin
            reg_data_out = l2_miss_counter_reg_f;
        end
        else if (reg_rd_addr_type == 8'ha8)
        begin
            reg_data_out = error_status_reg_f;
        end
        else
        begin
            reg_data_out = 0;
        end
    end
    else
    begin
        reg_data_out = 0;
    end
end
always @ * 
begin
    csm_en = ctrl_reg_f[0];
    error_status_en = ctrl_reg_f[1];
    l2_access_counter_inc_en = ctrl_reg_f[2];
    l2_miss_counter_inc_en = ctrl_reg_f[3];
    smt_base_addr = ctrl_reg_f[22+32-1 : 32];
end
always @ * 
begin
    my_nodeid = coreid_reg_f[34-1 : 0]; 
    core_max = coreid_reg_f[14+8+8+34-1 : 34];
end
endmodule
      
 
module l2_data(
    input wire clk,
    input wire rst_n,
    input wire clk_en,
    input wire rdw_en,
    input wire pdout_en,
    input wire deepsleep,
    input wire [8+2+2-1:0] addr,
    input wire [144-1:0] data_in,
    input wire [144-1:0] data_mask_in,
    output wire [144-1:0] data_out,
    output wire [144-1:0] pdata_out,
    
    output wire [4-1:0] srams_rtap_data,
    input wire  [4-1:0] rtap_srams_bist_command,
    input wire  [4-1:0] rtap_srams_bist_data
);
sram_l2_data l2_data_array(
    .MEMCLK     (clk),
    .RESET_N(rst_n),
    .CE         (clk_en),
    .A          (addr),
    .DIN        (data_in),
    .RDWEN      (rdw_en),
    .BW         (data_mask_in),
    .DOUT       (data_out),
    .BIST_COMMAND(rtap_srams_bist_command),
    .BIST_DIN(rtap_srams_bist_data),
    .BIST_DOUT(srams_rtap_data),
    .SRAMID(8'd13)
);
endmodule
      
 
module l2_data_wrap(
    input wire clk,
    input wire rst_n,
    input wire clk_en1,
    input wire clk_en2,
    input wire rdw_en1,
    input wire rdw_en2,
    input wire pdout_en,
    input wire deepsleep,
    input wire pipe_sel,
    input wire [8+2+2-1:0] addr1,
    input wire [144-1:0] data_in1,
    input wire [144-1:0] data_mask_in1,
    input wire [8+2+2-1:0] addr2,
    input wire [144-1:0] data_in2,
    input wire [144-1:0] data_mask_in2,
    output wire [144-1:0] data_out,
    output wire [144-1:0] pdata_out,
    
    output wire [4-1:0] srams_rtap_data,
    input wire  [4-1:0] rtap_srams_bist_command,
    input wire  [4-1:0] rtap_srams_bist_data
);
reg clk_en;
reg rdw_en;
reg [8+2+2-1:0] addr;
reg [144-1:0] data_in;
reg [144-1:0] data_mask_in;
always @ *
begin
    if (pipe_sel)
    begin
        clk_en = clk_en2;
        rdw_en = rdw_en2;
        addr = addr2;
        data_in = data_in2;
        data_mask_in = data_mask_in2;
    end
    else
    begin
        clk_en = clk_en1;
        rdw_en = rdw_en1;
        addr = addr1;
        data_in = data_in1;
        data_mask_in = data_mask_in1;
    end
end
l2_data l2_data(
    .clk            (clk),
    .rst_n          (rst_n),
    .clk_en         (clk_en),
    .rdw_en         (rdw_en),
    .pdout_en       (pdout_en),
    .deepsleep      (deepsleep),
    .addr           (addr),
    .data_in        (data_in),
    .data_mask_in   (data_mask_in),
    .data_out       (data_out),
    .pdata_out      (pdata_out),
    
    .srams_rtap_data (srams_rtap_data),
    .rtap_srams_bist_command (rtap_srams_bist_command),
    .rtap_srams_bist_data (rtap_srams_bist_data)
);
endmodule
      
 
module l2_decoder(
    input wire [192-1:0] msg_header,
    output reg [8-1:0] msg_type,
    output reg [8-1:0] msg_length,
    output reg [8-1:0] msg_mshrid,
    output reg [3-1:0] msg_data_size,
    output reg [1-1:0] msg_cache_type,
    output reg [4-1:0] msg_subline_vector,
    output reg [2-1:0] msg_mesi,
    output reg [1-1:0] msg_l2_miss,
    output reg [2-1:0] msg_subline_id,
    output reg [1-1:0] msg_last_subline,
    output reg [40-1:0] msg_addr,
    output reg [14-1:0] msg_src_chipid,
    output reg [8-1:0] msg_src_x,
    output reg [8-1:0] msg_src_y,
    output reg [4-1:0] msg_src_fbits,
    output reg [10-1:0] msg_sdid,
    output reg [6-1:0] msg_lsid
);
always @ *
begin
    msg_type = msg_header[21:14];
    msg_length = msg_header[29:22];
    msg_mshrid = msg_header[13:6];
    msg_data_size = msg_header[74:72];
    msg_cache_type = msg_header[75];
    msg_subline_vector = msg_header[79:76];
    msg_mesi = msg_header[5:4];
    msg_l2_miss = msg_header[3];
    msg_subline_id = msg_header[2:1];
    msg_last_subline = msg_header[0];
    msg_addr = msg_header[119:80];
    msg_src_chipid = msg_header[191:178];
    msg_src_x = msg_header[177:170];
    msg_src_y = msg_header[169:162];
    msg_src_fbits = msg_header[161:158];
    msg_sdid = msg_header[157:148];
    msg_lsid = msg_header[147:142];
end
endmodule
      
 
module l2_dir(
    input wire clk,
    input wire rst_n,
    input wire clk_en,
    input wire rdw_en,
    input wire pdout_en,
    input wire deepsleep,
    input wire [8+2-1:0] addr,
    input wire [64-1:0] data_in,
    input wire [64-1:0] data_mask_in,
    output wire [64-1:0] data_out,
    output wire [64-1:0] pdata_out,
    
    output wire [4-1:0] srams_rtap_data,
    input wire  [4-1:0] rtap_srams_bist_command,
    input wire  [4-1:0] rtap_srams_bist_data
);
sram_l2_dir l2_dir_array(
    .MEMCLK     (clk),
    .RESET_N(rst_n),
    .CE         (clk_en),
    .A          (addr),
    .DIN        (data_in),
    .RDWEN      (rdw_en),
    .BW         (data_mask_in),
    .DOUT       (data_out),
    .BIST_COMMAND(rtap_srams_bist_command),
    .BIST_DIN(rtap_srams_bist_data),
    .BIST_DOUT(srams_rtap_data),
    .SRAMID(8'd14)
);
endmodule
      
 
module l2_dir_wrap(
    input wire clk,
    input wire rst_n,
    input wire clk_en1,
    input wire clk_en2,
    input wire rdw_en1,
    input wire rdw_en2,
    input wire pdout_en,
    input wire deepsleep,
    input wire pipe_sel,
    input wire [8+2-1:0] addr1,
    input wire [64-1:0] data_in1,
    input wire [64-1:0] data_mask_in1,
    input wire [8+2-1:0] addr2,
    input wire [64-1:0] data_in2,
    input wire [64-1:0] data_mask_in2,
    output wire [64-1:0] data_out,
    output wire [64-1:0] pdata_out,
    
    output wire [4-1:0] srams_rtap_data,
    input wire  [4-1:0] rtap_srams_bist_command,
    input wire  [4-1:0] rtap_srams_bist_data
);
reg clk_en;
reg rdw_en;
reg [8+2-1:0] addr;
reg [64-1:0] data_in;
reg [64-1:0] data_mask_in;
always @ *
begin
    if (pipe_sel)
    begin
        clk_en = clk_en2;
        rdw_en = rdw_en2;
        addr = addr2;
        data_in = data_in2;
        data_mask_in = data_mask_in2;
    end
    else
    begin
        clk_en = clk_en1;
        rdw_en = rdw_en1;
        addr = addr1;
        data_in = data_in1;
        data_mask_in = data_mask_in1;
    end
end
l2_dir l2_dir(
    .clk            (clk),
    .rst_n          (rst_n),
    .clk_en         (clk_en),
    .rdw_en         (rdw_en),
    .pdout_en       (pdout_en),
    .deepsleep      (deepsleep),
    .addr           (addr),
    .data_in        (data_in),
    .data_mask_in   (data_mask_in),
    .data_out       (data_out),
    .pdata_out      (pdata_out),
    
    .srams_rtap_data (srams_rtap_data),
    .rtap_srams_bist_command (rtap_srams_bist_command),
    .rtap_srams_bist_data (rtap_srams_bist_data)
);
endmodule
      
 
module l2_encoder(
    input wire [14-1:0] msg_dst_chipid,
    input wire [8-1:0] msg_dst_x,
    input wire [8-1:0] msg_dst_y,
    input wire [4-1:0] msg_dst_fbits,
    input wire [8-1:0] msg_length,
    input wire [8-1:0] msg_type,
    input wire [8-1:0] msg_mshrid,
    input wire [3-1:0] msg_data_size,
    input wire [1-1:0] msg_cache_type,
    input wire [4-1:0] msg_subline_vector,
    input wire [2-1:0] msg_mesi,
    input wire [1-1:0] msg_l2_miss,
    input wire [1-1:0] msg_last_subline,
    input wire [2-1:0] msg_subline_id,
    input wire [40-1:0] msg_addr,
    input wire [14-1:0] msg_src_chipid,
    input wire [8-1:0] msg_src_x,
    input wire [8-1:0] msg_src_y,
    input wire [4-1:0] msg_src_fbits,
    input wire [10-1:0] msg_sdid,
    input wire [6-1:0] msg_lsid,
    output reg [192-1:0] msg_header
);
always @ *
begin
    msg_header = {msg_src_chipid,
                  msg_src_x,
                  msg_src_y,
                  msg_src_fbits,
                  msg_sdid,
                  msg_lsid,
                  14'd0,
                  8'd0,
                  msg_addr,
                  msg_subline_vector,
                  msg_cache_type,
                  msg_data_size,
                  8'd0,
                  msg_dst_chipid,
                  msg_dst_x,
                  msg_dst_y,
                  msg_dst_fbits,
                  msg_length,
                  msg_type,
                  msg_mshrid,
                  msg_mesi,
                  msg_l2_miss,
                  msg_subline_id,
                  msg_last_subline};
end
endmodule
      
 
module l2_mshr_decoder(
    input wire [120+2-1:0] data_in,
    output reg [40-1:0] addr_out,
    output reg [2-1:0] way_out,
    output reg [8-1:0] mshrid_out,
    output reg [1-1:0] cache_type_out,
    output reg [3-1:0] data_size_out,
    output reg [8-1:0] msg_type_out,
    output reg [1-1:0] msg_l2_miss_out,
    output reg [14-1:0] src_chipid_out,
    output reg [8-1:0] src_x_out,
    output reg [8-1:0] src_y_out,
    output reg [4-1:0] src_fbits_out,
    output reg [10-1:0] sdid_out,
    output reg [6-1:0] lsid_out,
    output reg [6-1:0] miss_lsid_out,
    output reg smc_miss_out,
    output reg recycled,
    output reg inv_fwd_pending
);
always @ *
begin
    addr_out = data_in[39:0];
    way_out = data_in[39+2:40];
    mshrid_out = data_in[47+2:40+2];
    cache_type_out = data_in[48+2];
    data_size_out = data_in[51+2:49+2];
    msg_type_out = data_in[59+2:52+2];
    msg_l2_miss_out = data_in[60+2];
    src_chipid_out = data_in[74+2:61+2];
    src_x_out = data_in[82+2:75+2];
    src_y_out = data_in[90+2:83+2];
    src_fbits_out = data_in[94+2:91+2];
    sdid_out = data_in[104+2:95+2];
    lsid_out = data_in[110+2:105+2];
    miss_lsid_out = data_in[116+2:111+2];
    smc_miss_out = data_in[117+2];
    recycled = data_in[118+2];
    inv_fwd_pending = data_in[119+2];
end
endmodule
      
 
module l2_pipe1(
    input wire clk,
    input wire rst_n,
    input wire [34-1:0] my_nodeid,
    
    input wire csm_en,
    
    input wire [22-1:0] smt_base_addr,
  
   
   
    input wire noc_valid_in,
    input wire [64-1:0] noc_data_in,
    output wire noc_ready_in,
    
    
   
    output wire noc_valid_out,
    output wire [64-1:0] noc_data_out,
    input wire  noc_ready_out,
    input wire pipe2_valid_S1,
    input wire pipe2_valid_S2,
    input wire pipe2_valid_S3,
    input wire [8-1:0] pipe2_msg_type_S1,
    input wire [8-1:0] pipe2_msg_type_S2,
    input wire [8-1:0] pipe2_msg_type_S3,
    input wire [40-1:0] pipe2_addr_S1,
    input wire [40-1:0] pipe2_addr_S2,
    input wire [40-1:0] pipe2_addr_S3,
    input wire global_stall_S1,
    input wire global_stall_S2,
    input wire global_stall_S4,
    input wire mshr_hit,
    input wire [120+2-1:0] cam_mshr_data_out,
    input wire [120+2-1:0] pending_mshr_data_out,
 
    input wire [6-1:0] mshr_inv_counter_out,
    input wire [3:0] mshr_empty_slots,
    input wire mshr_pending,
    input wire [3-1:0] mshr_pending_index,
    input wire [3-1:0] mshr_empty_index,
    
    input wire broadcast_counter_zero,
    input wire broadcast_counter_max,
    input wire broadcast_counter_avail,
    input wire [14-1:0] broadcast_chipid_out,
    input wire [8-1:0] broadcast_x_out,
    input wire [8-1:0] broadcast_y_out,
    
    input wire [15*4+2+4-1:0] state_data_out,
    
    input wire [104-1:0] tag_data_out,
    input wire [64-1:0] dir_data_out,
    input wire [144-1:0] data_data_out,
    
    input wire smc_hit,
    input wire [30-1:0] smc_data_out,
    input wire [4-1:0] smc_valid_out,
    input wire [14-1:0] smc_tag_out,
    
    input wire [64-1:0] reg_data_out,
    output wire mshr_cam_en,
    output wire mshr_wr_state_en,
    output wire mshr_wr_data_en,
    output wire mshr_pending_ready,
    output wire [2-1:0] mshr_state_in,
    output wire [120+2-1:0] mshr_data_in,
    output wire [120+2-1:0] mshr_data_mask_in,
    output wire [3-1:0] mshr_inv_counter_rd_index_in,
    output wire [3-1:0] mshr_wr_index_in,
    output wire [8-1:0] mshr_addr_in,
    output wire state_rd_en,
    output wire state_wr_en,
    output wire [8-1:0] state_rd_addr,
    output wire [8-1:0] state_wr_addr,
    output wire [15*4+2+4-1:0] state_data_in,
    output wire [15*4+2+4-1:0] state_data_mask_in,
    output wire tag_clk_en,
    output wire tag_rdw_en,
    output wire [8-1:0] tag_addr,
    output wire [104-1:0] tag_data_in,
    output wire [104-1:0] tag_data_mask_in,
    output wire dir_clk_en,
    output wire dir_rdw_en,
    output wire [8+2-1:0] dir_addr,
    output wire [64-1:0] dir_data_in,
    output wire [64-1:0] dir_data_mask_in,
    output wire data_clk_en,
    output wire data_rdw_en,
    output wire [8+2+2-1:0] data_addr,
    output wire [144-1:0] data_data_in,
    output wire [144-1:0] data_data_mask_in,
    
    output wire [2-1:0] broadcast_counter_op,
    output wire broadcast_counter_op_val,
    
    
    output wire smc_rd_en,
    output wire [16-1:0] smc_rd_addr_in,
    output wire smc_rd_diag_en,
    output wire smc_flush_en,
    output wire [2-1:0] smc_addr_op,
    output wire smc_wr_en,
    output wire smc_wr_diag_en,
    output wire [16-1:0] smc_wr_addr_in,
    output wire [128-1:0] smc_data_in,
    
    output wire l2_access_valid,
    output wire l2_miss_valid,
    output wire data_ecc_corr_error,
    output wire data_ecc_uncorr_error,
    output wire [8+2+2-1:0] data_ecc_addr,
    output wire [40-1:0] error_addr,
    output wire reg_rd_en,
    output wire reg_wr_en,
    output wire [8-1:0] reg_rd_addr_type,
    output wire [8-1:0] reg_wr_addr_type,
    output wire [64-1:0] reg_data_in
);
wire [8-1:0] msg_type;
wire [8-1:0] msg_length;
wire [8-1:0] msg_mshrid;
wire [3-1:0] msg_data_size;
wire [1-1:0] msg_cache_type;
wire [40-1:0] msg_addr;
wire [14-1:0] msg_src_chipid;
wire [8-1:0] msg_src_x;
wire [8-1:0] msg_src_y;
wire [4-1:0] msg_src_fbits;
wire [10-1:0] msg_sdid;
wire [6-1:0] msg_lsid;
wire [8-1:0] cam_mshr_msg_type;
wire [8-1:0] cam_mshr_mshrid;
wire [3-1:0] cam_mshr_data_size;
wire [1-1:0] cam_mshr_cache_type;
wire [40-1:0] cam_mshr_addr;
wire [2-1:0] cam_mshr_way;
wire [1-1:0] cam_mshr_l2_miss;
wire [14-1:0] cam_mshr_src_chipid;
wire [8-1:0] cam_mshr_src_x;
wire [8-1:0] cam_mshr_src_y;
wire [4-1:0] cam_mshr_src_fbits;
wire [10-1:0] cam_mshr_sdid;
wire [6-1:0] cam_mshr_lsid;
wire [6-1:0] cam_mshr_miss_lsid;
 
wire cam_mshr_smc_miss;
 
wire cam_mshr_recycled;
wire [8-1:0] pending_mshr_msg_type;
wire [8-1:0] pending_mshr_mshrid;
wire [3-1:0] pending_mshr_data_size;
wire [1-1:0] pending_mshr_cache_type;
wire [40-1:0] pending_mshr_addr;
wire [2-1:0] pending_mshr_way;
wire [1-1:0] pending_mshr_l2_miss;
wire [14-1:0] pending_mshr_src_chipid;
wire [8-1:0] pending_mshr_src_x;
wire [8-1:0] pending_mshr_src_y;
wire [4-1:0] pending_mshr_src_fbits;
wire [10-1:0] pending_mshr_sdid;
wire [6-1:0] pending_mshr_lsid;
wire [6-1:0] pending_mshr_miss_lsid;
wire pending_mshr_smc_miss;
wire pending_mshr_recycled;
 
wire msg_header_valid;
wire [192-1:0] msg_header;
wire msg_header_ready;
wire msg_data_valid;
wire [64-1:0] msg_data;
wire msg_data_ready;
wire valid_S1; 
wire stall_S1;  
wire msg_from_mshr_S1;
wire [40-1:0] addr_S1;
wire dis_flush_S1;
wire [4-1:0] amo_alu_op_S2;
wire valid_S2; 
wire stall_S2;  
wire stall_before_S2; 
wire stall_real_S2; 
wire msg_from_mshr_S2;
wire [8-1:0] msg_type_S2;
wire [3-1:0] data_size_S2;
wire [1-1:0] cache_type_S2;
wire state_owner_en_S2;
wire [2-1:0] state_owner_op_S2;
wire state_subline_en_S2;
wire [2-1:0] state_subline_op_S2;
wire state_di_en_S2;
wire state_vd_en_S2;
wire [2-1:0] state_vd_S2;
wire state_mesi_en_S2;
wire [2-1:0] state_mesi_S2;
wire state_lru_en_S2;
wire [1-1:0] state_lru_op_S2;
wire state_rb_en_S2;
wire l2_ifill_32B_S2;
wire [2-1:0] l2_load_data_subline_S2;
wire [40-1:0] addr_S2;
wire l2_tag_hit_S2;
wire l2_evict_S2;
wire l2_wb_S2;
wire [2-1:0] l2_way_state_mesi_S2;
wire [2-1:0] l2_way_state_vd_S2;
wire [1-1:0] l2_way_state_cache_type_S2;
wire [4-1:0] l2_way_state_subline_S2;
wire [2-1:0] dir_op_S2;
wire req_from_owner_S2;
wire addr_l2_aligned_S2;
wire special_addr_type_S2;
wire [6-1:0] lsid_S2;
wire state_load_sdid_S2;
wire valid_S3; 
wire stall_S3;  
wire stall_before_S3; 
wire [40-1:0] addr_S3;
wire valid_S4;    
wire stall_S4;
wire stall_before_S4; 
wire [6-1:0] dir_sharer_S4;
wire [6-1:0] dir_sharer_counter_S4;
wire cas_cmp_en_S4;
wire [3-1:0] cas_cmp_data_size_S4;
wire [40-1:0] addr_S4;
wire l2_evict_S4;
wire l2_tag_hit_S4;
wire [2-1:0] l2_way_state_mesi_S4;
wire [6-1:0] l2_way_state_owner_S4;
wire [2-1:0] l2_way_state_vd_S4;
wire [4-1:0] l2_way_state_subline_S4;
wire [1-1:0] l2_way_state_cache_type_S4;
wire [8-1:0] mshrid_S4;
wire req_from_owner_S4;
wire cas_cmp_S4;
wire atomic_read_data_en_S4;
wire [8-1:0] msg_type_S4;
wire [3-1:0] data_size_S4;
wire [1-1:0] cache_type_S4;
wire [1-1:0] l2_miss_S4;
wire [6-1:0] mshr_miss_lsid_S4;
wire [6-1:0] lsid_S4;
wire special_addr_type_S4;
wire state_wr_sel_S4;
wire [64-1:0] dir_data_S4;
wire [64-1:0] dir_data_sel_S4;
wire smc_miss_S4;
wire stall_smc_buf_S4;
    
wire msg_from_mshr_S4;
wire req_recycle_S4;
wire inv_fwd_pending_S4;
wire msg_send_valid;
wire msg_send_ready;
wire [3-1:0] msg_send_mode;
wire [8-1:0] msg_send_type;
wire [8-1:0] msg_send_type_pre;
wire [8-1:0] msg_send_length;
wire [3-1:0] msg_send_data_size;
wire [1-1:0] msg_send_cache_type;
wire [1-1:0] msg_send_l2_miss;
wire [2-1:0] msg_send_mesi;
wire [8-1:0] msg_send_mshrid;
wire [4-1:0] msg_send_subline_vector;
wire [40-1:0] msg_send_addr;
wire [14-1:0] msg_send_dst_chipid;
wire [8-1:0] msg_send_dst_x;
wire [8-1:0] msg_send_dst_y;
wire [4-1:0] msg_send_dst_fbits;
wire [64*2-1:0] msg_send_data;
wire [64*3-1:0] msg_send_header;
assign error_addr = addr_S4;
l2_pipe1_buf_in buf_in(
    .clk                    (clk),
    .rst_n                  (rst_n),
    .valid_in               (noc_valid_in),
    .data_in                (noc_data_in),
    .ready_in               (noc_ready_in),
    .msg_header_valid_out   (msg_header_valid),
    .msg_header_out         (msg_header),
    .msg_header_ready_out   (msg_header_ready),
    .msg_data_valid_out     (msg_data_valid),
    .msg_data_out           (msg_data),
    .msg_data_ready_out     (msg_data_ready)
);
l2_decoder decoder(
    .msg_header         (msg_header),
    .msg_type           (msg_type),
    .msg_length         (msg_length),
    .msg_mshrid         (msg_mshrid),
    .msg_data_size      (msg_data_size),
    .msg_cache_type     (msg_cache_type),
    .msg_subline_vector (),
    .msg_mesi           (),
    .msg_l2_miss        (),
    .msg_subline_id     (),
    .msg_last_subline   (),
    .msg_addr           (msg_addr),
    .msg_src_chipid     (msg_src_chipid),
    .msg_src_x          (msg_src_x),
    .msg_src_y          (msg_src_y),
    .msg_src_fbits      (msg_src_fbits),
    .msg_sdid           (msg_sdid),
    .msg_lsid           (msg_lsid)
);
    
    
    
l2_mshr_decoder cam_mshr_decoder(
    
    
    .data_in            (cam_mshr_data_out),
    .addr_out           (cam_mshr_addr),
    .way_out            (cam_mshr_way),
    .mshrid_out         (cam_mshr_mshrid),
    .cache_type_out     (cam_mshr_cache_type), 
    .data_size_out      (cam_mshr_data_size),
    .msg_type_out       (cam_mshr_msg_type),
    .msg_l2_miss_out    (cam_mshr_l2_miss),
    .src_chipid_out     (cam_mshr_src_chipid),
    .src_x_out          (cam_mshr_src_x),
    .src_y_out          (cam_mshr_src_y),
    .src_fbits_out      (cam_mshr_src_fbits),
    .sdid_out           (cam_mshr_sdid),
    .lsid_out           (cam_mshr_lsid),
    .miss_lsid_out      (cam_mshr_miss_lsid),
    
    .smc_miss_out       (cam_mshr_smc_miss),
    
    
    .recycled           (cam_mshr_recycled),
    .inv_fwd_pending    ()
);
l2_mshr_decoder pending_mshr_decoder(
    
    
    .data_in            (pending_mshr_data_out),
    .addr_out           (pending_mshr_addr),
    .way_out            (pending_mshr_way),
    .mshrid_out         (pending_mshr_mshrid),
    .cache_type_out     (pending_mshr_cache_type), 
    .data_size_out      (pending_mshr_data_size),
    .msg_type_out       (pending_mshr_msg_type),
    .msg_l2_miss_out    (pending_mshr_l2_miss),
    .src_chipid_out     (pending_mshr_src_chipid),
    .src_x_out          (pending_mshr_src_x),
    .src_y_out          (pending_mshr_src_y),
    .src_fbits_out      (pending_mshr_src_fbits),
    .sdid_out           (pending_mshr_sdid),
    .lsid_out           (pending_mshr_lsid),
    .miss_lsid_out      (pending_mshr_miss_lsid),
    
    .smc_miss_out       (pending_mshr_smc_miss),
    
    
    .recycled           (pending_mshr_recycled),
    .inv_fwd_pending    ()
);
 
l2_pipe1_ctrl ctrl(
    .clk                        (clk),
    .rst_n                      (rst_n),
    
    .csm_en                     (csm_en),
    
    .pipe2_valid_S1             (pipe2_valid_S1),
    .pipe2_valid_S2             (pipe2_valid_S2),
    .pipe2_valid_S3             (pipe2_valid_S3),
    .pipe2_msg_type_S1          (pipe2_msg_type_S1),
    .pipe2_msg_type_S2          (pipe2_msg_type_S2),
    .pipe2_msg_type_S3          (pipe2_msg_type_S3),
    .pipe2_addr_S1              (pipe2_addr_S1),
    .pipe2_addr_S2              (pipe2_addr_S2),
    .pipe2_addr_S3              (pipe2_addr_S3),
    .global_stall_S1            (global_stall_S1),
    .msg_header_valid_S1        (msg_header_valid),
    .msg_type_S1                (msg_type),
    .msg_data_size_S1           (msg_data_size),
    .msg_cache_type_S1          (msg_cache_type),
    .mshr_hit_S1                (mshr_hit),
    .cam_mshr_msg_type_S1       (cam_mshr_msg_type),
    .cam_mshr_l2_miss_S1        (cam_mshr_l2_miss),
    .cam_mshr_data_size_S1      (cam_mshr_data_size),
    .cam_mshr_cache_type_S1     (cam_mshr_cache_type), 
 
    .mshr_pending_S1            (mshr_pending),
    .mshr_pending_index_S1      (mshr_pending_index),
    .mshr_empty_slots_S1        (mshr_empty_slots),
    
    .cam_mshr_smc_miss_S1       (cam_mshr_smc_miss),
 
    
    .pending_mshr_msg_type_S1           (pending_mshr_msg_type),
    .pending_mshr_l2_miss_S1            (pending_mshr_l2_miss),
    .pending_mshr_data_size_S1          (pending_mshr_data_size),
    .pending_mshr_cache_type_S1         (pending_mshr_cache_type), 
    
    .pending_mshr_smc_miss_S1           (pending_mshr_smc_miss),
    
 
    .msg_data_valid_S1          (msg_data_valid),
    .addr_S1                    (addr_S1),
   
    .global_stall_S2            (global_stall_S2),
    .l2_tag_hit_S2              (l2_tag_hit_S2),
    .l2_evict_S2                (l2_evict_S2),
    .l2_wb_S2                   (l2_wb_S2),
    .l2_way_state_mesi_S2       (l2_way_state_mesi_S2),
    .l2_way_state_vd_S2         (l2_way_state_vd_S2),
    .l2_way_state_cache_type_S2 (l2_way_state_cache_type_S2),
    .l2_way_state_subline_S2    (l2_way_state_subline_S2),
    .req_from_owner_S2          (req_from_owner_S2),
    .addr_l2_aligned_S2         (addr_l2_aligned_S2),
    .lsid_S2                    (lsid_S2),
    .msg_data_valid_S2          (msg_data_valid),
    .addr_S2                    (addr_S2),
    .dir_data_S3                (dir_data_out),
    .addr_S3                    (addr_S3),
    .global_stall_S4            (global_stall_S4),
    .l2_evict_S4                (l2_evict_S4),
    .l2_tag_hit_S4              (l2_tag_hit_S4),
    .l2_way_state_mesi_S4       (l2_way_state_mesi_S4),
    .l2_way_state_owner_S4      (l2_way_state_owner_S4),
    .l2_way_state_vd_S4         (l2_way_state_vd_S4),
    .l2_way_state_subline_S4    (l2_way_state_subline_S4),
    .l2_way_state_cache_type_S4 (l2_way_state_cache_type_S4),
    .mshrid_S4                  (mshrid_S4),
    .req_from_owner_S4          (req_from_owner_S4),
    .mshr_miss_lsid_S4          (mshr_miss_lsid_S4),
    .lsid_S4                    (lsid_S4),
    .addr_S4                    (addr_S4),
    .cas_cmp_S4                 (cas_cmp_S4),
    .msg_send_ready_S4          (msg_send_ready),
    .mshr_empty_index_S4        (mshr_empty_index),
    
    
    .smc_hit_S4                 (smc_hit),
    .broadcast_counter_zero_S4  (broadcast_counter_zero),
    .broadcast_counter_max_S4   (broadcast_counter_max),
    .broadcast_counter_avail_S4 (broadcast_counter_avail),
    .broadcast_chipid_out_S4    (broadcast_chipid_out),
    .broadcast_x_out_S4         (broadcast_x_out),
    .broadcast_y_out_S4         (broadcast_y_out),
    
    .valid_S1                   (valid_S1),  
    .stall_S1                   (stall_S1),    
    .msg_from_mshr_S1           (msg_from_mshr_S1), 
    .dis_flush_S1               (dis_flush_S1),
    .mshr_cam_en_S1             (mshr_cam_en),
    .mshr_pending_ready_S1      (mshr_pending_ready),
    .msg_header_ready_S1        (msg_header_ready),
    .tag_clk_en_S1              (tag_clk_en),
    .tag_rdw_en_S1              (tag_rdw_en),
    .state_rd_en_S1             (state_rd_en),
    .reg_wr_en_S1               (reg_wr_en),
    .reg_wr_addr_type_S1        (reg_wr_addr_type),
    .valid_S2                   (valid_S2),    
    .stall_S2                   (stall_S2), 
    .stall_before_S2            (stall_before_S2), 
    .stall_real_S2              (stall_real_S2),
    .msg_type_S2                (msg_type_S2),
    .msg_from_mshr_S2           (msg_from_mshr_S2),
    .special_addr_type_S2       (special_addr_type_S2),
    .dir_clk_en_S2              (dir_clk_en),
    .dir_rdw_en_S2              (dir_rdw_en),
    .dir_op_S2                  (dir_op_S2),
    .data_clk_en_S2             (data_clk_en),
    .data_rdw_en_S2             (data_rdw_en),
    .amo_alu_op_S2              (amo_alu_op_S2),
    .data_size_S2               (data_size_S2),
    .cache_type_S2              (cache_type_S2),
    .state_owner_en_S2          (state_owner_en_S2),
    .state_owner_op_S2          (state_owner_op_S2),
    .state_subline_en_S2        (state_subline_en_S2),
    .state_subline_op_S2        (state_subline_op_S2),   
    .state_di_en_S2             (state_di_en_S2),
    .state_vd_en_S2             (state_vd_en_S2),
    .state_vd_S2                (state_vd_S2),
    .state_mesi_en_S2           (state_mesi_en_S2),
    .state_mesi_S2              (state_mesi_S2),
    .state_lru_en_S2            (state_lru_en_S2),
    .state_lru_op_S2            (state_lru_op_S2),
    .state_rb_en_S2             (state_rb_en_S2),
    .state_load_sdid_S2         (state_load_sdid_S2),
    .l2_ifill_32B_S2            (l2_ifill_32B_S2),
    .l2_load_data_subline_S2    (l2_load_data_subline_S2),
    .msg_data_ready_S2          (msg_data_ready),
    
    .smc_wr_en_S2               (smc_wr_en),
    .smc_wr_diag_en_S2          (smc_wr_diag_en),
    .smc_flush_en_S2            (smc_flush_en),
    .smc_addr_op_S2             (smc_addr_op),
        
    .valid_S3                   (valid_S3),    
    .stall_S3                   (stall_S3), 
    .stall_before_S3            (stall_before_S3), 
    .valid_S4                   (valid_S4),    
    .stall_S4                   (stall_S4), 
    .stall_before_S4            (stall_before_S4),
     
    .stall_smc_buf_S4           (stall_smc_buf_S4),
    
    .msg_from_mshr_S4           (msg_from_mshr_S4),
    .req_recycle_S4             (req_recycle_S4),
    .inv_fwd_pending_S4         (inv_fwd_pending_S4),
    .dir_sharer_S4              (dir_sharer_S4),
    .dir_sharer_counter_S4      (dir_sharer_counter_S4),
    .cas_cmp_en_S4              (cas_cmp_en_S4),
    .atomic_read_data_en_S4     (atomic_read_data_en_S4),
    .cas_cmp_data_size_S4       (cas_cmp_data_size_S4),
    .msg_send_valid_S4          (msg_send_valid),
    .msg_send_mode_S4           (msg_send_mode),
    .msg_send_type_S4           (msg_send_type),
    .msg_send_type_pre_S4       (msg_send_type_pre),
    .msg_send_length_S4         (msg_send_length),
    .msg_send_data_size_S4      (msg_send_data_size),
    .msg_send_cache_type_S4     (msg_send_cache_type),
    .msg_send_mesi_S4           (msg_send_mesi),
    .msg_send_l2_miss_S4        (msg_send_l2_miss),
    .msg_send_mshrid_S4         (msg_send_mshrid),
    .msg_send_subline_vector_S4 (msg_send_subline_vector),
    .special_addr_type_S4       (special_addr_type_S4),
    .dir_data_sel_S4            (dir_data_sel_S4),
    .dir_data_S4                (dir_data_S4),
    .msg_type_S4                (msg_type_S4),
    .data_size_S4               (data_size_S4),
    .cache_type_S4              (cache_type_S4),
    .l2_miss_S4                 (l2_miss_S4),
    
    .smc_miss_S4                (smc_miss_S4),
    
    .mshr_wr_data_en_S4         (mshr_wr_data_en),
    .mshr_wr_state_en_S4        (mshr_wr_state_en),
    .mshr_state_in_S4           (mshr_state_in),
    .mshr_wr_index_in_S4        (mshr_wr_index_in),    
    .mshr_inv_counter_rd_index_in_S4(mshr_inv_counter_rd_index_in),    
    .state_wr_sel_S4            (state_wr_sel_S4),
    .state_wr_en_S4             (state_wr_en),
    
    .broadcast_counter_op_S4    (broadcast_counter_op),
    .broadcast_counter_op_val_S4(broadcast_counter_op_val),
    
    
    
    .smc_rd_diag_en_buf_S4      (smc_rd_diag_en),
    .smc_rd_en_buf_S4           (smc_rd_en),
    
    .l2_access_valid_S4         (l2_access_valid),
    .l2_miss_valid_S4           (l2_miss_valid),
    .reg_rd_en_S4               (reg_rd_en),
    .reg_rd_addr_type_S4        (reg_rd_addr_type)
);
l2_pipe1_dpath dpath(
    .clk                        (clk),
    .rst_n                      (rst_n),
    
    .csm_en                     (csm_en),
    
    .smt_base_addr              (smt_base_addr),
    
    .cam_mshr_addr_S1           (cam_mshr_addr),
    .cam_mshr_mshrid_S1         (cam_mshr_mshrid),
    .cam_mshr_way_S1            (cam_mshr_way),
    .cam_mshr_src_chipid_S1     (cam_mshr_src_chipid),
    .cam_mshr_src_x_S1          (cam_mshr_src_x),
    .cam_mshr_src_y_S1          (cam_mshr_src_y),
    .cam_mshr_src_fbits_S1      (cam_mshr_src_fbits),
    .cam_mshr_sdid_S1           (cam_mshr_sdid),
    .cam_mshr_lsid_S1           (cam_mshr_lsid),
    .cam_mshr_miss_lsid_S1      (cam_mshr_miss_lsid),
    .cam_mshr_recycled_S1       (cam_mshr_recycled),
    
    .mshr_pending_S1            (mshr_pending),
    .pending_mshr_addr_S1       (pending_mshr_addr),
    .pending_mshr_mshrid_S1     (pending_mshr_mshrid),
    .pending_mshr_way_S1        (pending_mshr_way),
    .pending_mshr_src_chipid_S1 (pending_mshr_src_chipid),
    .pending_mshr_src_x_S1      (pending_mshr_src_x),
    .pending_mshr_src_y_S1      (pending_mshr_src_y),
    .pending_mshr_src_fbits_S1  (pending_mshr_src_fbits),
    .pending_mshr_sdid_S1       (pending_mshr_sdid),
    .pending_mshr_lsid_S1       (pending_mshr_lsid),
    .pending_mshr_miss_lsid_S1  (pending_mshr_miss_lsid),
    .pending_mshr_recycled_S1   (pending_mshr_recycled),
 
    .dis_flush_S1               (dis_flush_S1),
    .msg_addr_S1                (msg_addr),
    .msg_mshrid_S1              (msg_mshrid),
    .msg_src_chipid_S1          (msg_src_chipid),
    .msg_src_x_S1               (msg_src_x),
    .msg_src_y_S1               (msg_src_y),
    .msg_src_fbits_S1           (msg_src_fbits),
    .msg_sdid_S1                (msg_sdid),
    .msg_lsid_S1                (msg_lsid),
    .msg_data_S1                (msg_data),
    .valid_S1                   (valid_S1),
    .stall_S1                   (stall_S1),
    .msg_from_mshr_S1           (msg_from_mshr_S1), 
    .state_data_S2              (state_data_out),
    .tag_data_S2                (tag_data_out),
    .msg_data_S2                (msg_data),
    .msg_type_S2                (msg_type_S2),
    .msg_from_mshr_S2           (msg_from_mshr_S2),
    .special_addr_type_S2       (special_addr_type_S2),
    .data_size_S2               (data_size_S2),
    .cache_type_S2              (cache_type_S2),
    .state_owner_en_S2          (state_owner_en_S2),
    .state_owner_op_S2          (state_owner_op_S2), 
    .state_subline_en_S2        (state_subline_en_S2),
    .state_subline_op_S2        (state_subline_op_S2),
    .state_di_en_S2             (state_di_en_S2),
    .state_vd_en_S2             (state_vd_en_S2),
    .state_vd_S2                (state_vd_S2),
    .state_mesi_en_S2           (state_mesi_en_S2),
    .state_mesi_S2              (state_mesi_S2),
    .state_lru_en_S2            (state_lru_en_S2),
    .state_lru_op_S2            (state_lru_op_S2),
    .state_rb_en_S2             (state_rb_en_S2),
    .state_load_sdid_S2         (state_load_sdid_S2),
    .dir_op_S2                  (dir_op_S2),
    .l2_ifill_32B_S2            (l2_ifill_32B_S2),
    .l2_load_data_subline_S2    (l2_load_data_subline_S2),
    .valid_S2                   (valid_S2),
    .stall_S2                   (stall_S2),
    .stall_before_S2            (stall_before_S2), 
    .data_clk_en_S2             (data_clk_en),
    .stall_real_S2              (stall_real_S2),
    .amo_alu_op_S2              (amo_alu_op_S2),
    .valid_S3                   (valid_S3),
    .stall_S3                   (stall_S3),
    .stall_before_S3            (stall_before_S3), 
    .data_data_S3               (data_data_out),
    .valid_S4                   (valid_S4),
    .stall_S4                   (stall_S4),
    .stall_before_S4            (stall_before_S4),
     
    .stall_smc_buf_S4           (stall_smc_buf_S4),
    
    .msg_from_mshr_S4           (msg_from_mshr_S4),
    .req_recycle_S4             (req_recycle_S4),
    .inv_fwd_pending_S4         (inv_fwd_pending_S4),
    .cas_cmp_en_S4              (cas_cmp_en_S4),    
    .atomic_read_data_en_S4     (atomic_read_data_en_S4),
    .cas_cmp_data_size_S4       (cas_cmp_data_size_S4),
    .dir_sharer_S4              (dir_sharer_S4),
    .dir_sharer_counter_S4      (dir_sharer_counter_S4),
    .mshr_inv_counter_out_S4    (mshr_inv_counter_out),
    .special_addr_type_S4       (special_addr_type_S4),
    .dir_data_sel_S4            (dir_data_sel_S4),
    .dir_data_S4                (dir_data_S4),
    .msg_send_type_S4           (msg_send_type),
    .msg_send_length_S4         (msg_send_length),
    .my_nodeid_chipid_S4        (my_nodeid[33:20]),
    .my_nodeid_x_S4             (my_nodeid[19:12]),
    .my_nodeid_y_S4             (my_nodeid[11:4]),
    .state_wr_sel_S4            (state_wr_sel_S4),
    .msg_type_S4                (msg_type_S4),
    .msg_send_type_pre_S4       (msg_send_type_pre),
    .data_size_S4               (data_size_S4),
    .cache_type_S4              (cache_type_S4),
    .l2_miss_S4                 (l2_miss_S4),
    
    .smc_miss_S4                (smc_miss_S4),
    .smc_data_out_S4            (smc_data_out),
    .smc_valid_out_S4           (smc_valid_out),
    .smc_tag_out_S4             (smc_tag_out),
    
    .reg_data_out_S4            (reg_data_out),
    
    .broadcast_chipid_out_S4    (broadcast_chipid_out),
    .broadcast_x_out_S4         (broadcast_x_out),
    .broadcast_y_out_S4         (broadcast_y_out),
    
 
    .addr_S1                    (addr_S1),
    .mshr_addr_in_S1            (mshr_addr_in),
    .tag_addr_S1                (tag_addr),
    .tag_data_in_S1             (tag_data_in),  
    .tag_data_mask_in_S1        (tag_data_mask_in),
    .state_rd_addr_S1           (state_rd_addr),
    .reg_data_in_S1             (reg_data_in),
    .addr_S2                    (addr_S2),
    .l2_tag_hit_S2              (l2_tag_hit_S2),
    .l2_evict_S2                (l2_evict_S2),
    .l2_wb_S2                   (l2_wb_S2),
    .l2_way_state_mesi_S2       (l2_way_state_mesi_S2),
    .l2_way_state_vd_S2         (l2_way_state_vd_S2),    
    .l2_way_state_cache_type_S2 (l2_way_state_cache_type_S2),
    .l2_way_state_subline_S2    (l2_way_state_subline_S2),
    .req_from_owner_S2          (req_from_owner_S2),
    .addr_l2_aligned_S2         (addr_l2_aligned_S2),
    .lsid_S2                    (lsid_S2),
    .dir_addr_S2                (dir_addr),
    .dir_data_in_S2             (dir_data_in),
    .dir_data_mask_in_S2        (dir_data_mask_in),
    .data_addr_S2               (data_addr),
    .data_data_in_S2            (data_data_in),
    .data_data_mask_in_S2       (data_data_mask_in),
    
    .smc_wr_addr_in_S2          (smc_wr_addr_in),
    .smc_data_in_S2             (smc_data_in),
    
    .addr_S3                    (addr_S3),
    .addr_S4                    (addr_S4),
    .data_addr_S4               (data_ecc_addr),
    .l2_evict_S4                (l2_evict_S4),
    .l2_tag_hit_S4              (l2_tag_hit_S4),
    .l2_way_state_mesi_S4       (l2_way_state_mesi_S4),
    .l2_way_state_owner_S4      (l2_way_state_owner_S4),
    .l2_way_state_vd_S4         (l2_way_state_vd_S4),
    .l2_way_state_subline_S4    (l2_way_state_subline_S4),
    .l2_way_state_cache_type_S4 (l2_way_state_cache_type_S4),
    .mshrid_S4                  (mshrid_S4),
    .req_from_owner_S4          (req_from_owner_S4),
    .mshr_miss_lsid_S4          (mshr_miss_lsid_S4),
    .lsid_S4                    (lsid_S4),
    .corr_error_S4              (data_ecc_corr_error),
    .uncorr_error_S4            (data_ecc_uncorr_error),
    .cas_cmp_S4                 (cas_cmp_S4),
    .msg_send_addr_S4           (msg_send_addr),
    .msg_send_dst_chipid_S4     (msg_send_dst_chipid),
    .msg_send_dst_x_S4          (msg_send_dst_x),
    .msg_send_dst_y_S4          (msg_send_dst_y),
    .msg_send_dst_fbits_S4      (msg_send_dst_fbits),
    .msg_send_data_S4           (msg_send_data),
    .mshr_data_in_S4            (mshr_data_in),
    .mshr_data_mask_in_S4       (mshr_data_mask_in),
    
    .smc_rd_addr_in_buf_S4      (smc_rd_addr_in),
    
    .state_wr_addr_S4           (state_wr_addr),
    .state_data_in_S4           (state_data_in),
    .state_data_mask_in_S4      (state_data_mask_in)
);
l2_encoder encoder(
    .msg_dst_chipid             (msg_send_dst_chipid),
    .msg_dst_x                  (msg_send_dst_x),
    .msg_dst_y                  (msg_send_dst_y),
    .msg_dst_fbits              (msg_send_dst_fbits),
    .msg_length                 (msg_send_length),
    .msg_type                   (msg_send_type),
    .msg_mshrid                 (msg_send_mshrid),
    .msg_data_size              (msg_send_data_size),
    .msg_cache_type             (msg_send_cache_type),
    .msg_subline_vector         (msg_send_subline_vector),
    .msg_mesi                   (msg_send_mesi),
    .msg_l2_miss                (msg_send_l2_miss),
    .msg_subline_id             ({2{1'b0}}),
    .msg_last_subline           ({1{1'b0}}),
    .msg_addr                   (msg_send_addr),
    .msg_src_chipid             (my_nodeid[33:20]),
    .msg_src_x                  (my_nodeid[19:12]),
    .msg_src_y                  (my_nodeid[11:4]),
    .msg_src_fbits              (my_nodeid[3:0]),
    .msg_sdid                   ({10{1'b0}}),
    .msg_lsid                   ({6{1'b0}}),
    .msg_header                 (msg_send_header)
);
l2_pipe1_buf_out buf_out(
    .clk                (clk),
    .rst_n              (rst_n),
    .mode_in            (msg_send_mode),
    .valid_in           (msg_send_valid),
    .data_in            ({msg_send_data, msg_send_header}),
    .ready_in           (msg_send_ready),
    .valid_out          (noc_valid_out),
    .data_out           (noc_data_out),
    .ready_out          (noc_ready_out)
);
endmodule
      
 
module l2_pipe2(
    input wire clk,
    input wire rst_n,
    
    input wire csm_en,
    
    
   
    input wire noc_valid_in,
    input wire [64-1:0] noc_data_in,
    output wire noc_ready_in,
    input wire [2-1:0] mshr_state_out,
    input wire [120+2-1:0] mshr_data_out,
    
    input wire broadcast_counter_zero,
    input wire broadcast_counter_max,
    input wire [14-1:0] broadcast_chipid_out,
    input wire [8-1:0] broadcast_x_out,
    input wire [8-1:0] broadcast_y_out,
    
    input wire [15*4+2+4-1:0] state_data_out,
    
    input wire [104-1:0] tag_data_out,
    input wire [64-1:0] dir_data_out,
    output wire mshr_rd_en,
    output wire mshr_wr_state_en,
    output wire mshr_wr_data_en,
    output wire [2-1:0] mshr_state_in,
    output wire [120+2-1:0] mshr_data_in,
    output wire [120+2-1:0] mshr_data_mask_in,
    output wire [3-1:0] mshr_rd_index_in,
    output wire [3-1:0] mshr_wr_index_in,
    output wire mshr_inc_counter_en,
    output wire state_rd_en,
    output wire state_wr_en,
    output wire [8-1:0] state_rd_addr,
    output wire [8-1:0] state_wr_addr,
    output wire [15*4+2+4-1:0] state_data_in,
    output wire [15*4+2+4-1:0] state_data_mask_in,
    output wire tag_clk_en,
    output wire tag_rdw_en,
    output wire [8-1:0] tag_addr,
    output wire [104-1:0] tag_data_in,
    output wire [104-1:0] tag_data_mask_in,
    output wire dir_clk_en,
    output wire dir_rdw_en,
    output wire [8+2-1:0] dir_addr,
    output wire [64-1:0] dir_data_in,
    output wire [64-1:0] dir_data_mask_in,
    output wire data_clk_en,
    output wire data_rdw_en,
    output wire [8+2+2-1:0] data_addr,
    output wire [144-1:0] data_data_in,
    output wire [144-1:0] data_data_mask_in,
    
    output wire [2-1:0] broadcast_counter_op,
    output wire broadcast_counter_op_val,
    output wire smc_wr_en,
    output wire [16-1:0] smc_wr_addr_in,
    output wire [128-1:0] smc_data_in,
    
    output wire valid_S1,
    output wire valid_S2,
    output wire valid_S3,
    output wire [8-1:0] msg_type_S1,
    output wire [8-1:0] msg_type_S2,
    output wire [8-1:0] msg_type_S3,
    output wire [40-1:0] addr_S1,
    output wire [40-1:0] addr_S2,
    output wire [40-1:0] addr_S3,
    output wire active_S1,
    output wire active_S2,
    output wire active_S3
);
wire [8-1:0] msg_type;
wire [8-1:0] msg_length;
wire [8-1:0] msg_mshrid;
wire [3-1:0] msg_data_size;
wire [1-1:0] msg_cache_type;
wire [2-1:0] msg_subline_id;
wire [1-1:0] msg_last_subline;
wire [2-1:0] msg_mesi;
wire [40-1:0] msg_addr;
wire [14-1:0] msg_src_chipid;
wire [8-1:0] msg_src_x;
wire [8-1:0] msg_src_y;
wire [4-1:0] msg_src_fbits;
wire [10-1:0] msg_sdid;
wire [6-1:0] msg_lsid;
wire [8-1:0] mshr_msg_type;
wire [8-1:0] mshr_mshrid;
wire [3-1:0] mshr_data_size;
wire [1-1:0] mshr_cache_type;
wire [40-1:0] mshr_addr;
wire [2-1:0] mshr_way;
wire [1-1:0] mshr_l2_miss;
wire [14-1:0] mshr_src_chipid;
wire [8-1:0] mshr_src_x;
wire [8-1:0] mshr_src_y;
wire [4-1:0] mshr_src_fbits;
wire [10-1:0] mshr_sdid;
wire [6-1:0] mshr_lsid;
wire [6-1:0] mshr_miss_lsid;
wire mshr_smc_miss;
wire mshr_recycled;
wire mshr_inv_fwd_pending;
wire msg_header_valid;
wire [192-1:0] msg_header;
wire msg_header_ready;
wire msg_data_valid;
wire [128-1:0] msg_data;
wire msg_data_ready;
wire stall_S1;
wire msg_from_mshr_S1;
wire is_same_address_S1;
wire stall_S2;
wire stall_before_S2;
wire msg_from_mshr_S2;
wire [3-1:0] data_size_S2;
wire [1-1:0] cache_type_S2;
wire state_owner_en_S2;
wire [2-1:0] state_owner_op_S2;
wire state_subline_en_S2;
wire [2-1:0] state_subline_op_S2;
wire state_di_en_S2;
wire state_vd_en_S2;
wire [2-1:0] state_vd_S2;
wire state_mesi_en_S2;
wire [2-1:0] state_mesi_S2;
wire state_lru_en_S2;
wire [1-1:0] state_lru_op_S2;
wire state_rb_en_S2;
wire dir_clr_en_S2;
wire l2_load_64B_S2;
wire l2_load_32B_S2;
wire [2-1:0] l2_load_data_subline_S2;
wire l2_tag_hit_S2;
wire [2-1:0] l2_way_sel_S2;
wire l2_evict_S2;
wire l2_wb_S2;
wire [6-1:0] l2_way_state_owner_S2;
wire [2-1:0] l2_way_state_mesi_S2;
wire [2-1:0] l2_way_state_vd_S2;
wire [4-1:0] l2_way_state_subline_S2;
wire [1-1:0] l2_way_state_cache_type_S2;
wire addr_l2_aligned_S2;
wire subline_valid_S2;
wire [6-1:0] lsid_S2;
wire stall_S3;
assign msg_type_S1 = msg_type;
l2_pipe2_buf_in buf_in(
    .clk                    (clk),
    .rst_n                  (rst_n),
    .valid_in               (noc_valid_in),
    .data_in                (noc_data_in),
    .ready_in               (noc_ready_in),
    .msg_header_valid_out   (msg_header_valid),
    .msg_header_out         (msg_header),
    .msg_header_ready_out   (msg_header_ready),
    .msg_data_valid_out     (msg_data_valid),
    .msg_data_out           (msg_data),
    .msg_data_ready_out     (msg_data_ready)
);
l2_decoder decoder(
    .msg_header         (msg_header),
    .msg_type           (msg_type),
    .msg_length         (msg_length),
    .msg_mshrid         (msg_mshrid),
    .msg_data_size      (msg_data_size),
    .msg_cache_type     (msg_cache_type),
    .msg_subline_vector (),
    .msg_mesi           (msg_mesi),
    .msg_l2_miss        (),
    .msg_subline_id     (msg_subline_id),
    .msg_last_subline   (msg_last_subline),
    .msg_addr           (msg_addr),
    .msg_src_chipid     (msg_src_chipid),
    .msg_src_x          (msg_src_x),
    .msg_src_y          (msg_src_y),
    .msg_src_fbits      (msg_src_fbits),
    .msg_sdid           (msg_sdid),
    .msg_lsid           (msg_lsid)
);
l2_mshr_decoder mshr_decoder(
    .data_in            (mshr_data_out),
    .addr_out           (mshr_addr),
    .way_out            (mshr_way),
    .mshrid_out         (mshr_mshrid),
    .cache_type_out     (mshr_cache_type), 
    .data_size_out      (mshr_data_size),
    .msg_type_out       (mshr_msg_type),
    .msg_l2_miss_out    (mshr_l2_miss),
    .src_chipid_out     (mshr_src_chipid),
    .src_x_out          (mshr_src_x),
    .src_y_out          (mshr_src_y),
    .src_fbits_out      (mshr_src_fbits),
    .sdid_out           (mshr_sdid),
    .lsid_out           (mshr_lsid),
    .miss_lsid_out      (mshr_miss_lsid),
    
    .smc_miss_out       (mshr_smc_miss),
    
        
    .recycled           (mshr_recycled),
    .inv_fwd_pending    (mshr_inv_fwd_pending)
);
l2_pipe2_ctrl ctrl(
    .clk                        (clk),
    .rst_n                      (rst_n),
    
    .csm_en                     (csm_en),
    
    .msg_header_valid_S1        (msg_header_valid),
    .msg_type_S1                (msg_type),
    .msg_length_S1              (msg_length),
    .msg_data_size_S1           (msg_data_size),
    .msg_cache_type_S1          (msg_cache_type),
    .msg_last_subline_S1        (msg_last_subline),
    .msg_mesi_S1                (msg_mesi),
    .mshr_msg_type_S1           (mshr_msg_type),
    .mshr_l2_miss_S1            (mshr_l2_miss),
    .mshr_data_size_S1          (mshr_data_size),
    .mshr_cache_type_S1         (mshr_cache_type),
     
    .mshr_smc_miss_S1           (mshr_smc_miss),
    
    .mshr_state_out_S1          (mshr_state_out),
    .mshr_inv_fwd_pending_S1    (mshr_inv_fwd_pending),
    .addr_S1                    (addr_S1),
    .is_same_address_S1         (is_same_address_S1),
   
    .l2_tag_hit_S2              (l2_tag_hit_S2),
    .l2_way_sel_S2              (l2_way_sel_S2),
    .l2_wb_S2                   (l2_wb_S2),
    .l2_way_state_owner_S2      (l2_way_state_owner_S2),
    .l2_way_state_mesi_S2       (l2_way_state_mesi_S2),
    .l2_way_state_vd_S2         (l2_way_state_vd_S2),
    .l2_way_state_subline_S2    (l2_way_state_subline_S2),
    .l2_way_state_cache_type_S2 (l2_way_state_cache_type_S2),
    .addr_l2_aligned_S2         (addr_l2_aligned_S2),
    .subline_valid_S2           (subline_valid_S2),
    .msg_data_valid_S2          (msg_data_valid),
    
    .broadcast_counter_zero_S2  (broadcast_counter_zero),
    .broadcast_counter_max_S2   (broadcast_counter_max),
    .broadcast_chipid_out_S2    (broadcast_chipid_out),
    .broadcast_x_out_S2         (broadcast_x_out),
    .broadcast_y_out_S2         (broadcast_y_out),
    
    .lsid_S2                    (lsid_S2),
    .addr_S2                    (addr_S2),
    .addr_S3                    (addr_S3),
    .valid_S1                   (valid_S1),  
    .stall_S1                   (stall_S1), 
    .active_S1                  (active_S1),   
    .msg_from_mshr_S1           (msg_from_mshr_S1), 
    .mshr_rd_en_S1              (mshr_rd_en),
    .msg_header_ready_S1        (msg_header_ready),
    .tag_clk_en_S1              (tag_clk_en),
    .tag_rdw_en_S1              (tag_rdw_en),
    .state_rd_en_S1             (state_rd_en),
    .valid_S2                   (valid_S2),    
    .stall_S2                   (stall_S2), 
    .stall_before_S2            (stall_before_S2), 
    .active_S2                  (active_S2), 
    .msg_from_mshr_S2           (msg_from_mshr_S2),
    .msg_type_S2                (msg_type_S2),
    .data_size_S2               (data_size_S2),
    .cache_type_S2              (cache_type_S2),
    .dir_clk_en_S2              (dir_clk_en),
    .dir_rdw_en_S2              (dir_rdw_en),
    .dir_clr_en_S2              (dir_clr_en_S2),
    .data_clk_en_S2             (data_clk_en),
    .data_rdw_en_S2             (data_rdw_en),
    .state_owner_en_S2          (state_owner_en_S2),
    .state_owner_op_S2          (state_owner_op_S2),
    .state_subline_en_S2        (state_subline_en_S2),
    .state_subline_op_S2        (state_subline_op_S2),   
    .state_di_en_S2             (state_di_en_S2),
    .state_vd_en_S2             (state_vd_en_S2),
    .state_vd_S2                (state_vd_S2),
    .state_mesi_en_S2           (state_mesi_en_S2),
    .state_mesi_S2              (state_mesi_S2),
    .state_lru_en_S2            (state_lru_en_S2),
    .state_lru_op_S2            (state_lru_op_S2),
    .state_rb_en_S2             (state_rb_en_S2),
    .l2_load_64B_S2             (l2_load_64B_S2),
    .l2_load_32B_S2             (l2_load_32B_S2),
    .l2_load_data_subline_S2    (l2_load_data_subline_S2),
    .msg_data_ready_S2          (msg_data_ready),
    
    .smc_wr_en_S2               (smc_wr_en),
    .broadcast_counter_op_S2    (broadcast_counter_op),
    .broadcast_counter_op_val_S2(broadcast_counter_op_val),
    
    .valid_S3                   (valid_S3),    
    .stall_S3                   (stall_S3), 
    .active_S3                  (active_S3),   
    .msg_type_S3                (msg_type_S3),
    .mshr_wr_state_en_S3        (mshr_wr_state_en),
    .mshr_wr_data_en_S3         (mshr_wr_data_en),
    .mshr_state_in_S3           (mshr_state_in),
    .mshr_inc_counter_en_S3     (mshr_inc_counter_en),
    .state_wr_en_S3             (state_wr_en)
);
l2_pipe2_dpath dpath(
    .clk                        (clk),
    .rst_n                      (rst_n),
    .mshr_addr_S1               (mshr_addr),
    .mshr_mshrid_S1             (mshr_mshrid),
    .mshr_way_S1                (mshr_way),
    .mshr_src_chipid_S1         (mshr_src_chipid),
    .mshr_src_x_S1              (mshr_src_x),
    .mshr_src_y_S1              (mshr_src_y),
    .mshr_src_fbits_S1          (mshr_src_fbits),
    .mshr_sdid_S1               (mshr_sdid),
    .mshr_lsid_S1               (mshr_lsid),
    .mshr_miss_lsid_S1          (mshr_miss_lsid),
    .msg_addr_S1                (msg_addr),
    .msg_type_S1                (msg_type),
    .msg_subline_id_S1          (msg_subline_id),
    .msg_mshrid_S1              (msg_mshrid),
    .msg_src_chipid_S1          (msg_src_chipid),
    .msg_src_x_S1               (msg_src_x),
    .msg_src_y_S1               (msg_src_y),
    .msg_src_fbits_S1           (msg_src_fbits),
    .msg_sdid_S1                (msg_sdid),
    .msg_lsid_S1                (msg_lsid),
    .valid_S1                   (valid_S1),
    .stall_S1                   (stall_S1),
    .msg_from_mshr_S1           (msg_from_mshr_S1), 
    .state_data_S2              (state_data_out),
    .tag_data_S2                (tag_data_out),
    .msg_data_S2                (msg_data),
    .msg_from_mshr_S2           (msg_from_mshr_S2),
    .msg_type_S2                (msg_type_S2),
    .data_size_S2               (data_size_S2),
    .cache_type_S2              (cache_type_S2),
    .state_owner_en_S2          (state_owner_en_S2),
    .state_owner_op_S2          (state_owner_op_S2), 
    .state_subline_en_S2        (state_subline_en_S2),
    .state_subline_op_S2        (state_subline_op_S2),
    .state_di_en_S2             (state_di_en_S2),
    .state_vd_en_S2             (state_vd_en_S2),
    .state_vd_S2                (state_vd_S2),
    .state_mesi_en_S2           (state_mesi_en_S2),
    .state_mesi_S2              (state_mesi_S2),
    .state_lru_en_S2            (state_lru_en_S2),
    .state_lru_op_S2            (state_lru_op_S2),
    .state_rb_en_S2             (state_rb_en_S2),
    .dir_clr_en_S2              (dir_clr_en_S2),
    .l2_load_64B_S2             (l2_load_64B_S2),
    .l2_load_32B_S2             (l2_load_32B_S2),
    .l2_load_data_subline_S2    (l2_load_data_subline_S2),
    .valid_S2                   (valid_S2),
    .stall_S2                   (stall_S2),
    .stall_before_S2            (stall_before_S2), 
    .valid_S3                   (valid_S3),
    .stall_S3                   (stall_S3),
    .addr_S1                    (addr_S1),
    .mshr_rd_index_S1           (mshr_rd_index_in),
    .tag_addr_S1                (tag_addr),
    .state_rd_addr_S1           (state_rd_addr),
    .tag_data_in_S1             (tag_data_in),  
    .tag_data_mask_in_S1        (tag_data_mask_in),
    .is_same_address_S1         (is_same_address_S1),
    .addr_S2                    (addr_S2),
    .l2_tag_hit_S2              (l2_tag_hit_S2),
    .l2_way_sel_S2              (l2_way_sel_S2),
    .l2_wb_S2                   (l2_wb_S2),
    .l2_way_state_owner_S2      (l2_way_state_owner_S2),
    .l2_way_state_mesi_S2       (l2_way_state_mesi_S2),
    .l2_way_state_vd_S2         (l2_way_state_vd_S2),    
    .l2_way_state_subline_S2    (l2_way_state_subline_S2),
    .l2_way_state_cache_type_S2 (l2_way_state_cache_type_S2),
    .addr_l2_aligned_S2         (addr_l2_aligned_S2),
    .subline_valid_S2           (subline_valid_S2),
    .lsid_S2                    (lsid_S2),
    .dir_addr_S2                (dir_addr),
    .dir_data_in_S2             (dir_data_in),
    .dir_data_mask_in_S2        (dir_data_mask_in),
    .data_addr_S2               (data_addr),
    .data_data_in_S2            (data_data_in),
    .data_data_mask_in_S2       (data_data_mask_in),
    
    .smc_wr_addr_in_S2          (smc_wr_addr_in),
    .smc_data_in_S2             (smc_data_in),
    
    .addr_S3                    (addr_S3),
    .mshr_wr_index_S3           (mshr_wr_index_in),
    .mshr_data_in_S3            (mshr_data_in),
    .mshr_data_mask_in_S3       (mshr_data_mask_in),
    .state_wr_addr_S3           (state_wr_addr),
    .state_data_in_S3           (state_data_in),
    .state_data_mask_in_S3      (state_data_mask_in)
);
endmodule
      
 
module l2_smc_wrap(
    input wire clk,
    input wire rst_n,
    input wire pipe_sel,
    input wire rd_en,
    input wire rd_diag_en,
    input wire flush_en,
    input wire [2-1:0] addr_op,
    input wire [16-1:0] rd_addr_in,
    input wire wr_en1,
    input wire [16-1:0] wr_addr_in1,
    input wire [128-1:0] data_in1,
    input wire wr_diag_en1,
    input wire wr_en2,
    input wire [16-1:0] wr_addr_in2,
    input wire [128-1:0] data_in2,
    input wire wr_diag_en2,
    output wire hit,
    output wire [30-1:0] data_out,
    output wire [4-1:0] valid_out,
    output wire [14-1:0] tag_out
);
reg wr_en;
reg [16-1:0] wr_addr_in;
reg [128-1:0] data_in;
reg wr_diag_en;
always @ *
begin
    if (pipe_sel)
    begin
        wr_en = wr_en2;
        wr_addr_in = wr_addr_in2;
        data_in = data_in2;
        wr_diag_en = wr_diag_en2;
    end
    else
    begin
        wr_en = wr_en1;
        wr_addr_in = wr_addr_in1;
        data_in = data_in1;
        wr_diag_en = wr_diag_en1;
    end
end
l2_smc l2_smc(
    .clk            (clk),
    .rst_n          (rst_n),
    .rd_en          (rd_en),
    .wr_en          (wr_en),
    .rd_diag_en     (rd_diag_en),
    .wr_diag_en     (wr_diag_en),
    .flush_en       (flush_en),
    .addr_op        (addr_op),
    .rd_addr_in     (rd_addr_in),
    .wr_addr_in     (wr_addr_in),
    .data_in        (data_in),
    .hit            (hit),
    .data_out       (data_out),
    .valid_out      (valid_out),
    .tag_out        (tag_out)
);
endmodule
      
 
module l2_state_wrap(
    input wire clk,
    input wire rst_n,
    input wire pipe_rd_sel,
    input wire pipe_wr_sel,
    input wire pdout_en,
    input wire deepsleep,
    input wire rd_en1,
    input wire wr_en1,
    input wire [8-1:0] rd_addr1,
    input wire [8-1:0] wr_addr1,
    input wire [15*4+2+4-1:0] data_in1,
    input wire [15*4+2+4-1:0] data_mask_in1,
    input wire rd_en2,
    input wire wr_en2,
    input wire [8-1:0] rd_addr2,
    input wire [8-1:0] wr_addr2,
    input wire [15*4+2+4-1:0] data_in2,
    input wire [15*4+2+4-1:0] data_mask_in2,
    output wire [15*4+2+4-1:0] data_out,
    output wire [15*4+2+4-1:0] pdata_out,
    
    output wire [4-1:0] srams_rtap_data,
    input wire  [4-1:0] rtap_srams_bist_command,
    input wire  [4-1:0] rtap_srams_bist_data
);
reg rd_en;
reg wr_en;
reg [8-1:0] rd_addr;
reg [8-1:0] wr_addr;
reg [15*4+2+4-1:0] data_in;
reg [15*4+2+4-1:0] data_mask_in;
always @ *
begin
    if (pipe_rd_sel)
    begin
        rd_en = rd_en2;
        rd_addr = rd_addr2;
    end
    else
    begin
        rd_en = rd_en1;
        rd_addr = rd_addr1;
    end
end
always @ *
begin
    if (pipe_wr_sel)
    begin
        wr_en = wr_en2;
        wr_addr = wr_addr2;
        data_in = data_in2;
        data_mask_in = data_mask_in2;
     end
    else
    begin
        wr_en = wr_en1;
        wr_addr = wr_addr1;
        data_in = data_in1;
        data_mask_in = data_mask_in1;
    end
end
l2_state l2_state(
    .clk            (clk),
    .rst_n          (rst_n),
    .rd_en          (rd_en),
    .wr_en          (wr_en),
    .pdout_en       (pdout_en),
    .deepsleep      (deepsleep),
    .rd_addr        (rd_addr),
    .wr_addr        (wr_addr),
    .data_in        (data_in),
    .data_mask_in   (data_mask_in),
    .data_out       (data_out),
    .pdata_out      (pdata_out),
    
    .srams_rtap_data (srams_rtap_data),
    .rtap_srams_bist_command (rtap_srams_bist_command),
    .rtap_srams_bist_data (rtap_srams_bist_data)
);
endmodule
      
 
module l2_tag(
    input wire clk,
    input wire rst_n,
    input wire clk_en,
    
    input wire rdw_en,
    input wire pdout_en,
    input wire deepsleep,
    input wire [8-1:0] addr,
    input wire [104-1:0] data_in,
    input wire [104-1:0] data_mask_in,
    output wire [104-1:0] data_out,
    output wire [104-1:0] pdata_out,
    
    output wire [4-1:0] srams_rtap_data,
    input wire  [4-1:0] rtap_srams_bist_command,
    input wire  [4-1:0] rtap_srams_bist_data
);
sram_l2_tag l2_tag_array(
    .MEMCLK     (clk),
    .RESET_N(rst_n),
    .CE         (clk_en),
    .A          (addr),
    .DIN        (data_in),
    .RDWEN      (rdw_en),
    .BW         (data_mask_in),
    .DOUT       (data_out),
    .BIST_COMMAND(rtap_srams_bist_command),
    .BIST_DIN(rtap_srams_bist_data),
    .BIST_DOUT(srams_rtap_data),
    .SRAMID(8'd16)
);
endmodule
      
 
module l2_tag_wrap(
    input wire clk,
    input wire rst_n,
    input wire clk_en1,
    input wire clk_en2,
    input wire rdw_en1,
    input wire rdw_en2,
    input wire pdout_en,
    input wire deepsleep,
    input wire pipe_sel,
    input wire [8-1:0] addr1,
    input wire [104-1:0] data_in1,
    input wire [104-1:0] data_mask_in1,
    input wire [8-1:0] addr2,
    input wire [104-1:0] data_in2,
    input wire [104-1:0] data_mask_in2,
    output wire [104-1:0] data_out,
    output wire [104-1:0] pdata_out,
    
    output wire [4-1:0] srams_rtap_data,
    input wire  [4-1:0] rtap_srams_bist_command,
    input wire  [4-1:0] rtap_srams_bist_data
);
reg clk_en;
reg rdw_en;
reg [8-1:0] addr;
reg [104-1:0] data_in;
reg [104-1:0] data_mask_in;
always @ *
begin
    if (pipe_sel)
    begin
        clk_en = clk_en2;
        rdw_en = rdw_en2;
        addr = addr2;
        data_in = data_in2;
        data_mask_in = data_mask_in2;
    end
    else
    begin
        clk_en = clk_en1;
        rdw_en = rdw_en1;
        addr = addr1;
        data_in = data_in1;
        data_mask_in = data_mask_in1;
    end
end
l2_tag l2_tag(
    .clk            (clk),
    .rst_n          (rst_n),
    .clk_en         (clk_en),
    .rdw_en         (rdw_en),
    .pdout_en       (pdout_en),
    .deepsleep      (deepsleep),
    .addr           (addr),
    .data_in        (data_in),
    .data_mask_in   (data_mask_in),
    .data_out       (data_out),
    .pdata_out      (pdata_out),
    
    .srams_rtap_data (srams_rtap_data),
    .rtap_srams_bist_command (rtap_srams_bist_command),
    .rtap_srams_bist_data (rtap_srams_bist_data)
);
endmodule
      
 
module l2_data_ecc ( 
   input  [64-1:0]      din,
   input  [8-1:0]	 parity,
   output [64-1:0]      dout,
   output                                    corr_error,
   output                                    uncorr_error
);
   
wire [64-1:0] 	err_bit_pos;
wire [8-2:0]    cflag;
wire 	                                pflag;
assign cflag[0] = parity[0]  ^ din[0] ^ din[1] ^ din[3] ^ din[4] ^ din[6] ^ din[8] ^ din[10] ^ din[11] ^ din[13] ^ din[15] ^ din[17] ^ din[19] ^ din[21] ^ din[23] ^ din[25] ^ din[26] ^ din[28] ^ din[30] ^ din[32] ^ din[34] ^ din[36] ^ din[38] ^ din[40] ^ din[42] ^ din[44] ^ din[46] ^ din[48] ^ din[50] ^ din[52] ^ din[54] ^ din[56] ^ din[57] ^ din[59] ^ din[61] ^ din[63] ;
assign cflag[1] = parity[1]  ^ din[0] ^ din[2] ^ din[3] ^ din[5] ^ din[6] ^ din[9] ^ din[10] ^ din[12] ^ din[13] ^ din[16] ^ din[17] ^ din[20] ^ din[21] ^ din[24] ^ din[25] ^ din[27] ^ din[28] ^ din[31] ^ din[32] ^ din[35] ^ din[36] ^ din[39] ^ din[40] ^ din[43] ^ din[44] ^ din[47] ^ din[48] ^ din[51] ^ din[52] ^ din[55] ^ din[56] ^ din[58] ^ din[59] ^ din[62] ^ din[63] ;
assign cflag[2] = parity[2]  ^ din[1] ^ din[2] ^ din[3] ^ din[7] ^ din[8] ^ din[9] ^ din[10] ^ din[14] ^ din[15] ^ din[16] ^ din[17] ^ din[22] ^ din[23] ^ din[24] ^ din[25] ^ din[29] ^ din[30] ^ din[31] ^ din[32] ^ din[37] ^ din[38] ^ din[39] ^ din[40] ^ din[45] ^ din[46] ^ din[47] ^ din[48] ^ din[53] ^ din[54] ^ din[55] ^ din[56] ^ din[60] ^ din[61] ^ din[62] ^ din[63] ;
assign cflag[3] = parity[3]  ^ din[4] ^ din[5] ^ din[6] ^ din[7] ^ din[8] ^ din[9] ^ din[10] ^ din[18] ^ din[19] ^ din[20] ^ din[21] ^ din[22] ^ din[23] ^ din[24] ^ din[25] ^ din[33] ^ din[34] ^ din[35] ^ din[36] ^ din[37] ^ din[38] ^ din[39] ^ din[40] ^ din[49] ^ din[50] ^ din[51] ^ din[52] ^ din[53] ^ din[54] ^ din[55] ^ din[56] ;
assign cflag[4] = parity[4]  ^ din[11] ^ din[12] ^ din[13] ^ din[14] ^ din[15] ^ din[16] ^ din[17] ^ din[18] ^ din[19] ^ din[20] ^ din[21] ^ din[22] ^ din[23] ^ din[24] ^ din[25] ^ din[41] ^ din[42] ^ din[43] ^ din[44] ^ din[45] ^ din[46] ^ din[47] ^ din[48] ^ din[49] ^ din[50] ^ din[51] ^ din[52] ^ din[53] ^ din[54] ^ din[55] ^ din[56] ;
assign cflag[5] = parity[5]  ^ din[26] ^ din[27] ^ din[28] ^ din[29] ^ din[30] ^ din[31] ^ din[32] ^ din[33] ^ din[34] ^ din[35] ^ din[36] ^ din[37] ^ din[38] ^ din[39] ^ din[40] ^ din[41] ^ din[42] ^ din[43] ^ din[44] ^ din[45] ^ din[46] ^ din[47] ^ din[48] ^ din[49] ^ din[50] ^ din[51] ^ din[52] ^ din[53] ^ din[54] ^ din[55] ^ din[56] ;
assign cflag[6] = parity[6]  ^ din[57] ^ din[58] ^ din[59] ^ din[60] ^ din[61] ^ din[62] ^ din[63] ;
assign pflag = cflag[0]
 ^ parity[1]  ^ parity[2]  ^ parity[3]  ^ parity[4]  ^ parity[5]  ^ parity[6] 
^ din[2] ^ din[5] ^ din[7] ^ din[9] ^ din[12] ^ din[14] ^ din[16] ^ din[18] ^ din[20] ^ din[22] ^ din[24] ^ din[27] ^ din[29] ^ din[31] ^ din[33] ^ din[35] ^ din[37] ^ din[39] ^ din[41] ^ din[43] ^ din[45] ^ din[47] ^ din[49] ^ din[51] ^ din[53] ^ din[55] ^ din[58] ^ din[60] ^ din[62] ;
assign err_bit_pos[0] =  (cflag[0]) & (cflag[1]) & (~cflag[2]) & (~cflag[3]) & (~cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[1] =  (cflag[0]) & (~cflag[1]) & (cflag[2]) & (~cflag[3]) & (~cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[2] =  (~cflag[0]) & (cflag[1]) & (cflag[2]) & (~cflag[3]) & (~cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[3] =  (cflag[0]) & (cflag[1]) & (cflag[2]) & (~cflag[3]) & (~cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[4] =  (cflag[0]) & (~cflag[1]) & (~cflag[2]) & (cflag[3]) & (~cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[5] =  (~cflag[0]) & (cflag[1]) & (~cflag[2]) & (cflag[3]) & (~cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[6] =  (cflag[0]) & (cflag[1]) & (~cflag[2]) & (cflag[3]) & (~cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[7] =  (~cflag[0]) & (~cflag[1]) & (cflag[2]) & (cflag[3]) & (~cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[8] =  (cflag[0]) & (~cflag[1]) & (cflag[2]) & (cflag[3]) & (~cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[9] =  (~cflag[0]) & (cflag[1]) & (cflag[2]) & (cflag[3]) & (~cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[10] =  (cflag[0]) & (cflag[1]) & (cflag[2]) & (cflag[3]) & (~cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[11] =  (cflag[0]) & (~cflag[1]) & (~cflag[2]) & (~cflag[3]) & (cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[12] =  (~cflag[0]) & (cflag[1]) & (~cflag[2]) & (~cflag[3]) & (cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[13] =  (cflag[0]) & (cflag[1]) & (~cflag[2]) & (~cflag[3]) & (cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[14] =  (~cflag[0]) & (~cflag[1]) & (cflag[2]) & (~cflag[3]) & (cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[15] =  (cflag[0]) & (~cflag[1]) & (cflag[2]) & (~cflag[3]) & (cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[16] =  (~cflag[0]) & (cflag[1]) & (cflag[2]) & (~cflag[3]) & (cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[17] =  (cflag[0]) & (cflag[1]) & (cflag[2]) & (~cflag[3]) & (cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[18] =  (~cflag[0]) & (~cflag[1]) & (~cflag[2]) & (cflag[3]) & (cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[19] =  (cflag[0]) & (~cflag[1]) & (~cflag[2]) & (cflag[3]) & (cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[20] =  (~cflag[0]) & (cflag[1]) & (~cflag[2]) & (cflag[3]) & (cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[21] =  (cflag[0]) & (cflag[1]) & (~cflag[2]) & (cflag[3]) & (cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[22] =  (~cflag[0]) & (~cflag[1]) & (cflag[2]) & (cflag[3]) & (cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[23] =  (cflag[0]) & (~cflag[1]) & (cflag[2]) & (cflag[3]) & (cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[24] =  (~cflag[0]) & (cflag[1]) & (cflag[2]) & (cflag[3]) & (cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[25] =  (cflag[0]) & (cflag[1]) & (cflag[2]) & (cflag[3]) & (cflag[4]) & (~cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[26] =  (cflag[0]) & (~cflag[1]) & (~cflag[2]) & (~cflag[3]) & (~cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[27] =  (~cflag[0]) & (cflag[1]) & (~cflag[2]) & (~cflag[3]) & (~cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[28] =  (cflag[0]) & (cflag[1]) & (~cflag[2]) & (~cflag[3]) & (~cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[29] =  (~cflag[0]) & (~cflag[1]) & (cflag[2]) & (~cflag[3]) & (~cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[30] =  (cflag[0]) & (~cflag[1]) & (cflag[2]) & (~cflag[3]) & (~cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[31] =  (~cflag[0]) & (cflag[1]) & (cflag[2]) & (~cflag[3]) & (~cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[32] =  (cflag[0]) & (cflag[1]) & (cflag[2]) & (~cflag[3]) & (~cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[33] =  (~cflag[0]) & (~cflag[1]) & (~cflag[2]) & (cflag[3]) & (~cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[34] =  (cflag[0]) & (~cflag[1]) & (~cflag[2]) & (cflag[3]) & (~cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[35] =  (~cflag[0]) & (cflag[1]) & (~cflag[2]) & (cflag[3]) & (~cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[36] =  (cflag[0]) & (cflag[1]) & (~cflag[2]) & (cflag[3]) & (~cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[37] =  (~cflag[0]) & (~cflag[1]) & (cflag[2]) & (cflag[3]) & (~cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[38] =  (cflag[0]) & (~cflag[1]) & (cflag[2]) & (cflag[3]) & (~cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[39] =  (~cflag[0]) & (cflag[1]) & (cflag[2]) & (cflag[3]) & (~cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[40] =  (cflag[0]) & (cflag[1]) & (cflag[2]) & (cflag[3]) & (~cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[41] =  (~cflag[0]) & (~cflag[1]) & (~cflag[2]) & (~cflag[3]) & (cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[42] =  (cflag[0]) & (~cflag[1]) & (~cflag[2]) & (~cflag[3]) & (cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[43] =  (~cflag[0]) & (cflag[1]) & (~cflag[2]) & (~cflag[3]) & (cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[44] =  (cflag[0]) & (cflag[1]) & (~cflag[2]) & (~cflag[3]) & (cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[45] =  (~cflag[0]) & (~cflag[1]) & (cflag[2]) & (~cflag[3]) & (cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[46] =  (cflag[0]) & (~cflag[1]) & (cflag[2]) & (~cflag[3]) & (cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[47] =  (~cflag[0]) & (cflag[1]) & (cflag[2]) & (~cflag[3]) & (cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[48] =  (cflag[0]) & (cflag[1]) & (cflag[2]) & (~cflag[3]) & (cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[49] =  (~cflag[0]) & (~cflag[1]) & (~cflag[2]) & (cflag[3]) & (cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[50] =  (cflag[0]) & (~cflag[1]) & (~cflag[2]) & (cflag[3]) & (cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[51] =  (~cflag[0]) & (cflag[1]) & (~cflag[2]) & (cflag[3]) & (cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[52] =  (cflag[0]) & (cflag[1]) & (~cflag[2]) & (cflag[3]) & (cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[53] =  (~cflag[0]) & (~cflag[1]) & (cflag[2]) & (cflag[3]) & (cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[54] =  (cflag[0]) & (~cflag[1]) & (cflag[2]) & (cflag[3]) & (cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[55] =  (~cflag[0]) & (cflag[1]) & (cflag[2]) & (cflag[3]) & (cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[56] =  (cflag[0]) & (cflag[1]) & (cflag[2]) & (cflag[3]) & (cflag[4]) & (cflag[5]) & (~cflag[6]) ;
assign err_bit_pos[57] =  (cflag[0]) & (~cflag[1]) & (~cflag[2]) & (~cflag[3]) & (~cflag[4]) & (~cflag[5]) & (cflag[6]) ;
assign err_bit_pos[58] =  (~cflag[0]) & (cflag[1]) & (~cflag[2]) & (~cflag[3]) & (~cflag[4]) & (~cflag[5]) & (cflag[6]) ;
assign err_bit_pos[59] =  (cflag[0]) & (cflag[1]) & (~cflag[2]) & (~cflag[3]) & (~cflag[4]) & (~cflag[5]) & (cflag[6]) ;
assign err_bit_pos[60] =  (~cflag[0]) & (~cflag[1]) & (cflag[2]) & (~cflag[3]) & (~cflag[4]) & (~cflag[5]) & (cflag[6]) ;
assign err_bit_pos[61] =  (cflag[0]) & (~cflag[1]) & (cflag[2]) & (~cflag[3]) & (~cflag[4]) & (~cflag[5]) & (cflag[6]) ;
assign err_bit_pos[62] =  (~cflag[0]) & (cflag[1]) & (cflag[2]) & (~cflag[3]) & (~cflag[4]) & (~cflag[5]) & (cflag[6]) ;
assign err_bit_pos[63] =  (cflag[0]) & (cflag[1]) & (cflag[2]) & (~cflag[3]) & (~cflag[4]) & (~cflag[5]) & (cflag[6]) ;
assign dout = din ^ err_bit_pos;
assign corr_error = pflag;
assign uncorr_error = |(cflag[8-2:0]) & ~pflag;
endmodule
      
 
module l2_data_pgen ( 
   input    [64-1:0]   din,
   output   [8-1:0] parity
);
assign parity[0] =  din[0] ^ din[1] ^ din[3] ^ din[4] ^ din[6] ^ din[8] ^ din[10] ^ din[11] ^ din[13] ^ din[15] ^ din[17] ^ din[19] ^ din[21] ^ din[23] ^ din[25] ^ din[26] ^ din[28] ^ din[30] ^ din[32] ^ din[34] ^ din[36] ^ din[38] ^ din[40] ^ din[42] ^ din[44] ^ din[46] ^ din[48] ^ din[50] ^ din[52] ^ din[54] ^ din[56] ^ din[57] ^ din[59] ^ din[61] ^ din[63] ;
assign parity[1] =  din[0] ^ din[2] ^ din[3] ^ din[5] ^ din[6] ^ din[9] ^ din[10] ^ din[12] ^ din[13] ^ din[16] ^ din[17] ^ din[20] ^ din[21] ^ din[24] ^ din[25] ^ din[27] ^ din[28] ^ din[31] ^ din[32] ^ din[35] ^ din[36] ^ din[39] ^ din[40] ^ din[43] ^ din[44] ^ din[47] ^ din[48] ^ din[51] ^ din[52] ^ din[55] ^ din[56] ^ din[58] ^ din[59] ^ din[62] ^ din[63] ;
assign parity[2] =  din[1] ^ din[2] ^ din[3] ^ din[7] ^ din[8] ^ din[9] ^ din[10] ^ din[14] ^ din[15] ^ din[16] ^ din[17] ^ din[22] ^ din[23] ^ din[24] ^ din[25] ^ din[29] ^ din[30] ^ din[31] ^ din[32] ^ din[37] ^ din[38] ^ din[39] ^ din[40] ^ din[45] ^ din[46] ^ din[47] ^ din[48] ^ din[53] ^ din[54] ^ din[55] ^ din[56] ^ din[60] ^ din[61] ^ din[62] ^ din[63] ;
assign parity[3] =  din[4] ^ din[5] ^ din[6] ^ din[7] ^ din[8] ^ din[9] ^ din[10] ^ din[18] ^ din[19] ^ din[20] ^ din[21] ^ din[22] ^ din[23] ^ din[24] ^ din[25] ^ din[33] ^ din[34] ^ din[35] ^ din[36] ^ din[37] ^ din[38] ^ din[39] ^ din[40] ^ din[49] ^ din[50] ^ din[51] ^ din[52] ^ din[53] ^ din[54] ^ din[55] ^ din[56] ;
assign parity[4] =  din[11] ^ din[12] ^ din[13] ^ din[14] ^ din[15] ^ din[16] ^ din[17] ^ din[18] ^ din[19] ^ din[20] ^ din[21] ^ din[22] ^ din[23] ^ din[24] ^ din[25] ^ din[41] ^ din[42] ^ din[43] ^ din[44] ^ din[45] ^ din[46] ^ din[47] ^ din[48] ^ din[49] ^ din[50] ^ din[51] ^ din[52] ^ din[53] ^ din[54] ^ din[55] ^ din[56] ;
assign parity[5] =  din[26] ^ din[27] ^ din[28] ^ din[29] ^ din[30] ^ din[31] ^ din[32] ^ din[33] ^ din[34] ^ din[35] ^ din[36] ^ din[37] ^ din[38] ^ din[39] ^ din[40] ^ din[41] ^ din[42] ^ din[43] ^ din[44] ^ din[45] ^ din[46] ^ din[47] ^ din[48] ^ din[49] ^ din[50] ^ din[51] ^ din[52] ^ din[53] ^ din[54] ^ din[55] ^ din[56] ;
assign parity[6] =  din[57] ^ din[58] ^ din[59] ^ din[60] ^ din[61] ^ din[62] ^ din[63] ;
assign parity[7] =  din[0] ^ din[1] ^ din[2] ^ din[4] ^ din[5] ^ din[7] ^ din[10] ^ din[11] ^ din[12] ^ din[14] ^ din[17] ^ din[18] ^ din[21] ^ din[23] ^ din[24] ^ din[26] ^ din[27] ^ din[29] ^ din[32] ^ din[33] ^ din[36] ^ din[38] ^ din[39] ^ din[41] ^ din[44] ^ din[46] ^ din[47] ^ din[50] ^ din[51] ^ din[53] ^ din[56] ^ din[57] ^ din[58] ^ din[60] ^ din[63] ;
endmodule 
      
 
module l2_mshr(
    input wire clk,
    input wire rst_n,
    
    input wire rd_en,
    
    input wire cam_en,
    
    input wire wr_state_en,
    
    input wire wr_data_en,
    
    input wire pending_ready,
    
    input wire inc_counter_en,
    
    input wire [2-1:0] state_in,
    
    input wire [120+2-1:0] data_in,
    input wire [120+2-1:0] data_mask_in,
    
    input wire [3-1:0] rd_index_in,
    
    input wire [3-1:0] inv_counter_rd_index_in,
    
    input wire [3-1:0] wr_index_in,
    
    input wire [8-1:0] addr_in,
    output reg hit,
    output reg [3-1:0] hit_index,
    
    
    output reg [2-1:0] state_out,
    output reg [120+2-1:0] data_out,
    output reg [6-1:0] inv_counter_out,
    
    output reg [3:0] empty_slots,
    output reg pending,
    output reg [3-1:0] pending_index,
    output reg [3-1:0] empty_index
);
reg [2-1:0] state_mem_f [8-1:0];
reg [120+2-1:0] data_mem_f [8-1:0];
reg [6-1:0] counter_mem_f [8-1:0];
reg [3-1:0] wbg_counter_f;
reg [3-1:0] wbg_counter_next;
always @ *
begin
    empty_slots = 0;
    if (state_mem_f[0] == 2'd0)
    begin
        empty_slots = empty_slots + 1;
    end
    if (state_mem_f[1] == 2'd0)
    begin
        empty_slots = empty_slots + 1;
    end
    if (state_mem_f[2] == 2'd0)
    begin
        empty_slots = empty_slots + 1;
    end
    if (state_mem_f[3] == 2'd0)
    begin
        empty_slots = empty_slots + 1;
    end
    if (state_mem_f[4] == 2'd0)
    begin
        empty_slots = empty_slots + 1;
    end
    if (state_mem_f[5] == 2'd0)
    begin
        empty_slots = empty_slots + 1;
    end
    if (state_mem_f[6] == 2'd0)
    begin
        empty_slots = empty_slots + 1;
    end
    if (state_mem_f[7] == 2'd0)
    begin
        empty_slots = empty_slots + 1;
    end
end
always @ *
begin
    if (state_mem_f[0] == 2'd2)
    begin
        pending = 1'b1;
        pending_index = 3'd0;
    end
    else if (state_mem_f[1] == 2'd2)
    begin
        pending = 1'b1;
        pending_index = 3'd1;
    end
    else if (state_mem_f[2] == 2'd2)
    begin
        pending = 1'b1;
        pending_index = 3'd2;
    end
    else if (state_mem_f[3] == 2'd2)
    begin
        pending = 1'b1;
        pending_index = 3'd3;
    end
    else if (state_mem_f[4] == 2'd2)
    begin
        pending = 1'b1;
        pending_index = 3'd4;
    end
    else if (state_mem_f[5] == 2'd2)
    begin
        pending = 1'b1;
        pending_index = 3'd5;
    end
    else if (state_mem_f[6] == 2'd2)
    begin
        pending = 1'b1;
        pending_index = 3'd6;
    end
    else if (state_mem_f[7] == 2'd2)
    begin
        pending = 1'b1;
        pending_index = 3'd7;
    end
    else
    begin
        pending = 1'b0;
        pending_index = 3'd0;
    end
end
always @ *
begin
    if (state_mem_f[0] == 2'd0)
    begin
        empty_index = 3'd0;
    end
    else if (state_mem_f[1] == 2'd0)
    begin
        empty_index = 3'd1;
    end
    else if (state_mem_f[2] == 2'd0)
    begin
        empty_index = 3'd2;
    end
    else if (state_mem_f[3] == 2'd0)
    begin
        empty_index = 3'd3;
    end
    else if (state_mem_f[4] == 2'd0)
    begin
        empty_index = 3'd4;
    end
    else if (state_mem_f[5] == 2'd0)
    begin
        empty_index = 3'd5;
    end
    else if (state_mem_f[6] == 2'd0)
    begin
        empty_index = 3'd6;
    end
    else if (state_mem_f[7] == 2'd0)
    begin
        empty_index = 3'd7;
    end
    else
    begin
        empty_index = 3'd0;
    end
end
always @ *
begin
    if (rd_en)
    begin
        state_out = state_mem_f[rd_index_in];
        data_out = data_mem_f[rd_index_in];
    end
    else if (cam_en && hit)
    begin
        state_out = state_mem_f[hit_index];
        data_out = data_mem_f[hit_index];
    end
    else if (pending)
    begin
        state_out = state_mem_f[pending_index];
        data_out = data_mem_f[pending_index];
    end
    else
    begin
        state_out = 2'd0;
        data_out = 0;
    end
end
always @ *
begin
    inv_counter_out = counter_mem_f[inv_counter_rd_index_in];
end
always @ *
begin
    if(cam_en)
    begin
        if ((data_mem_f[0][6+8-1:6] == addr_in) && (state_mem_f[0] != 2'd0))
        begin
            hit = 1'b1;
            hit_index = 3'd0;
        end
        else if ((data_mem_f[1][6+8-1:6] == addr_in) && (state_mem_f[1] != 2'd0))
        begin
            hit = 1'b1;
            hit_index = 3'd1;
        end
        else if ((data_mem_f[2][6+8-1:6] == addr_in) && (state_mem_f[2] != 2'd0))
        begin
            hit = 1'b1;
            hit_index = 3'd2;
        end
        else if ((data_mem_f[3][6+8-1:6] == addr_in) && (state_mem_f[3] != 2'd0))
        begin
            hit = 1'b1;
            hit_index = 3'd3;
        end
        else if ((data_mem_f[4][6+8-1:6] == addr_in) && (state_mem_f[4] != 2'd0))
        begin
            hit = 1'b1;
            hit_index = 3'd4;
        end
        else if ((data_mem_f[5][6+8-1:6] == addr_in) && (state_mem_f[5] != 2'd0))
        begin
            hit = 1'b1;
            hit_index = 3'd5;
        end
        else if ((data_mem_f[6][6+8-1:6] == addr_in) && (state_mem_f[6] != 2'd0))
        begin
            hit = 1'b1;
            hit_index = 3'd6;
        end
        else if ((data_mem_f[7][6+8-1:6] == addr_in) && (state_mem_f[7] != 2'd0))
        begin
            hit = 1'b1;
            hit_index = 3'd7;
        end
        else
        begin
            hit = 1'b0;
            hit_index = 3'd0;
        end
    end
    else
    begin
        hit = 1'b0;
        hit_index = 3'd0;
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        state_mem_f[0] <= 2'd0;
        state_mem_f[1] <= 2'd0;
        state_mem_f[2] <= 2'd0;
        state_mem_f[3] <= 2'd0;
        state_mem_f[4] <= 2'd0;
        state_mem_f[5] <= 2'd0;
        state_mem_f[6] <= 2'd0;
        state_mem_f[7] <= 2'd0;
    end
    else if (wr_state_en)
    begin
        state_mem_f[wr_index_in] <= state_in;
        if (pending && pending_ready && (pending_index != wr_index_in))
        begin
            
            if (data_mem_f[pending_index][117+2])
            begin
                state_mem_f[pending_index] <= 2'd1;
            end
            else
            begin
                state_mem_f[pending_index] <= 2'd0;
            end
        end
    end
    else if (pending && pending_ready)
    begin
        if (data_mem_f[pending_index][117+2])
        begin
            state_mem_f[pending_index] <= 2'd1;
        end
        else
        begin
            state_mem_f[pending_index] <= 2'd0;
        end
    end
    else if (cam_en && hit && (data_mem_f[hit_index][59+2:52+2] == 8'd13))
    begin
        state_mem_f[hit_index] <= 2'd2;
    end
    
    else if (wbg_counter_f > 4)
    begin
        if ((state_mem_f[0] == 2'd1) && (data_mem_f[0][59+2:52+2] == 8'd13))
        begin
            state_mem_f[0] <= 2'd2;
        end
        if ((state_mem_f[1] == 2'd1) && (data_mem_f[1][59+2:52+2] == 8'd13))
        begin
            state_mem_f[1] <= 2'd2;
        end
        if ((state_mem_f[2] == 2'd1) && (data_mem_f[2][59+2:52+2] == 8'd13))
        begin
            state_mem_f[2] <= 2'd2;
        end
        if ((state_mem_f[3] == 2'd1) && (data_mem_f[3][59+2:52+2] == 8'd13))
        begin
            state_mem_f[3] <= 2'd2;
        end
        if ((state_mem_f[4] == 2'd1) && (data_mem_f[4][59+2:52+2] == 8'd13))
        begin
            state_mem_f[4] <= 2'd2;
        end
        if ((state_mem_f[5] == 2'd1) && (data_mem_f[5][59+2:52+2] == 8'd13))
        begin
            state_mem_f[5] <= 2'd2;
        end
        if ((state_mem_f[6] == 2'd1) && (data_mem_f[6][59+2:52+2] == 8'd13))
        begin
            state_mem_f[6] <= 2'd2;
        end
        if ((state_mem_f[7] == 2'd1) && (data_mem_f[7][59+2:52+2] == 8'd13))
        begin
            state_mem_f[7] <= 2'd2;
        end
    end
end
always @ *
begin
    if(wr_state_en && wr_data_en && (state_in == 2'd1) 
    && (data_in[59+2:52+2] == 8'd13) && (data_mask_in[59+2:52+2] == {8{1'b1}}))
    begin
        wbg_counter_next = wbg_counter_f + 1;
    end
    else if ((~wr_state_en) && (~(pending && pending_ready)) 
          && (cam_en && hit && (data_mem_f[hit_index][59+2:52+2] == 8'd13)))
    begin
        wbg_counter_next = wbg_counter_f - 1;
    end
    else
    begin
        wbg_counter_next = wbg_counter_f;
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        wbg_counter_f <= 0;
    end
    else   
    begin
        wbg_counter_f <= wbg_counter_next;
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        counter_mem_f[0] <= {6{1'b0}};
        counter_mem_f[1] <= {6{1'b0}};
        counter_mem_f[2] <= {6{1'b0}};
        counter_mem_f[3] <= {6{1'b0}};
        counter_mem_f[4] <= {6{1'b0}};
        counter_mem_f[5] <= {6{1'b0}};
        counter_mem_f[6] <= {6{1'b0}};
        counter_mem_f[7] <= {6{1'b0}};
    end
    else if (pending && pending_ready)
    begin
        counter_mem_f[pending_index] <= {6{1'b0}};
        if (inc_counter_en && (pending_index != wr_index_in))
        begin
            counter_mem_f[wr_index_in] <= counter_mem_f[wr_index_in] + 1;
        end
    end
    else if (inc_counter_en)
    begin
        counter_mem_f[wr_index_in] <= counter_mem_f[wr_index_in] + 1;
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        data_mem_f[0] <= {120+2{1'b0}};
        data_mem_f[1] <= {120+2{1'b0}};
        data_mem_f[2] <= {120+2{1'b0}};
        data_mem_f[3] <= {120+2{1'b0}};
        data_mem_f[4] <= {120+2{1'b0}};
        data_mem_f[5] <= {120+2{1'b0}};
        data_mem_f[6] <= {120+2{1'b0}};
        data_mem_f[7] <= {120+2{1'b0}};
    end
    else if (wr_data_en)
    begin
        data_mem_f[wr_index_in] <= (data_mem_f[wr_index_in] & (~data_mask_in))
                                 | (data_in & data_mask_in);
    end
    else
    begin
        data_mem_f[wr_index_in] <= data_mem_f[wr_index_in];
    end
end
endmodule
      
 
module l2_mshr_wrap(
    input wire clk,
    input wire rst_n,
 
    input wire pipe_wr_sel,
 
    input wire cam_en1,
    input wire wr_state_en1,
    input wire wr_data_en1,
    input wire pending_ready1,
    input wire [2-1:0] state_in1,
    input wire [120+2-1:0] data_in1,
    input wire [120+2-1:0] data_mask_in1,
 
    input wire [3-1:0] inv_counter_rd_index_in1,
    input wire [3-1:0] wr_index_in1,
    input wire [8-1:0] addr_in1,
 
    input wire wr_state_en2,
    input wire wr_data_en2,
 
    input wire inc_counter_en2,
    input wire [2-1:0] state_in2,
    input wire [120+2-1:0] data_in2,
    input wire [120+2-1:0] data_mask_in2,
    input wire [3-1:0] rd_index_in2,
    input wire [3-1:0] wr_index_in2,
 
    output reg hit,
    output reg [3-1:0] hit_index,
    output reg [2-1:0] rd_state_out,
    output reg [120+2-1:0] rd_data_out,
    
    output reg [120+2-1:0] cam_data_out,
    output reg [120+2-1:0] pending_data_out,
    output reg [6-1:0] inv_counter_out,
    output reg [3:0] empty_slots,
    output reg pending,
    output reg [3-1:0] pending_index,
    output reg [3-1:0] empty_index
 
);
 
reg wr_state_en;
reg wr_data_en;
 
reg [2-1:0] state_in;
reg [120+2-1:0] data_in;
reg [120+2-1:0] data_mask_in;
 
reg [3-1:0] wr_index_in;
 
 
always @ *
begin
    if (pipe_wr_sel)
    begin
        wr_state_en = wr_state_en2;
        wr_data_en = wr_data_en2;
        state_in = state_in2;
        data_in = data_in2;
        data_mask_in = data_mask_in2;
        wr_index_in = wr_index_in2;
    end
    else
    begin
        wr_state_en = wr_state_en1;
        wr_data_en = wr_data_en1;
        state_in = state_in1;
        data_in = data_in1;
        data_mask_in = data_mask_in1;
        wr_index_in = wr_index_in1;
    end
end
reg [2-1:0] state_mem_f [8-1:0];
reg [120+2-1:0] data_mem_f [8-1:0];
reg [6-1:0] counter_mem_f [8-1:0];
reg [3-1:0] wbg_counter_f;
reg [3-1:0] wbg_counter_next;
always @ *
begin
    empty_slots = 0;
    if (state_mem_f[0] == 2'd0)
    begin
        empty_slots = empty_slots + 1;
    end
    if (state_mem_f[1] == 2'd0)
    begin
        empty_slots = empty_slots + 1;
    end
    if (state_mem_f[2] == 2'd0)
    begin
        empty_slots = empty_slots + 1;
    end
    if (state_mem_f[3] == 2'd0)
    begin
        empty_slots = empty_slots + 1;
    end
    if (state_mem_f[4] == 2'd0)
    begin
        empty_slots = empty_slots + 1;
    end
    if (state_mem_f[5] == 2'd0)
    begin
        empty_slots = empty_slots + 1;
    end
    if (state_mem_f[6] == 2'd0)
    begin
        empty_slots = empty_slots + 1;
    end
    if (state_mem_f[7] == 2'd0)
    begin
        empty_slots = empty_slots + 1;
    end
end
always @ *
begin
    if (state_mem_f[0] == 2'd2)
    begin
        pending = 1'b1;
        pending_index = 3'd0;
    end
    else if (state_mem_f[1] == 2'd2)
    begin
        pending = 1'b1;
        pending_index = 3'd1;
    end
    else if (state_mem_f[2] == 2'd2)
    begin
        pending = 1'b1;
        pending_index = 3'd2;
    end
    else if (state_mem_f[3] == 2'd2)
    begin
        pending = 1'b1;
        pending_index = 3'd3;
    end
    else if (state_mem_f[4] == 2'd2)
    begin
        pending = 1'b1;
        pending_index = 3'd4;
    end
    else if (state_mem_f[5] == 2'd2)
    begin
        pending = 1'b1;
        pending_index = 3'd5;
    end
    else if (state_mem_f[6] == 2'd2)
    begin
        pending = 1'b1;
        pending_index = 3'd6;
    end
    else if (state_mem_f[7] == 2'd2)
    begin
        pending = 1'b1;
        pending_index = 3'd7;
    end
    else
    begin
        pending = 1'b0;
        pending_index = 3'd0;
    end
end
always @ *
begin
    if (state_mem_f[0] == 2'd0)
    begin
        empty_index = 3'd0;
    end
    else if (state_mem_f[1] == 2'd0)
    begin
        empty_index = 3'd1;
    end
    else if (state_mem_f[2] == 2'd0)
    begin
        empty_index = 3'd2;
    end
    else if (state_mem_f[3] == 2'd0)
    begin
        empty_index = 3'd3;
    end
    else if (state_mem_f[4] == 2'd0)
    begin
        empty_index = 3'd4;
    end
    else if (state_mem_f[5] == 2'd0)
    begin
        empty_index = 3'd5;
    end
    else if (state_mem_f[6] == 2'd0)
    begin
        empty_index = 3'd6;
    end
    else if (state_mem_f[7] == 2'd0)
    begin
        empty_index = 3'd7;
    end
    else
    begin
        empty_index = 3'd0;
    end
end
always @ *
begin
    
    
    rd_state_out = state_mem_f[rd_index_in2];
    rd_data_out = data_mem_f[rd_index_in2];
    
    
    
    
    
    cam_data_out = data_mem_f[hit_index];
    
    
    
    
    pending_data_out = data_mem_f[pending_index];
    
    
    
    
    
    
end
always @ *
begin
    inv_counter_out = counter_mem_f[inv_counter_rd_index_in1];
end
always @ *
begin
    if(cam_en1)
    begin
        if ((data_mem_f[0][6+8-1:6] == addr_in1) && (state_mem_f[0] != 2'd0))
        begin
            hit = 1'b1;
            hit_index = 3'd0;
        end
        else if ((data_mem_f[1][6+8-1:6] == addr_in1) && (state_mem_f[1] != 2'd0))
        begin
            hit = 1'b1;
            hit_index = 3'd1;
        end
        else if ((data_mem_f[2][6+8-1:6] == addr_in1) && (state_mem_f[2] != 2'd0))
        begin
            hit = 1'b1;
            hit_index = 3'd2;
        end
        else if ((data_mem_f[3][6+8-1:6] == addr_in1) && (state_mem_f[3] != 2'd0))
        begin
            hit = 1'b1;
            hit_index = 3'd3;
        end
        else if ((data_mem_f[4][6+8-1:6] == addr_in1) && (state_mem_f[4] != 2'd0))
        begin
            hit = 1'b1;
            hit_index = 3'd4;
        end
        else if ((data_mem_f[5][6+8-1:6] == addr_in1) && (state_mem_f[5] != 2'd0))
        begin
            hit = 1'b1;
            hit_index = 3'd5;
        end
        else if ((data_mem_f[6][6+8-1:6] == addr_in1) && (state_mem_f[6] != 2'd0))
        begin
            hit = 1'b1;
            hit_index = 3'd6;
        end
        else if ((data_mem_f[7][6+8-1:6] == addr_in1) && (state_mem_f[7] != 2'd0))
        begin
            hit = 1'b1;
            hit_index = 3'd7;
        end
        else
        begin
            hit = 1'b0;
            hit_index = 3'd0;
        end
    end
    else
    begin
        hit = 1'b0;
        hit_index = 3'd0;
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        state_mem_f[0] <= 2'd0;
        state_mem_f[1] <= 2'd0;
        state_mem_f[2] <= 2'd0;
        state_mem_f[3] <= 2'd0;
        state_mem_f[4] <= 2'd0;
        state_mem_f[5] <= 2'd0;
        state_mem_f[6] <= 2'd0;
        state_mem_f[7] <= 2'd0;
    end
    else if (wr_state_en)
    begin
        state_mem_f[wr_index_in] <= state_in;
        if (pending && pending_ready1 && (pending_index != wr_index_in))
        begin
            
            if (data_mem_f[pending_index][117+2])
            begin
                state_mem_f[pending_index] <= 2'd1;
            end
            else
            begin
                state_mem_f[pending_index] <= 2'd0;
            end
        end
    end
    else if (pending && pending_ready1)
    begin
        if (data_mem_f[pending_index][117+2])
        begin
            state_mem_f[pending_index] <= 2'd1;
        end
        else
        begin
            state_mem_f[pending_index] <= 2'd0;
        end
    end
    else if (cam_en1 && hit && (data_mem_f[hit_index][59+2:52+2] == 8'd13))
    begin
        state_mem_f[hit_index] <= 2'd2;
    end
    
    else if (wbg_counter_f > 4)
    begin
        if ((state_mem_f[0] == 2'd1) && (data_mem_f[0][59+2:52+2] == 8'd13))
        begin
            state_mem_f[0] <= 2'd2;
        end
        if ((state_mem_f[1] == 2'd1) && (data_mem_f[1][59+2:52+2] == 8'd13))
        begin
            state_mem_f[1] <= 2'd2;
        end
        if ((state_mem_f[2] == 2'd1) && (data_mem_f[2][59+2:52+2] == 8'd13))
        begin
            state_mem_f[2] <= 2'd2;
        end
        if ((state_mem_f[3] == 2'd1) && (data_mem_f[3][59+2:52+2] == 8'd13))
        begin
            state_mem_f[3] <= 2'd2;
        end
        if ((state_mem_f[4] == 2'd1) && (data_mem_f[4][59+2:52+2] == 8'd13))
        begin
            state_mem_f[4] <= 2'd2;
        end
        if ((state_mem_f[5] == 2'd1) && (data_mem_f[5][59+2:52+2] == 8'd13))
        begin
            state_mem_f[5] <= 2'd2;
        end
        if ((state_mem_f[6] == 2'd1) && (data_mem_f[6][59+2:52+2] == 8'd13))
        begin
            state_mem_f[6] <= 2'd2;
        end
        if ((state_mem_f[7] == 2'd1) && (data_mem_f[7][59+2:52+2] == 8'd13))
        begin
            state_mem_f[7] <= 2'd2;
        end
    end
end
always @ *
begin
    if(wr_state_en && wr_data_en && (state_in == 2'd1) 
    && (data_in[59+2:52+2] == 8'd13) && (data_mask_in[59+2:52+2] == {8{1'b1}}))
    begin
        wbg_counter_next = wbg_counter_f + 1;
    end
    else if ((~wr_state_en) && (~(pending && pending_ready1)) 
          && (cam_en1 && hit && (data_mem_f[hit_index][59+2:52+2] == 8'd13)))
    begin
        wbg_counter_next = wbg_counter_f - 1;
    end
    else
    begin
        wbg_counter_next = wbg_counter_f;
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        wbg_counter_f <= 0;
    end
    else   
    begin
        wbg_counter_f <= wbg_counter_next;
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        counter_mem_f[0] <= {6{1'b0}};
        counter_mem_f[1] <= {6{1'b0}};
        counter_mem_f[2] <= {6{1'b0}};
        counter_mem_f[3] <= {6{1'b0}};
        counter_mem_f[4] <= {6{1'b0}};
        counter_mem_f[5] <= {6{1'b0}};
        counter_mem_f[6] <= {6{1'b0}};
        counter_mem_f[7] <= {6{1'b0}};
    end
    else if (pending && pending_ready1)
    begin
        counter_mem_f[pending_index] <= {6{1'b0}};
        if (inc_counter_en2 && (pending_index != wr_index_in))
        begin
            counter_mem_f[wr_index_in] <= counter_mem_f[wr_index_in] + 1;
        end
    end
    else if (inc_counter_en2)
    begin
        counter_mem_f[wr_index_in] <= counter_mem_f[wr_index_in] + 1;
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        data_mem_f[0] <= {120+2{1'b0}};
        data_mem_f[1] <= {120+2{1'b0}};
        data_mem_f[2] <= {120+2{1'b0}};
        data_mem_f[3] <= {120+2{1'b0}};
        data_mem_f[4] <= {120+2{1'b0}};
        data_mem_f[5] <= {120+2{1'b0}};
        data_mem_f[6] <= {120+2{1'b0}};
        data_mem_f[7] <= {120+2{1'b0}};
    end
    else if (wr_data_en)
    begin
        data_mem_f[wr_index_in] <= (data_mem_f[wr_index_in] & (~data_mask_in))
                                 | (data_in & data_mask_in);
    end
    else
    begin
        data_mem_f[wr_index_in] <= data_mem_f[wr_index_in];
    end
end
 
endmodule
      
 
module l2_pipe1_buf_in(
    input wire clk,
    input wire rst_n,
    input wire valid_in,
    input wire [64-1:0] data_in,
    output reg ready_in,
   
    output reg msg_header_valid_out,
    output reg [192-1:0] msg_header_out,
    input wire msg_header_ready_out,
    output reg msg_data_valid_out,
    output reg [64-1:0] msg_data_out,
    input wire msg_data_ready_out
);
localparam msg_data_state0 = 2'd0;
localparam msg_data_state1 = 2'd1;
localparam msg_data_state2 = 2'd2;
localparam msg_state_header0 = 3'd0;
localparam msg_state_header1 = 3'd1;
localparam msg_state_header2 = 3'd2;
localparam msg_state_data0 = 3'd3;
localparam msg_state_data1 = 3'd4;
reg [2:0] msg_state_f;
reg [2:0] msg_state_next;
reg real_ready_in;
reg [1:0] msg_data_state_f;
reg [1:0] msg_data_state_next;
reg [2:0] msg_int_state_f;
reg [2:0] msg_int_state_next;
reg int_stall;
always @ *
begin
    if (!rst_n)
    begin
        msg_data_state_next = msg_data_state0;
    end
    else if((msg_state_f == msg_state_header0) && valid_in)
    begin
        if (data_in[21:14] == 8'd32)
        begin
            msg_data_state_next = msg_data_state1;
        end
        else
        begin
            msg_data_state_next = data_in[29:22] - 2;
        end
    end
    else
    begin
        msg_data_state_next = msg_data_state_f;
    end
end
always @ (posedge clk)
begin
    msg_data_state_f <= msg_data_state_next;
end
always @ *
begin
    if (!rst_n)
    begin
        msg_state_next = msg_state_header0;
    end
    else if (valid_in && real_ready_in)
    begin
        if ((msg_state_f == msg_state_header2) && (msg_data_state_f == msg_data_state0))
        begin
            msg_state_next = msg_state_header0;
        end
        else if ((msg_state_f == msg_state_data0) && (msg_data_state_f == msg_data_state1))
        begin
            msg_state_next = msg_state_header0;
        end
        else
        begin
            if (msg_state_f == msg_state_data1)
            begin
                msg_state_next = msg_state_header0;
            end
            else
            begin
                msg_state_next = msg_state_f + 3'd1;
            end
        end
    end
    else
    begin
        msg_state_next = msg_state_f;
    end 
end
always @ (posedge clk)
begin
    msg_state_f <= msg_state_next;
end
always @ *
begin
    if (!rst_n)
    begin
        msg_int_state_next = msg_state_header0;
    end
    else if (valid_in && real_ready_in && (data_in[21:14] == 8'd32) 
         && (msg_state_f == msg_state_header0))
    begin
        msg_int_state_next = msg_state_header1;
    end
    else if (valid_in && real_ready_in && (msg_int_state_f == msg_state_header1))
    begin
        msg_int_state_next = msg_state_header2;
    end
    else if (valid_in && real_ready_in && (msg_int_state_f == msg_state_header2))
    begin
        msg_int_state_next = msg_state_header0;
    end
    else
    begin
        msg_int_state_next = msg_int_state_f;
    end 
end
always @ (posedge clk)
begin
    msg_int_state_f <= msg_int_state_next;
end
always @ *
begin
    if ((valid_in && (data_in[21:14] == 8'd32) && (msg_state_f == msg_state_header0))
    || (msg_int_state_f == msg_state_header1))
    begin
        int_stall = 1'b1;
    end
    else
    begin
        int_stall = 1'b0;
    end
end
localparam msg_mux_header = 1'b0;
localparam msg_mux_data = 1'b1;
reg msg_mux_sel;
always @ *
begin
    if ((msg_state_f == msg_state_header0)
    ||  (msg_state_f == msg_state_header1)
    ||  (msg_state_f == msg_state_header2))
    begin
        msg_mux_sel = msg_mux_header;
    end
    else
        msg_mux_sel = msg_mux_data;
end
reg msg_header_valid_in;
reg [64-1:0] msg_header_in;
reg msg_header_ready_in;
reg msg_data_valid_in;
reg [64-1:0] msg_data_in;
reg msg_data_ready_in;
always @ *
begin
    if (msg_mux_sel == msg_mux_header)
    begin
        msg_header_valid_in = valid_in;
        msg_header_in = data_in;
    end
    else
    begin
        msg_header_valid_in = 0;
        msg_header_in = 0;
    end
end
always @ *
begin
    if (msg_mux_sel == msg_mux_data)
    begin
        msg_data_valid_in = valid_in;
        msg_data_in = data_in;
    end
    else
    begin
        msg_data_valid_in = 0;
        msg_data_in = 0;
    end
end
always @ *
begin
    if (msg_mux_sel == msg_mux_data)
    begin
        real_ready_in = msg_data_ready_in; 
    end
    else
    begin
        real_ready_in = msg_header_ready_in;
    end
end
always @ *
begin
    ready_in = real_ready_in && (!int_stall);
end
reg [64-1:0] header_buf_mem_f [8-1:0];
reg header_buf_empty;
reg header_buf_full;
reg [3:0] header_buf_counter_f;
reg [3:0] header_buf_counter_next;
reg [3-1:0] header_rd_ptr_f;
reg [3-1:0] header_rd_ptr_next;
reg [3-1:0] header_rd_ptr_plus1;
reg [3-1:0] header_rd_ptr_plus2;
reg [3-1:0] header_wr_ptr_f;
reg [3-1:0] header_wr_ptr_next;
always @ *
begin
    header_buf_empty = (header_buf_counter_f == 0);
    header_buf_full = (header_buf_counter_f ==  8);
end
always @ *
begin
    if ((msg_header_valid_in && msg_header_ready_in) && (msg_header_valid_out && msg_header_ready_out))
    begin
        header_buf_counter_next = header_buf_counter_f + 1 - 3;
    end
    else if (msg_header_valid_in && msg_header_ready_in)
    begin 
        header_buf_counter_next = header_buf_counter_f + 1;
    end
    else if (msg_header_valid_out && msg_header_ready_out)
    begin 
        header_buf_counter_next = header_buf_counter_f - 3;
    end
    else
    begin
        header_buf_counter_next = header_buf_counter_f;
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        header_buf_counter_f <= 0;
    end
    else
    begin
        header_buf_counter_f <= header_buf_counter_next;
    end
end
always @ *
begin
    if (!rst_n)
    begin   
        header_rd_ptr_next = 0;
    end
    else if (msg_header_valid_out && msg_header_ready_out)
    begin
        header_rd_ptr_next = header_rd_ptr_f + 3;
    end
    else
    begin
        header_rd_ptr_next = header_rd_ptr_f;
    end
end
always @ (posedge clk)
begin
    header_rd_ptr_f <= header_rd_ptr_next;
end
always @ *
begin
    if (!rst_n)
    begin   
        header_wr_ptr_next = 0;
    end
    else if (msg_header_valid_in && msg_header_ready_in)
    begin
        header_wr_ptr_next = header_wr_ptr_f + 1;
    end
    else
    begin
        header_wr_ptr_next = header_wr_ptr_f;
    end
end
always @ (posedge clk)
begin
    header_wr_ptr_f <= header_wr_ptr_next;
end
always @ *
begin
    header_rd_ptr_plus1 = header_rd_ptr_f + 1;
    header_rd_ptr_plus2 = header_rd_ptr_f + 2;
end
always @ *
begin
   msg_header_ready_in = !header_buf_full;
end
always @ *
begin
    msg_header_valid_out = (header_buf_counter_f >= 3);
    msg_header_out = {header_buf_mem_f[header_rd_ptr_plus2], 
                      header_buf_mem_f[header_rd_ptr_plus1], 
                      header_buf_mem_f[header_rd_ptr_f]};
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin   
        header_buf_mem_f[0] <= 0;
        header_buf_mem_f[1] <= 0;
        header_buf_mem_f[2] <= 0;
        header_buf_mem_f[3] <= 0;
        header_buf_mem_f[4] <= 0;
        header_buf_mem_f[5] <= 0;
        header_buf_mem_f[6] <= 0;
        header_buf_mem_f[7] <= 0;
    end
    else if (msg_header_valid_in && msg_header_ready_in)
    begin
        header_buf_mem_f[header_wr_ptr_f] <= msg_header_in;
    end
    else
    begin 
        header_buf_mem_f[header_wr_ptr_f] <= header_buf_mem_f[header_wr_ptr_f];
    end
end
reg [64-1:0] data_buf_mem_f [4-1:0];
reg data_buf_empty;
reg data_buf_full;
reg [2:0] data_buf_counter_f;
reg [2:0] data_buf_counter_next;
reg [2-1:0] data_rd_ptr_f;
reg [2-1:0] data_rd_ptr_next;
reg [2-1:0] data_wr_ptr_f;
reg [2-1:0] data_wr_ptr_next;
always @ *
begin
    data_buf_empty = (data_buf_counter_f == 0);
    data_buf_full = (data_buf_counter_f ==  4);
end
always @ *
begin
    if (!rst_n)
    begin
        data_buf_counter_next = 0;
    end
    else if ((msg_data_valid_in && msg_data_ready_in) && (msg_data_valid_out && msg_data_ready_out))
    begin
        data_buf_counter_next = data_buf_counter_f + 1 - 1;
    end
    else if (msg_data_valid_in && msg_data_ready_in)
    begin 
        data_buf_counter_next = data_buf_counter_f + 1;
    end
    else if (msg_data_valid_out && msg_data_ready_out)
    begin 
        data_buf_counter_next = data_buf_counter_f - 1;
    end
    else
    begin
        data_buf_counter_next = data_buf_counter_f;
    end
end
always @ (posedge clk)
begin
    data_buf_counter_f <= data_buf_counter_next;
end
always @ *
begin
    if (!rst_n)
    begin   
        data_rd_ptr_next = 0;
    end
    else if (msg_data_valid_out && msg_data_ready_out)
    begin
        data_rd_ptr_next = data_rd_ptr_f + 1;
    end
    else
    begin
        data_rd_ptr_next = data_rd_ptr_f;
    end
end
always @ (posedge clk)
begin
    data_rd_ptr_f <= data_rd_ptr_next;
end
always @ *
begin
    if (!rst_n)
    begin   
        data_wr_ptr_next = 0;
    end
    else if (msg_data_valid_in && msg_data_ready_in)
    begin
        data_wr_ptr_next = data_wr_ptr_f + 1;
    end
    else
    begin
        data_wr_ptr_next = data_wr_ptr_f;
    end
end
always @ (posedge clk)
begin
    data_wr_ptr_f <= data_wr_ptr_next;
end
always @ *
begin
   msg_data_ready_in = !data_buf_full;
end
always @ *
begin
    msg_data_valid_out = !data_buf_empty;
    msg_data_out = data_buf_mem_f[data_rd_ptr_f]; 
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin   
        data_buf_mem_f[0] <= 0;
        data_buf_mem_f[1] <= 0;
        data_buf_mem_f[2] <= 0;
        data_buf_mem_f[3] <= 0;
    end
    else if (msg_data_valid_in && msg_data_ready_in)
    begin
        data_buf_mem_f[data_wr_ptr_f] <= msg_data_in;
    end
    else
    begin 
        data_buf_mem_f[data_wr_ptr_f] <= data_buf_mem_f[data_wr_ptr_f];
    end
end
endmodule
      
 
module l2_pipe1_buf_out(
    input wire clk,
    input wire rst_n,
    input wire [3-1:0] mode_in,
    input wire valid_in,
    input wire [320 -1:0] data_in,
    output reg ready_in,
   
    output reg valid_out,
    output reg [64-1:0] data_out,
    input wire ready_out
);
reg [64-1:0] buf_mem_f [16-1:0];
reg buf_empty;
reg buf_full;
reg [4:0] buf_counter_f;
reg [4:0] buf_counter_next;
reg [4-1:0] rd_ptr_f;
reg [4-1:0] rd_ptr_next;
reg [4-1:0] wr_ptr_f;
reg [4-1:0] wr_ptr_next;
reg [4-1:0] wr_ptr_plus1;
reg [4-1:0] wr_ptr_plus2;
reg [4-1:0] wr_ptr_plus3;
reg [4-1:0] wr_ptr_plus4;
reg [4:0] buf_rd_flits;
always @ *
begin
    if (mode_in == 3'd1)
    begin
        buf_rd_flits = 1;
    end
    else if (mode_in == 3'd2)
    begin
        buf_rd_flits = 2;
    end
    else if (mode_in == 3'd3)
    begin
        buf_rd_flits = 3;
    end
    else if (mode_in == 3'd4)
    begin
        buf_rd_flits = 3;
    end
    else if (mode_in == 3'd5)
    begin
        buf_rd_flits = 4;
    end
    else if (mode_in == 3'd6)
    begin
        buf_rd_flits = 5;
    end
    else if (mode_in == 3'd7)
    begin
        buf_rd_flits = 2;
    end
    else
    begin
        buf_rd_flits = 0;
    end
end
always @ *
begin
   buf_empty = (buf_counter_f == 0);
   buf_full = (buf_counter_f ==  16);
end
always @ *
begin
    if (!rst_n)
    begin
        buf_counter_next = 0;
    end
    else if ((valid_in && ready_in) && (valid_out && ready_out))
    begin
        buf_counter_next = buf_counter_f + buf_rd_flits - 1;
    end
    else if (valid_in && ready_in)
    begin 
        buf_counter_next = buf_counter_f + buf_rd_flits;
    end
    else if (valid_out && ready_out)
    begin 
        buf_counter_next = buf_counter_f - 1;
    end
    else
    begin
        buf_counter_next = buf_counter_f;
    end
end
always @ (posedge clk)
begin
    buf_counter_f <= buf_counter_next;
end
always @ *
begin
    if (!rst_n)
    begin   
        rd_ptr_next = 0;
    end
    else if (valid_out && ready_out)
    begin
        rd_ptr_next = rd_ptr_f + 1;
    end
    else
    begin
        rd_ptr_next = rd_ptr_f;
    end
end
always @ (posedge clk)
begin
    rd_ptr_f <= rd_ptr_next;
end
always @ *
begin
    if (!rst_n)
    begin   
        wr_ptr_next = 0;
    end
    else if (valid_in && ready_in)
    begin
        wr_ptr_next = wr_ptr_f + buf_rd_flits;
    end
    else
    begin
        wr_ptr_next = wr_ptr_f;
    end
end
always @ (posedge clk)
begin
    wr_ptr_f <= wr_ptr_next;
end
always @ *
begin
    wr_ptr_plus1 = wr_ptr_f + 1;
    wr_ptr_plus2 = wr_ptr_f + 2;
    wr_ptr_plus3 = wr_ptr_f + 3;
    wr_ptr_plus4 = wr_ptr_f + 4;
end
always @ *
begin
    ready_in = (buf_counter_f <= 16 - buf_rd_flits);
end
always @ *
begin
    valid_out = !buf_empty;
    data_out = buf_mem_f[rd_ptr_f]; 
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin  
        buf_mem_f[0] <= 0;
        buf_mem_f[1] <= 0;
        buf_mem_f[2] <= 0;
        buf_mem_f[3] <= 0;
        buf_mem_f[4] <= 0;
        buf_mem_f[5] <= 0;
        buf_mem_f[6] <= 0;
        buf_mem_f[7] <= 0;
        buf_mem_f[8] <= 0;
        buf_mem_f[9] <= 0;
        buf_mem_f[10] <= 0;
        buf_mem_f[11] <= 0;
        buf_mem_f[12] <= 0;
        buf_mem_f[13] <= 0;
        buf_mem_f[14] <= 0;
        buf_mem_f[15] <= 0;
    end
    else if (valid_in && ready_in)
    begin
        if (mode_in == 3'd1)
        begin
            buf_mem_f[wr_ptr_f] <= data_in[64-1:0];
        end
        else if (mode_in == 3'd2)
        begin
            buf_mem_f[wr_ptr_f] <= data_in[64-1:0];
            buf_mem_f[wr_ptr_plus1] <= data_in[64*4-1:64*3];
        end
        else if (mode_in == 3'd7)
        begin
            buf_mem_f[wr_ptr_f] <= data_in[64*4-1:64*3];
            buf_mem_f[wr_ptr_plus1] <= data_in[64*5-1:64*4];
        end
        else if (mode_in == 3'd4)
        begin
            buf_mem_f[wr_ptr_f] <= data_in[64-1:0];
            buf_mem_f[wr_ptr_plus1] <= data_in[64*2-1:64];
            buf_mem_f[wr_ptr_plus2] <= data_in[64*3-1:64*2];
        end
        else if (mode_in == 3'd3)
        begin
            buf_mem_f[wr_ptr_f] <= data_in[64-1:0];
            buf_mem_f[wr_ptr_plus1] <= data_in[64*4-1:64*3];
            buf_mem_f[wr_ptr_plus2] <= data_in[64*5-1:64*4];
        end
        else if (mode_in == 3'd5)
        begin
            buf_mem_f[wr_ptr_f] <= data_in[64-1:0];
            buf_mem_f[wr_ptr_plus1] <= data_in[64*2-1:64];
            buf_mem_f[wr_ptr_plus2] <= data_in[64*3-1:64*2];
            buf_mem_f[wr_ptr_plus3] <= data_in[64*4-1:64*3];
        end
        else if (mode_in == 3'd6)
        begin
            buf_mem_f[wr_ptr_f] <= data_in[64-1:0];
            buf_mem_f[wr_ptr_plus1] <= data_in[64*2-1:64];
            buf_mem_f[wr_ptr_plus2] <= data_in[64*3-1:64*2];
            buf_mem_f[wr_ptr_plus3] <= data_in[64*4-1:64*3];
            buf_mem_f[wr_ptr_plus4] <= data_in[64*5-1:64*4];
        end
    end
end
endmodule
      
 
module l2_pipe1_ctrl(
    input wire clk,
    input wire rst_n,
    
    input wire csm_en,
    
    
    input wire pipe2_valid_S1,
    input wire pipe2_valid_S2,
    input wire pipe2_valid_S3,
    input wire [8-1:0] pipe2_msg_type_S1,
    input wire [8-1:0] pipe2_msg_type_S2,
    input wire [8-1:0] pipe2_msg_type_S3,
    input wire [40-1:0] pipe2_addr_S1,
    input wire [40-1:0] pipe2_addr_S2,
    input wire [40-1:0] pipe2_addr_S3,
    
    input wire global_stall_S1,
    
    input wire msg_header_valid_S1,
    input wire [8-1:0] msg_type_S1,
    input wire [3-1:0] msg_data_size_S1,
    input wire [1-1:0] msg_cache_type_S1,
    
    input wire mshr_hit_S1,
 
    input wire mshr_pending_S1,
    input wire [3-1:0] mshr_pending_index_S1,
    input wire [3:0] mshr_empty_slots_S1,
    
 
    
    
    input wire [8-1:0] cam_mshr_msg_type_S1,
    input wire [1-1:0] cam_mshr_l2_miss_S1,
    input wire [3-1:0] cam_mshr_data_size_S1,
    input wire [1-1:0] cam_mshr_cache_type_S1,
    
    input wire cam_mshr_smc_miss_S1,
    
    
    input wire [8-1:0] pending_mshr_msg_type_S1,
    input wire [1-1:0] pending_mshr_l2_miss_S1,
    input wire [3-1:0] pending_mshr_data_size_S1,
    input wire [1-1:0] pending_mshr_cache_type_S1,
    
    input wire pending_mshr_smc_miss_S1,
    
 
    
    input wire msg_data_valid_S1,
    input wire [40-1:0] addr_S1,
    
    
    input wire global_stall_S2,
    
    input wire l2_tag_hit_S2,
    input wire l2_evict_S2,
    input wire l2_wb_S2,
    input wire [2-1:0] l2_way_state_mesi_S2,
    input wire [2-1:0] l2_way_state_vd_S2,
    input wire [1-1:0] l2_way_state_cache_type_S2,
    input wire [4-1:0] l2_way_state_subline_S2,
    input wire req_from_owner_S2,
    input wire addr_l2_aligned_S2,
    input wire [6-1:0] lsid_S2,
    
    input wire msg_data_valid_S2,
    input wire [40-1:0] addr_S2,
    
    
    
    
    input wire [64-1:0] dir_data_S3,
    input wire [40-1:0] addr_S3,
    
    
    input wire global_stall_S4,
    
    input wire [3-1:0] mshr_empty_index_S4,
    
    input wire l2_tag_hit_S4,
    input wire l2_evict_S4,
    input wire [2-1:0] l2_way_state_mesi_S4,
    input wire [6-1:0] l2_way_state_owner_S4,
    input wire [2-1:0] l2_way_state_vd_S4,
    input wire [4-1:0] l2_way_state_subline_S4,
    input wire [1-1:0] l2_way_state_cache_type_S4,
    input wire [8-1:0] mshrid_S4,
    input wire req_from_owner_S4,
    input wire [6-1:0] mshr_miss_lsid_S4,
    input wire [6-1:0] lsid_S4,
    
    input wire broadcast_counter_zero_S4,
    input wire broadcast_counter_max_S4,
    input wire broadcast_counter_avail_S4,
    input wire [14-1:0] broadcast_chipid_out_S4,
    input wire [8-1:0] broadcast_x_out_S4,
    input wire [8-1:0] broadcast_y_out_S4,
    
    input wire [40-1:0] addr_S4,
    
    input wire cas_cmp_S4,
    
    input wire msg_send_ready_S4,
    
    
    input wire smc_hit_S4,
    
    
    output reg valid_S1,
    output reg stall_S1,
    output reg msg_from_mshr_S1,
    output reg dis_flush_S1,
    output reg mshr_cam_en_S1,
    output reg mshr_pending_ready_S1,
    output reg msg_header_ready_S1,
    output reg tag_clk_en_S1,
    output reg tag_rdw_en_S1,
    output reg state_rd_en_S1,
    output reg reg_wr_en_S1,
    output reg [8-1:0] reg_wr_addr_type_S1,
    
    output reg valid_S2,
    output reg stall_S2,
    output reg stall_before_S2,
    output reg stall_real_S2,
    output reg [8-1:0] msg_type_S2,
    output reg msg_from_mshr_S2,
    output reg special_addr_type_S2,
    output wire state_load_sdid_S2,
    output reg dir_clk_en_S2,
    output reg dir_rdw_en_S2,
    output reg [2-1:0] dir_op_S2,
    output reg data_clk_en_S2,
    output reg data_rdw_en_S2,
    output reg [4-1:0] amo_alu_op_S2,
    output reg [3-1:0] data_size_S2,
    output reg [1-1:0] cache_type_S2,
    output reg state_owner_en_S2,
    output reg [2-1:0] state_owner_op_S2,
    output reg state_subline_en_S2,
    output reg [2-1:0] state_subline_op_S2,
    output reg state_di_en_S2,
    output reg state_vd_en_S2,
    output reg [2-1:0] state_vd_S2,
    output reg state_mesi_en_S2,
    output reg [2-1:0] state_mesi_S2,
    output reg state_lru_en_S2,
    output reg [1-1:0] state_lru_op_S2,
    output reg state_rb_en_S2,
    output reg [2-1:0] l2_load_data_subline_S2,
    output reg l2_ifill_32B_S2,
    output reg msg_data_ready_S2,
    
    output reg smc_wr_en_S2,
    output reg smc_wr_diag_en_S2,
    output reg smc_flush_en_S2,
    output reg [2-1:0] smc_addr_op_S2,
    
    
    output reg valid_S3,
    output reg stall_S3,
    output reg stall_before_S3,
    
    output reg valid_S4,
    output reg stall_S4,
    output reg stall_before_S4,
    output reg [8-1:0] msg_type_S4,
    output reg [3-1:0] data_size_S4,
    output reg [1-1:0] cache_type_S4,
    output reg [1-1:0] l2_miss_S4,
    
    output reg smc_miss_S4,
    output reg stall_smc_buf_S4,
    
    output reg  msg_from_mshr_S4,
    output reg req_recycle_S4,
    output reg inv_fwd_pending_S4,
    output wire [6-1:0] dir_sharer_S4,
    output reg [6-1:0] dir_sharer_counter_S4,
    output reg [64-1:0] dir_data_sel_S4,
    output reg cas_cmp_en_S4,
    output reg atomic_read_data_en_S4,
    output reg [3-1:0] cas_cmp_data_size_S4,
    output reg [64-1:0] dir_data_S4,
    output reg msg_send_valid_S4,
    output reg [3-1:0] msg_send_mode_S4,
    output reg [8-1:0] msg_send_type_S4,
    output reg [8-1:0] msg_send_type_pre_S4,
    output reg [8-1:0] msg_send_length_S4,
    output reg [3-1:0] msg_send_data_size_S4,
    output reg [1-1:0] msg_send_cache_type_S4,
    output reg [2-1:0] msg_send_mesi_S4,
    output reg [1-1:0] msg_send_l2_miss_S4,
    output reg [8-1:0] msg_send_mshrid_S4,
    output reg [4-1:0] msg_send_subline_vector_S4,
    output reg special_addr_type_S4,
    output reg mshr_wr_data_en_S4,
    output reg mshr_wr_state_en_S4,
    output reg [2-1:0] mshr_state_in_S4,
    output reg [3-1:0] mshr_inv_counter_rd_index_in_S4,
    output reg [3-1:0] mshr_wr_index_in_S4,
    output reg state_wr_sel_S4,
    output reg state_wr_en_S4,
    
    output reg [2-1:0] broadcast_counter_op_S4,
    output reg broadcast_counter_op_val_S4,
    
    
    output reg smc_rd_diag_en_buf_S4,
    output reg smc_rd_en_buf_S4,
    
    output reg l2_access_valid_S4,
    output reg l2_miss_valid_S4,
    output reg reg_rd_en_S4,
    output reg [8-1:0] reg_rd_addr_type_S4
);
localparam y = 1'b1;
localparam n = 1'b0;
localparam rd = 1'b1;
localparam wr = 1'b0;
reg [8-1:0] msg_type_S2_f;
reg msg_from_mshr_S2_f;
reg [8-1:0] msg_type_S4_f;
reg stall_pre_S1;
reg stall_hazard_S1;
reg [8-1:0] msg_type_mux_S1;
reg [8-1:0] msg_type_trans_S1;
reg [3-1:0] data_size_S1;
reg [1-1:0] cache_type_S1;
reg msg_header_ready_real_S1;
reg msg_cas_cmp_S1_f;
reg msg_cas_cmp_S1_next;
reg msg_input_en_S1_f;
reg msg_input_en_S1_next;
reg [8-1:0] addr_type_S1;
reg [2-1:0] addr_op_S1;
reg special_addr_type_S1;
reg msg_data_rd_S1;
always @ *
begin
    valid_S1 = mshr_pending_S1 || (msg_header_valid_S1 && msg_input_en_S1_f);
end
always @ *
begin
    stall_pre_S1 = stall_S2 || global_stall_S1;
end
always @ *
begin
    mshr_pending_ready_S1 = mshr_pending_S1 && (!stall_S1);
end
always @ *
begin
    msg_from_mshr_S1 = mshr_pending_S1;
end
always @ *
begin
    if (msg_from_mshr_S1)
    begin
        msg_type_mux_S1 = pending_mshr_msg_type_S1;
 
    end
    else
    begin
        msg_type_mux_S1 = msg_type_S1;
    end
end
always @ *
begin
     
    
    
    mshr_cam_en_S1 = (!mshr_pending_S1) && msg_header_valid_S1 && (!global_stall_S1);
    
end
localparam atomic_state0 = 1'b0;
localparam atomic_state1 = 1'b1;
reg atomic_state_S1_f;
reg atomic_state_S1_next;
reg [4-1:0] amo_alu_op_S1;
reg [4-1:0] amo_alu_op_S2_f;
always @ *
begin
    amo_alu_op_S1 = 4'd0;
    if (!rst_n)
    begin
        atomic_state_S1_next = atomic_state0;
    end
    else if (valid_S1 && (!msg_from_mshr_S1) &&
       (msg_type_trans_S1 == 8'd6
        || msg_type_trans_S1 == 8'd10
        || msg_type_trans_S1 == 8'd44
        || msg_type_trans_S1 == 8'd45
        || msg_type_trans_S1 == 8'd46
        || msg_type_trans_S1 == 8'd47
        || msg_type_trans_S1 == 8'd48
        || msg_type_trans_S1 == 8'd49
        || msg_type_trans_S1 == 8'd50
        || msg_type_trans_S1 == 8'd51))
    begin
        atomic_state_S1_next = atomic_state1;
    end
    else if (valid_S1 && (!msg_from_mshr_S1) &&
            (msg_type_trans_S1 == 8'd7
            || msg_type_trans_S1 == 8'd8
            || msg_type_trans_S1 == 8'd11
            || msg_type_trans_S1 == 8'd52
            || msg_type_trans_S1 == 8'd53
            || msg_type_trans_S1 == 8'd54
            || msg_type_trans_S1 == 8'd55
            || msg_type_trans_S1 == 8'd56
            || msg_type_trans_S1 == 8'd57
            || msg_type_trans_S1 == 8'd58
            || msg_type_trans_S1 == 8'd59))
    begin
        atomic_state_S1_next = atomic_state0;
        case (msg_type_trans_S1)
            8'd52: begin
                amo_alu_op_S1 = 4'd1;
            end
            8'd53: begin
                amo_alu_op_S1 = 4'd2;
            end
            8'd54: begin
                amo_alu_op_S1 = 4'd3;
            end
            8'd55: begin
                amo_alu_op_S1 = 4'd4;
            end
            8'd56: begin
                amo_alu_op_S1 = 4'd5;
            end
            8'd57: begin
                amo_alu_op_S1 = 4'd6;
            end
            8'd58: begin
                amo_alu_op_S1 = 4'd7;
            end
            8'd59: begin
                amo_alu_op_S1 = 4'd8;
            end
        endcase
    end
    else
    begin
        atomic_state_S1_next = atomic_state_S1_f;
    end
end
always @ (posedge clk)
begin
    if (!stall_S1)
    begin
        atomic_state_S1_f <= atomic_state_S1_next;
    end
end
always @ *
begin
    case (msg_type_mux_S1)
    8'd14:
    begin
        case (addr_type_S1)
        8'hac, 8'had, 8'hae, 8'haf:
        begin
            msg_type_trans_S1 = 8'd35;
        end
        8'ha3:
        begin
            msg_type_trans_S1 = 8'd34;
        end
        default:
        begin
            msg_type_trans_S1 = msg_type_mux_S1;
        end
        endcase
    end
    8'd5:
    begin
        if (atomic_state_S1_f == atomic_state0)
        begin
            msg_type_trans_S1 = 8'd6;
        end
        else
        begin
            if (msg_cas_cmp_S1_f)
            begin
                msg_type_trans_S1 = 8'd7;
            end
            else
            begin
                msg_type_trans_S1 = 8'd8;
            end
        end
    end
    8'd9:
    begin
        if (atomic_state_S1_f == atomic_state0)
        begin
            msg_type_trans_S1 = 8'd10;
        end
        else
        begin
            msg_type_trans_S1 = 8'd11;
        end
    end
    8'd36:
    begin
        if (atomic_state_S1_f == atomic_state0)
        begin
            msg_type_trans_S1 = 8'd44;
        end
        else
        begin
            msg_type_trans_S1 = 8'd52;
        end
    end
    8'd37:
    begin
        if (atomic_state_S1_f == atomic_state0)
        begin
            msg_type_trans_S1 = 8'd45;
        end
        else
        begin
            msg_type_trans_S1 = 8'd53;
        end
    end
    8'd38:
    begin
        if (atomic_state_S1_f == atomic_state0)
        begin
            msg_type_trans_S1 = 8'd46;
        end
        else
        begin
            msg_type_trans_S1 = 8'd54;
        end
    end
    8'd39:
    begin
        if (atomic_state_S1_f == atomic_state0)
        begin
            msg_type_trans_S1 = 8'd47;
        end
        else
        begin
            msg_type_trans_S1 = 8'd55;
        end
    end
    8'd40:
    begin
        if (atomic_state_S1_f == atomic_state0)
        begin
            msg_type_trans_S1 = 8'd48;
        end
        else
        begin
            msg_type_trans_S1 = 8'd56;
        end
    end
    8'd41:
    begin
        if (atomic_state_S1_f == atomic_state0)
        begin
            msg_type_trans_S1 = 8'd49;
        end
        else
        begin
            msg_type_trans_S1 = 8'd57;
        end
    end
    8'd42:
    begin
        if (atomic_state_S1_f == atomic_state0)
        begin
            msg_type_trans_S1 = 8'd50;
        end
        else
        begin
            msg_type_trans_S1 = 8'd58;
        end
    end
    8'd43:
    begin
        if (atomic_state_S1_f == atomic_state0)
        begin
            msg_type_trans_S1 = 8'd51;
        end
        else
        begin
            msg_type_trans_S1 = 8'd59;
        end
    end
    default:
    begin
        msg_type_trans_S1 = msg_type_mux_S1;
    end
    endcase
end
always @ *
begin
    dis_flush_S1 = (msg_type_trans_S1 == 8'd35) && ~msg_from_mshr_S1;
end
always @ *
begin
    addr_type_S1 = addr_S1[39:32];
    addr_op_S1 = addr_S1[31:30];
end
always @ *
begin
    if ((msg_type_trans_S1 == 8'd14 || msg_type_trans_S1 == 8'd15)
    &&  (addr_type_S1 == 8'ha0
    ||   addr_type_S1 == 8'ha4
    ||   addr_type_S1 == 8'ha6
    ||   addr_type_S1 == 8'ha1
    ||   addr_type_S1 == 8'ha2
    ||   addr_type_S1 == 8'ha5
    ||   addr_type_S1 == 8'haa
    ||   addr_type_S1 == 8'hab
    ||   addr_type_S1 == 8'ha7
    ||   addr_type_S1 == 8'ha8
    ||   addr_type_S1 == 8'ha9))
    begin
        special_addr_type_S1 = 1'b1;
    end
    else
    begin
        special_addr_type_S1 = 1'b0;
    end
end
always @ *
begin
    if (msg_from_mshr_S1)
    begin
        data_size_S1 = pending_mshr_data_size_S1;
 
    end
    else
    begin
        data_size_S1 = msg_data_size_S1;
    end
end
always @ *
begin
    if (msg_from_mshr_S1)
    begin
        cache_type_S1 = pending_mshr_cache_type_S1;
 
    end
    else
    begin
        cache_type_S1 = msg_cache_type_S1;
    end
end
reg [3-1:0] cs_S1;
always @ *
begin
    cs_S1 = {3{1'bx}};
    if (valid_S1)
    begin
        if (special_addr_type_S1)
        begin
            case (addr_type_S1)
                8'ha4:
                begin
                    if (msg_type_trans_S1 == 8'd14)
                    begin
                        
                        cs_S1 = {y,             rd,       n};
                    end
                    else
                    begin
                        cs_S1 = {y,             wr,        n};
                    end
                end
                8'ha6:
                begin
                    if (msg_type_trans_S1 == 8'd14)
                    begin
                        
                        cs_S1 = {y,             rd,      y};
                    end
                    else
                    begin
                        cs_S1 = {n,             rd,       n};
                    end
                end
                default:
                begin
                    cs_S1 = {n,             rd,           n};
                end
            endcase
        end
        else
        begin
            case (msg_type_trans_S1)
                8'd31, 8'd14, 8'd15, 8'd1,
                8'd2,
                8'd60,
                8'd13, 8'd7, 8'd11,
                8'd6, 8'd10, 8'd35,8'd34,
                8'd44, 8'd52,
                8'd45, 8'd53,
                8'd46, 8'd54,
                8'd47, 8'd55,
                8'd48, 8'd56,
                8'd49, 8'd57,
                8'd50, 8'd58,
                8'd51, 8'd59:
                begin
                
                    cs_S1 = {y,             rd,     y};
                end
                8'd30, 8'd8, 8'd32:
                begin
                    cs_S1 = {n,             rd,          n};
                end
                default:
                begin
                    cs_S1 = {3{1'bx}};
                end
            endcase
        end
    end
    else
    begin
        cs_S1 = {3{1'b0}};
    end
end
always @ *
begin
    if (!rst_n)
    begin
        msg_input_en_S1_next = y;
    end
    else if ((valid_S1 && !stall_S1)
           &&((msg_type_trans_S1 == 8'd7)
           || (msg_type_trans_S1 == 8'd11)
           || (msg_type_trans_S1 == 8'd52)
           || (msg_type_trans_S1 == 8'd53)
           || (msg_type_trans_S1 == 8'd54)
           || (msg_type_trans_S1 == 8'd55)
           || (msg_type_trans_S1 == 8'd56)
           || (msg_type_trans_S1 == 8'd57)
           || (msg_type_trans_S1 == 8'd58)
           || (msg_type_trans_S1 == 8'd59)
           || (msg_type_trans_S1 == 8'd15))
           && !msg_from_mshr_S1)
    begin
        msg_input_en_S1_next = n;
    end
    else if ((valid_S2 && !stall_S2)
           &&((((msg_type_S2_f == 8'd7)
           || (msg_type_S2_f == 8'd11)
           || (msg_type_S2_f == 8'd52)
           || (msg_type_S2_f == 8'd53)
           || (msg_type_S2_f == 8'd54)
           || (msg_type_S2_f == 8'd55)
           || (msg_type_S2_f == 8'd56)
           || (msg_type_S2_f == 8'd57)
           || (msg_type_S2_f == 8'd58)
           || (msg_type_S2_f == 8'd59))
                && l2_tag_hit_S2 && (l2_way_state_mesi_S2 == 2'b00))
            ||((msg_type_S2_f == 8'd15)
                && ((!l2_tag_hit_S2 && !msg_from_mshr_S2_f) || (l2_tag_hit_S2 && (l2_way_state_mesi_S2 == 2'b00) && (l2_way_state_vd_S2 == 2'b10))))))
    begin
        msg_input_en_S1_next = y;
    end
    else
    begin
        msg_input_en_S1_next = msg_input_en_S1_f;
    end
end
always @ (posedge clk)
begin
    msg_input_en_S1_f <= msg_input_en_S1_next;
end
always @ *
begin
    msg_data_rd_S1 = valid_S1 && (msg_type_trans_S1 == 8'd15)
                  && (addr_type_S1 == 8'ha7
                  ||  addr_type_S1 == 8'ha9
                  ||  addr_type_S1 == 8'ha8
                  ||  addr_type_S1 == 8'haa
                  ||  addr_type_S1 == 8'hab
                  ||  addr_type_S1 == 8'ha4);
end
always @ *
begin
    reg_wr_en_S1 = valid_S1 && ~stall_S1 && (msg_type_trans_S1 == 8'd15)
               && ((addr_type_S1 == 8'ha9)
                || (addr_type_S1 == 8'ha7)
                || (addr_type_S1 == 8'ha8)
                || (addr_type_S1 == 8'haa)
                || (addr_type_S1 == 8'hab));
end
always @ *
begin
    reg_wr_addr_type_S1 = addr_type_S1;
end
always @ *
begin
    if (!rst_n)
    begin
        msg_cas_cmp_S1_next = n;
    end
    else if (msg_type_S4_f == 8'd6 && cas_cmp_en_S4)
    begin
        if (cas_cmp_S4)
        begin
            msg_cas_cmp_S1_next = y;
        end
        else
        begin
            msg_cas_cmp_S1_next = n;
        end
    end
    else
    begin
        msg_cas_cmp_S1_next = msg_cas_cmp_S1_f;
    end
end
always @ (posedge clk)
begin
    msg_cas_cmp_S1_f <= msg_cas_cmp_S1_next;
end
always @ *
begin
    stall_hazard_S1 = (valid_S2 && (addr_S1[6+8-1:6] == addr_S2[6+8-1:6]))
                   || (valid_S3 && (addr_S1[6+8-1:6] == addr_S3[6+8-1:6]))
                   || (valid_S4 && (addr_S1[6+8-1:6] == addr_S4[6+8-1:6]))
                   || (pipe2_valid_S1 && (addr_S1[39:6] == pipe2_addr_S1[39:6]))
                   || (pipe2_valid_S2 && (addr_S1[39:6] == pipe2_addr_S2[39:6]))
                   || (pipe2_valid_S3 && (addr_S1[39:6] == pipe2_addr_S3[39:6]));
end
reg stall_mshr_S1;
always @ *
begin
    
    
    stall_mshr_S1 = (mshr_cam_en_S1 && mshr_hit_S1)
                 || (~msg_from_mshr_S1
                 
                 &&((mshr_empty_slots_S1 <= 3 && (valid_S2 || valid_S3 || valid_S4))
                 ||  mshr_empty_slots_S1 == 0));
end
reg stall_msg_S1;
always @ *
begin
    stall_msg_S1 = msg_data_rd_S1 && ~msg_data_valid_S1;
end
always @ *
begin
    stall_S1 = valid_S1 && (stall_pre_S1 || stall_hazard_S1 || stall_mshr_S1 || stall_msg_S1);
end
always @ *
begin
    msg_header_ready_real_S1 = (!stall_S1) && (!msg_from_mshr_S1) && msg_input_en_S1_f;
end
always @ *
begin
    msg_header_ready_S1 = msg_header_ready_real_S1
        && ((msg_type_trans_S1 != 8'd6)
         && (msg_type_trans_S1 != 8'd10)
         && (msg_type_trans_S1 != 8'd44)
         && (msg_type_trans_S1 != 8'd45)
         && (msg_type_trans_S1 != 8'd46)
         && (msg_type_trans_S1 != 8'd47)
         && (msg_type_trans_S1 != 8'd48)
         && (msg_type_trans_S1 != 8'd49)
         && (msg_type_trans_S1 != 8'd50)
         && (msg_type_trans_S1 != 8'd51)
         );
end
always @ *
begin
    
    tag_clk_en_S1 = valid_S1 && cs_S1[2];
    
end
always @ *
begin
    
    tag_rdw_en_S1 = valid_S1 && cs_S1[1];
    
end
always @ *
begin
    
    state_rd_en_S1 = valid_S1 && cs_S1[0];
    
end
reg l2_miss_S1;
always @ *
begin
    if (msg_from_mshr_S1)
    begin
        l2_miss_S1 = pending_mshr_l2_miss_S1;
 
    end
    else
    begin
        l2_miss_S1 = 0;
    end
end
reg valid_S1_next;
always @ *
begin
    valid_S1_next = valid_S1 && !stall_S1;
end
reg valid_S2_f;
reg [3-1:0] data_size_S2_f;
reg [1-1:0] cache_type_S2_f;
reg [1-1:0] l2_miss_S2_f;
reg mshr_smc_miss_S2_f;
reg [3-1:0] mshr_pending_index_S2_f;
reg special_addr_type_S2_f;
reg msg_data_rd_S2_f;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        valid_S2_f <= 1'b0;
        msg_type_S2_f <= 0;
        data_size_S2_f <= 0;
        cache_type_S2_f <= 0;
        l2_miss_S2_f <= 0;
        
        mshr_smc_miss_S2_f <= 0;
        
        msg_from_mshr_S2_f <= 1'b0;
        mshr_pending_index_S2_f <= 0;
        special_addr_type_S2_f <= 0;
        msg_data_rd_S2_f <= 0;
        amo_alu_op_S2_f <= 4'b0;
    end
    else if (!stall_S2)
    begin
        valid_S2_f <= valid_S1_next;
        msg_type_S2_f <= msg_type_trans_S1;
        data_size_S2_f <= data_size_S1;
        cache_type_S2_f <= cache_type_S1;
        l2_miss_S2_f <= l2_miss_S1;
        
        mshr_smc_miss_S2_f <= (mshr_pending_S1 == 1'b1) ? pending_mshr_smc_miss_S1 : (mshr_hit_S1 && cam_mshr_smc_miss_S1);
 
        
        msg_from_mshr_S2_f <= msg_from_mshr_S1;
        mshr_pending_index_S2_f <= mshr_pending_index_S1;
        special_addr_type_S2_f <= special_addr_type_S1;
        msg_data_rd_S2_f <= msg_data_rd_S1;
        amo_alu_op_S2_f <= amo_alu_op_S1;
    end
end
reg stall_pre_S2;
reg stall_before_S2_f;
reg stall_before_S2_next;
reg state_wr_en_S2;
reg [1-1:0] l2_miss_S2;
reg req_recycle_S2;
reg req_recycle_cur_S2;
reg req_recycle_buf_S2_f;
reg req_recycle_buf_S2_next;
reg mshr_wr_data_en_S2;
reg mshr_wr_state_en_S2;
reg [2-1:0] mshr_state_in_S2;
reg [8-1:0] addr_type_S2;
reg [2-1:0] addr_op_S2;
always @ *
begin
    valid_S2 = valid_S2_f;
    data_size_S2 = data_size_S2_f;
    cache_type_S2 = cache_type_S2_f;
    msg_from_mshr_S2 = msg_from_mshr_S2_f;
    stall_before_S2 = stall_before_S2_f;
    msg_type_S2 = msg_type_S2_f;
    special_addr_type_S2 = special_addr_type_S2_f;
    amo_alu_op_S2 = amo_alu_op_S2_f;
end
always @ *
begin
    addr_type_S2 = addr_S2[39:32];
    addr_op_S2 = addr_S2[31:30];
end
always @ *
begin
    if (!rst_n)
    begin
        stall_before_S2_next = 0;
    end
    else
    begin
        stall_before_S2_next = stall_S2;
    end
end
always @ (posedge clk)
begin
    stall_before_S2_f <= stall_before_S2_next;
end
always @ *
begin
    stall_pre_S2 = stall_S3 || global_stall_S2;
end
reg [27-1:0] cs_S2;
always @ *
begin
    
    cs_S2 = {27{1'bx}};
    if (valid_S2)
    begin
        if (special_addr_type_S2_f)
        begin
            case (addr_type_S2)
                8'ha0:
                begin
                    if (msg_type_S2_f == 8'd14)
                    begin
                        
                        
                        cs_S2 = {4'd0, n,         rd,      2'd0, y,      rd,            n,       n,         2'd0,     n,          n,
                        
                        
                                 2'd0,    n,      n,      2'b01,  n,       2'b00, n,      1'b0};
                    end
                    else
                    begin
                        cs_S2 = {4'd0, n,         rd,      2'd0, y,      wr,            n,       n,         2'd0,     n,          y,
                                 2'd0,    n,      n,      2'b01,  n,       2'b00, n,      1'b0};
                    end
                end
                8'ha1:
                begin
                    if (msg_type_S2_f == 8'd14)
                    begin
                        cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            n,       n,         2'd0,     n,          n,
                                 2'd0,    n,      n,      2'b01,  n,       2'b00, n,      1'b0};
                    end
                    else
                    begin
                        cs_S2 = {4'd0, y,         wr,      2'd0, n,      rd,            n,       n,         2'd0,     n,          y,
                                 2'd0,    n,      n,      2'b01,  n,       2'b00, n,      1'b0};
                    end
                end
                8'ha6:
                begin
                    if (msg_type_S2_f == 8'd15)
                    begin
                        cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            n,       y,         2'd0,     y,          y,
                                 2'd0,    y,      y,      2'b00,  y,       2'b00, y,      1'b0};
                    end
                    else
                    begin
                        cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            n,       n,         2'd0,     n,          n,
                                 2'd0,    n,      n,      2'b01,  n,       2'b00, n,      1'b0};
                    end
                end
                8'ha2:
                begin
                    if (msg_type_S2_f == 8'd15)
                    begin
                        cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            n,       n,         2'd0,     n,          y,
                                 2'd0,    n,      n,      2'b01,  n,       2'b00, n,      1'b0};
                    end
                    else
                    begin
                        cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            n,       n,         2'd0,     n,          n,
                                 2'd0,    n,      n,      2'b01,  n,       2'b00, n,      1'b0};
                    end
                end
                default:
                begin
                    cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            n,       n,         2'd0,     n,          n,
                             2'd0,    n,      n,      2'b01,  n,       2'b00, n,      1'b0};
                end
            endcase
        end
        else if (req_recycle_S2)
        begin
            cs_S2 = {27{1'b0}};
        end
        else
        begin
            if ((msg_type_S2_f == 8'd8) || (msg_type_S2_f == 8'd32))
            begin
                cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            n,       n,         2'd0,     n,          y,
                         2'd0,    n,      n,      2'b01,  n,       2'b00, n,      1'b0};
            end
            else if (l2_evict_S2)
            begin
                case (l2_way_state_mesi_S2)
                2'b01:
                begin
                    cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,          n,
                             2'd0,   n,       n,      2'b01,  n,      2'b00, n,      1'b0};
                end
                
                2'b11:
                begin
                    cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,          n,
                             2'd0,   n,       n,      2'b01,  n,      2'b00, n,      1'b0};
                end
                
                2'b10:
                begin
                    
                    if (csm_en)
                    begin
                        cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,          n,
                                 2'd0,   n,       n,      2'b01,  n,      2'b00, n,      1'b0};
                    end
                    else
                    
                    begin
                        cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,          n,
                                 2'd0,   n,       n,      2'b01,  n,      2'b00, n,      1'b0};
                    end
                end
                2'b00:
                begin
                    case (l2_way_state_vd_S2)
                    2'b10:
                    begin
                        if (msg_type_S2_f == 8'd34)
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            n,       n,         2'd0,    n,          n,
                                    2'd0,   n,       y,      2'b00,  n,      2'b00, y,      1'b0};
                        end
                        else
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,          n,
                                    2'd0,   n,       y,      2'b00,  n,      2'b00, y,      1'b0};
                        end
                    end
                    2'b11:
                    begin
                        if (msg_type_S2_f == 8'd34)
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, y,      rd,            n,       n,         2'd0,    n,          n,
                                    2'd0,   n,       y,      2'b00,  n,      2'b00, y,      1'b0};
                        end
                        else
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, y,      rd,            y,       n,         2'd0,    n,          n,
                                     2'd0,   n,       y,      2'b00,  n,      2'b00, y,      1'b0};
                        end
                    end
                    default:
                    begin
                        cs_S2 = {27{1'bx}};
                    end
                    endcase
                end
                default:
                begin
                    cs_S2 = {27{1'bx}};
                end
                endcase
            end
            else if (!l2_tag_hit_S2)
            begin
                if (msg_type_S2_f == 8'd15)
                begin
                    if (msg_from_mshr_S2_f)
                    begin
                        
                        
                        cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            n,       n,         2'd0,     n,          n,
                        
                        
                                 2'd0,    n,      n,      2'b01,  n,       2'b00, n,      1'b0};
                    end
                    else
                    begin
                        cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,     n,          y,
                                 2'd0,    n,      n,      2'b01,  n,       2'b00, n,      1'b0};
                    end
                end
                else if (msg_type_S2_f == 8'd13
                 || msg_type_S2_f == 8'd34
                 || msg_type_S2_f == 8'd35)
                begin
                    cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            n,       n,         2'd0,    n,          n,
                             2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                end
                else
                begin
                    cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,          n,
                             2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                end
            end
            else begin
            case (msg_type_S2_f)
                8'd13:
                begin
                    
                    if (csm_en && (l2_way_state_mesi_S2 == 2'b10) && l2_way_state_subline_S2[addr_S2[5:4]])
                    begin
                        cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            n,       n,         2'd0,    n,          n,
                                2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                    end
                    else
                    
                    begin
                        cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            n,       n,         2'd0,    n,          n,
                                2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                    end
                end
                8'd35:
                begin
                    case (l2_way_state_mesi_S2)
                    2'b00:
                    begin
                        cs_S2 = {4'd0, n,         rd,      2'd0, y,      rd,            n,       n,         2'd0,    n,          n,
                                2'd0,   n,       y,      2'b00,  n,      2'b00, y,      1'b0};
                    end
                    2'b01:
                    begin
                        cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                 2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                    end
                    
                    2'b11:
                    begin
                        cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                 2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                    end
                    
                    2'b10:
                    begin
                        
                        if (csm_en)
                        begin
                            cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                     2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                        end
                        else
                        
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                     2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                        end
                    end
                    default:
                    begin
                        cs_S2 = {27{1'bx}};
                    end
                    endcase
                end
                8'd14:
                begin
                    case (l2_way_state_mesi_S2)
                    2'b00:
                    begin
                        case (l2_way_state_vd_S2)
                        2'b10:
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, y,      rd,            n,       n,         2'd0,    n,          n,
                                    2'd0,   n,       y,      2'b00,  n,      2'b00, y,      1'b0};
                        end
                        2'b11:
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, y,      rd,            y,       n,         2'd0,    n,          n,
                                    2'd0,   n,       y,      2'b10,  n,      2'b00, y,      1'b0};
                        end
                        default:
                        begin
                            cs_S2 = {27{1'bx}};
                        end
                        endcase
                    end
                    2'b01:
                    begin
                        cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                 2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                    end
                    
                    2'b11:
                    begin
                        cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                 2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                    end
                    
                    2'b10:
                    begin
                        
                        if (csm_en)
                        begin
                            cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                     2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                        end
                        else
                        
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                     2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                        end
                    end
                    default:
                    begin
                        cs_S2 = {27{1'bx}};
                    end
                    endcase
                end
                8'd15:
                begin
                    case (l2_way_state_mesi_S2)
                    2'b00:
                    begin
                        case (l2_way_state_vd_S2)
                        2'b10:
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, y,      rd,            y,       n,         2'd0,    n,          y,
                                    2'd0,   n,       y,      2'b00,  n,      2'b00, y,      1'b0};
                        end
                        2'b11:
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, y,      rd,            y,       n,         2'd0,    n,          n,
                                    2'd0,   n,       y,      2'b10,  n,      2'b00, y,      1'b0};
                        end
                        default:
                        begin
                            cs_S2 = {27{1'bx}};
                        end
                        endcase
                    end
                    2'b01:
                    begin
                        cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                 2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                    end
                    
                    2'b11:
                    begin
                        cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                 2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                    end
                    
                    2'b10:
                    begin
                        
                        if (csm_en)
                        begin
                            cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                     2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                        end
                        else
                        
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                     2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                        end
                    end
                    default:
                    begin
                        cs_S2 = {27{1'bx}};
                    end
                    endcase
                end
                8'd31:
                begin
                    case (l2_way_state_mesi_S2)
                    2'b00:
                    begin
                        if (cache_type_S2_f == 1'b0)
                        begin
                            
                            if (csm_en)
                            begin
                                cs_S2 = {4'd0, y,         wr,      2'd1, y,      rd,            n,       y,         2'd1,     y,      n,
                                         2'd2,   y,       n,      2'b00,  y,      2'b10,   y,     1'b1};
                            end
                            else
                            
                            begin
                                cs_S2 = {4'd0, n,         rd,      2'd0, y,      rd,            n,       y,         2'd1,     y,      n,
                                         2'd2,   y,       n,      2'b00,  y,      2'b10,   y,     1'b1};
                            end
                        end
                        else
                        begin
                            
                            if (csm_en)
                            begin
                                if (lsid_S2 == 6'd63)
                                begin
                                    cs_S2 = {4'd0, y,         wr,      2'd0, y,      rd,            n,       y,         2'd0,     y,      n,
                                            2'd1,   y,       n,      2'b00,  y,      2'b11,   y,     1'b1};
                                end
                                else
                                begin
                                    cs_S2 = {4'd0, y,         wr,      2'd0, y,      rd,            n,       y,         2'd1,     y,      n,
                                            2'd1,   y,       n,      2'b00,  y,      2'b01,   y,     1'b1};
                                end
                            end
                            else
                            
                            begin
                                cs_S2 = {4'd0, y,         wr,      2'd0, y,      rd,            n,       y,         2'd0,     y,      n,
                                         2'd2,   y,       n,      2'b00,  y,      2'b01,   y,     1'b1};
                            end
                        end
                    end
                    2'b01:
                    begin
                        if (cache_type_S2_f == l2_way_state_cache_type_S2)
                        begin
                            
                            if (csm_en)
                            begin
                                cs_S2 = {4'd0, y,         wr,      2'd0, y,      rd,            n,       n,         2'd0,    n,      n,
                                        2'd0,   n,       n,      2'b00,  n,      2'b00, y,     1'b1};
                            end
                            else
                            
                            begin
                                cs_S2 = {4'd0, y,         wr,      2'd0, y,      rd,            n,       n,         2'd0,    y,      n,
                                        2'd2,   n,       n,      2'b00,  n,      2'b00, y,     1'b1};
                            end
                        end
                        else
                        begin
                            cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                     2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                        end
                    end
                    
                    2'b11:
                    begin
                        if (cache_type_S2_f == l2_way_state_cache_type_S2)
                        begin
                            
                            if (csm_en)
                            begin
                                cs_S2 = {4'd0, n,         wr,      2'd0, y,      rd,            n,       n,         2'd0,    n,      n,
                                         2'd0,   n,       n,      2'b00,  n,      2'b00, y,     1'b1};
                            end
                            else
                            
                            begin
                                cs_S2 = {4'd0, n,         wr,      2'd0, y,      rd,            n,       n,         2'd0,    y,      n,
                                         2'd2,   n,       n,      2'b00,  n,      2'b00, y,     1'b1};
                            end
                        end
                        else
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                     2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                        end
                    end
                    
                    2'b10:
                    begin
                        if (req_from_owner_S2 && (cache_type_S2_f == l2_way_state_cache_type_S2))
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, y,      rd,            n,       n,         2'd0,    y,      n,
                                     2'd2,   n,       n,      2'b00,  n,      2'b00, y,      1'b1};
                        end
                        else
                        begin
                            
                            if (csm_en)
                            begin
                                cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                         2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                            end
                            else
                            
                            begin
                                cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                         2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                            end
                        end
                    end
                    default:
                    begin
                        cs_S2 = {27{1'bx}};
                    end
                    endcase
                end
                
                8'd60:
                begin
                    case (l2_way_state_mesi_S2)
                    2'b00:
                    begin
                        if (cache_type_S2_f == 1'b0)
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, y,      rd,            n,       y,         2'd1,     y,      n,
                                     2'd2,   y,       n,      2'b00,  y,      2'b10,   y,     1'b1};
                        end
                        else begin
                            cs_S2 = {27{1'bx}};
                        end
                    end
                    2'b01:   
                    begin
                        cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,          n,
                                 2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                    end
                    2'b10:
                    begin
                        if (req_from_owner_S2 && (cache_type_S2_f == l2_way_state_cache_type_S2))
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, y,      rd,            n,       n,         2'd0,    y,      n,
                                     2'd2,   n,       n,      2'b00,  n,      2'b00, y,      1'b1};
                        end
                        else
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                     2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                        end
                    end
                    default:
                    begin
                        cs_S2 = {27{1'bx}};
                    end
                    endcase
                end
                8'd1:
                begin
                    cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            n,       n,         2'd0,    n,      n,
                             2'd0,   n,       n,      2'b00,  n,      2'b00, y,      1'b1};
                end
                8'd2:
                begin
                    case (l2_way_state_mesi_S2)
                    2'b00:
                    begin
                        
                        if (csm_en)
                        begin
                            cs_S2 = {4'd0, y,         wr,      2'd1, y,      rd,            n,       y,         2'd1,     y,      n,
                                     2'd2,   y,       n,      2'b00,  y,      2'b10, y,     1'b1};
                        end
                        else
                        
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, y,      rd,            n,       y,         2'd1,     y,      n,
                                     2'd2,   y,       n,      2'b00,  y,      2'b10, y,     1'b1};
                        end
                    end
                    2'b01:
                    begin
                        cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,          n,
                                 2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                    end
                    
                    2'b11:
                    begin
                        cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,          n,
                                 2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                    end
                    
                    2'b10:
                    begin
                        if (req_from_owner_S2 && (cache_type_S2_f == l2_way_state_cache_type_S2))
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, y,      rd,            n,       n,         2'd0,    y,      n,
                                     2'd2,   n,       n,      2'b00,  n,      2'b00, y,      1'b1};
                        end
                        else
                        begin
                            
                            if (csm_en)
                            begin
                                cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                         2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                            end
                            else
                            
                            begin
                                cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                         2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                            end
                        end
                    end
                    default:
                    begin
                        cs_S2 = {27{1'bx}};
                    end
                    endcase
                end
                8'd6:
                begin
                    case (l2_way_state_mesi_S2)
                    2'b00:
                    begin
                        cs_S2 = {4'd0, n,         rd,      2'd0, y,      rd,            n,       n,         2'd0,     n,      y,
                                 2'd0,   n,       n,      2'b00,  n,      2'b00,   y,     1'b1};
                    end
                    2'b01:
                    begin
                        cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                 2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                    end
                    
                    2'b11:
                    begin
                        cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                 2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                    end
                    
                    2'b10:
                    begin
                        
                        if (csm_en)
                        begin
                            cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                     2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                        end
                        else
                        
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                     2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                        end
                    end
                    default:
                    begin
                        cs_S2 = {27{1'bx}};
                    end
                    endcase
                end
                8'd10,
                8'd44,
                8'd45,
                8'd46,
                8'd47,
                8'd48,
                8'd49,
                8'd50,
                8'd51:
                begin
                    case (l2_way_state_mesi_S2)
                    2'b00:
                    begin
                        cs_S2 = {4'd0, n,         rd,      2'd0, y,      rd,            n,       n,         2'd0,     n,      n,
                                 2'd0,   n,       n,      2'b00,  n,      2'b00,   y,     1'b1};
                    end
                    2'b01:
                    begin
                        cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                 2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                    end
                    
                    2'b11:
                    begin
                        cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                 2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                    end
                    
                    2'b10:
                    begin
                        
                        if (csm_en)
                        begin
                            cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                     2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                        end
                        else
                        
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                     2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                        end
                    end
                    default:
                    begin
                        cs_S2 = {27{1'bx}};
                    end
                    endcase
                end
                8'd7,
                8'd11,
                8'd52,
                8'd53,
                8'd54,
                8'd55,
                8'd56,
                8'd57,
                8'd58,
                8'd59:
                begin
                    case (l2_way_state_mesi_S2)
                    2'b00:
                    begin
                        case (msg_type_S2_f)
                        8'd7,
                        8'd11:
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, y,      wr,            n,       n,         2'd0,    n,      y,
                                 2'd0,   y,       y,      2'b11,  n,      2'b00, y,      1'b1};
                        end
                        8'd52:
                        begin
                            cs_S2 = {4'd1, n,         rd,      2'd0, y,      wr,            n,       n,         2'd0,    n,      y,
                                 2'd0,   y,       y,      2'b11,  n,      2'b00, y,      1'b1};
                        end
                        8'd53:
                        begin
                            cs_S2 = {4'd2, n,         rd,      2'd0, y,      wr,            n,       n,         2'd0,    n,      y,
                                 2'd0,   y,       y,      2'b11,  n,      2'b00, y,      1'b1};
                        end
                        8'd54:
                        begin
                            cs_S2 = {4'd3, n,         rd,      2'd0, y,      wr,            n,       n,         2'd0,    n,      y,
                                 2'd0,   y,       y,      2'b11,  n,      2'b00, y,      1'b1};
                        end
                        8'd55:
                        begin
                            cs_S2 = {4'd4, n,         rd,      2'd0, y,      wr,            n,       n,         2'd0,    n,      y,
                                 2'd0,   y,       y,      2'b11,  n,      2'b00, y,      1'b1};
                        end
                        8'd56:
                        begin
                            cs_S2 = {4'd5, n,         rd,      2'd0, y,      wr,            n,       n,         2'd0,    n,      y,
                                 2'd0,   y,       y,      2'b11,  n,      2'b00, y,      1'b1};
                        end
                        8'd57:
                        begin
                            cs_S2 = {4'd6, n,         rd,      2'd0, y,      wr,            n,       n,         2'd0,    n,      y,
                                 2'd0,   y,       y,      2'b11,  n,      2'b00, y,      1'b1};
                        end
                        8'd58:
                        begin
                            cs_S2 = {4'd7, n,         rd,      2'd0, y,      wr,            n,       n,         2'd0,    n,      y,
                                 2'd0,   y,       y,      2'b11,  n,      2'b00, y,      1'b1};
                        end
                        8'd59:
                        begin
                            cs_S2 = {4'd8, n,         rd,      2'd0, y,      wr,            n,       n,         2'd0,    n,      y,
                                 2'd0,   y,       y,      2'b11,  n,      2'b00, y,      1'b1};
                        end
                        endcase
                    end
                    2'b01:
                    begin
                        cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                 2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                    end
                    
                    2'b11:
                    begin
                        cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                 2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                    end
                    
                    2'b10:
                    begin
                        
                        if (csm_en)
                        begin
                            cs_S2 = {4'd0, y,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                     2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                        end
                        else
                        
                        begin
                            cs_S2 = {4'd0, n,         rd,      2'd0, n,      rd,            y,       n,         2'd0,    n,      n,
                                     2'd0,   n,       n,      2'b00,  n,      2'b00, n,      1'b0};
                        end
                    end
                    default:
                    begin
                        cs_S2 = {27{1'bx}};
                    end
                    endcase
                end
                default:
                begin
                    cs_S2 = {27{1'bx}};
                end
            endcase
            end
        end
    end
    else
    begin
        cs_S2 = {27{1'b0}};
    end
end
reg [2-1:0] l2_load_data_subline_S2_f;
reg [2-1:0] l2_load_data_subline_S2_next;
always @ *
begin
    dir_clk_en_S2 = !stall_S2 && cs_S2[22];
end
always @ *
begin
    dir_rdw_en_S2 = !stall_S2 && cs_S2[21];
end
always @ *
begin
    dir_op_S2 = cs_S2[20:19];
end
always @ *
begin
    data_clk_en_S2 = !stall_real_S2 && cs_S2[18];
end
always @ *
begin
    data_rdw_en_S2 = !stall_real_S2 && cs_S2[17];
end
always @ *
begin
    mshr_wr_data_en_S2 = !stall_S2 && cs_S2[16];
    mshr_wr_state_en_S2 = !stall_S2 && cs_S2[16];
end
always @ *
begin
    if ( l2_tag_hit_S2 && (msg_type_S2_f == 8'd14 || msg_type_S2_f == 8'd15)
    && (l2_way_state_mesi_S2 == 2'b00) && (l2_way_state_vd_S2 == 2'b11))
    begin
        mshr_state_in_S2 = 2'd2;
    end
    else
    begin
        mshr_state_in_S2 = 2'd1;
    end
end
always @ *
begin
    if (!l2_tag_hit_S2)
    begin
        l2_miss_S2 = 1;
    end
    else
    begin
        l2_miss_S2 = l2_miss_S2_f;
    end
end
always @ *
begin
    if (special_addr_type_S2_f && (addr_type_S2 == 8'ha2) && (msg_type_S2_f == 8'd15))
    begin
        smc_wr_en_S2 = 1'b1;
        smc_wr_diag_en_S2 = 1'b1;
    end
    else
    begin
        smc_wr_en_S2 = 1'b0;
        smc_wr_diag_en_S2 = 1'b0;
    end
end
always @ *
begin
    if (special_addr_type_S2_f && (addr_type_S2 == 8'ha5))
    begin
        smc_flush_en_S2 = 1'b1;
    end
    else
    begin
        smc_flush_en_S2 = 1'b0;
    end
end
always @ *
begin
    smc_addr_op_S2 = addr_op_S2;
end
always @ *
begin
    state_owner_en_S2 =  cs_S2[15];
end
always @ *
begin
    state_owner_op_S2 = cs_S2[14:13];
end
always @ *
begin
    state_subline_en_S2 =  cs_S2[12];
end
always @ *
begin
    state_subline_op_S2 = cs_S2[10:9];
end
assign state_load_sdid_S2 = csm_en && state_owner_en_S2 && (state_owner_op_S2 ==2'd1)
                                && state_subline_en_S2 && (state_subline_op_S2 == 2'd1);
always @ *
begin
    state_di_en_S2 = cs_S2[8];
end
always @ *
begin
    state_vd_en_S2 = cs_S2[7];
end
always @ *
begin
    state_vd_S2 = cs_S2[6:5];
end
always @ *
begin
    state_mesi_en_S2 = cs_S2[4];
end
always @ *
begin
    if (!cs_S2[4])
    begin
        state_mesi_S2 = l2_way_state_mesi_S2;
    end
    else
    begin
        state_mesi_S2 = cs_S2[3:2];
    end
end
always @ *
begin
    state_lru_en_S2 =  cs_S2[1];
end
always @ *
begin
    state_lru_op_S2 = cs_S2[0];
end
always @ *
begin
    state_rb_en_S2 =  l2_evict_S2  && (l2_way_state_mesi_S2 == 2'b00)
                 && (msg_type_S2_f != 8'd8);
end
always @ *
begin
    state_wr_en_S2 = valid_S2 && !stall_S2 && (
                          cs_S2[15]
                       || cs_S2[12]
                       || cs_S2[7]
                       || cs_S2[8]
                       || cs_S2[4]
                       || cs_S2[1]
                       || (state_rb_en_S2));
end
always @ *
begin
    req_recycle_cur_S2 = valid_S2
    &&  (~special_addr_type_S2_f)
    &&  ((pipe2_valid_S1 && (pipe2_msg_type_S1 == 8'd12)
        && (addr_S2[39:6] == pipe2_addr_S1[39:6]))
    ||   (pipe2_valid_S2 && (pipe2_msg_type_S1 == 8'd12)
        && (addr_S2[39:6] == pipe2_addr_S2[39:6]))
    ||   (pipe2_valid_S3 && (pipe2_msg_type_S3 == 8'd12)
        && (addr_S2[39:6] == pipe2_addr_S3[39:6])));
end
always @ *
begin
    if (!rst_n)
    begin
        req_recycle_buf_S2_next = 1'b0;
    end
    else
    begin
        if (!stall_S2)
        begin
            req_recycle_buf_S2_next = 1'b0;
        end
        else if (req_recycle_cur_S2)
        begin
            req_recycle_buf_S2_next = 1'b1;
        end
        else
        begin
            req_recycle_buf_S2_next = req_recycle_buf_S2_f;
        end
    end
end
always @ (posedge clk)
begin
    req_recycle_buf_S2_f <= req_recycle_buf_S2_next;
end
always @ *
begin
    req_recycle_S2 = req_recycle_cur_S2 | req_recycle_buf_S2_f;
end
always @ *
begin
    msg_data_ready_S2 = valid_S2 && !stall_S2 && (cs_S2[11] || msg_data_rd_S2_f);
end
always @ *
begin
    if (special_addr_type_S2)
    begin
        l2_ifill_32B_S2 = n;
    end
    else if (valid_S2 && l2_tag_hit_S2 && data_clk_en_S2 && (data_rdw_en_S2 == rd) && ~l2_wb_S2
    && (cache_type_S2_f == 1'b1))
    begin
        l2_ifill_32B_S2 = y;
    end
    else
    begin
        l2_ifill_32B_S2 = n;
    end
end
always @ *
begin
    if (!rst_n)
    begin
        l2_load_data_subline_S2_next = 2'd0;
    end
    else if (valid_S2 && !(stall_real_S2) && l2_ifill_32B_S2 && (l2_load_data_subline_S2_f == 2'd1))
    begin
        l2_load_data_subline_S2_next = 2'd0;
    end
    else if (valid_S2 && !(stall_real_S2) && (l2_wb_S2 || l2_ifill_32B_S2))
    begin
        l2_load_data_subline_S2_next = l2_load_data_subline_S2_f + 1;
    end
    else
    begin
        l2_load_data_subline_S2_next = l2_load_data_subline_S2_f;
    end
end
always @ (posedge clk)
begin
    l2_load_data_subline_S2_f <= l2_load_data_subline_S2_next;
end
reg stall_load_S2;
always @ *
begin
    if (l2_wb_S2)
    begin
        stall_load_S2 = (l2_load_data_subline_S2_f != 2'd3);
    end
    else if (l2_ifill_32B_S2)
    begin
        stall_load_S2 = (l2_load_data_subline_S2_f != 2'd1);
    end
    else
    begin
        stall_load_S2 = n;
    end
end
always @ *
begin
    l2_load_data_subline_S2 = l2_load_data_subline_S2_f;
end
reg stall_msg_S2;
always @ *
begin
    stall_msg_S2 = (cs_S2[11] || msg_data_rd_S2_f) && ~msg_data_valid_S2;
end
always @ *
begin
    stall_real_S2 = valid_S2 && (stall_pre_S2 || stall_msg_S2);
 end
always @ *
begin
    stall_S2 = valid_S2 && (stall_real_S2 || stall_load_S2);
end
reg valid_S2_next;
always @ *
begin
    valid_S2_next = valid_S2 && !stall_real_S2;
end
reg valid_S3_f;
reg [8-1:0] msg_type_S3_f;
reg [3-1:0] data_size_S3_f;
reg [1-1:0] cache_type_S3_f;
reg msg_from_mshr_S3_f;
reg [2-1:0] l2_load_data_subline_S3_f;
reg [2-1:0] state_mesi_S3_f;
reg [1-1:0] l2_miss_S3_f;
reg mshr_smc_miss_S3_f;
reg state_wr_en_S3_f;
reg mshr_wr_data_en_S3_f;
reg mshr_wr_state_en_S3_f;
reg [2-1:0] mshr_state_in_S3_f;
reg [3-1:0] mshr_pending_index_S3_f;
reg special_addr_type_S3_f;
reg req_recycle_S3_f;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        valid_S3_f <= 1'b0;
        msg_type_S3_f <= 0;
        data_size_S3_f <= 0;
        cache_type_S3_f <= 0;
        msg_from_mshr_S3_f <= 0;
        l2_load_data_subline_S3_f <= 0;
        state_mesi_S3_f <= 0;
        l2_miss_S3_f <= 0;
        
        mshr_smc_miss_S3_f <= 0;
        
        state_wr_en_S3_f <= 0;
        mshr_wr_data_en_S3_f <= 0;
        mshr_wr_state_en_S3_f <= 0;
        mshr_state_in_S3_f <= 0;
        mshr_pending_index_S3_f <= 0;
        special_addr_type_S3_f <= 0;
        req_recycle_S3_f <= 0;
    end
    else if (!stall_S3)
    begin
        valid_S3_f <= valid_S2_next;
        msg_type_S3_f <= msg_type_S2_f;
        data_size_S3_f <= data_size_S2_f;
        cache_type_S3_f <= cache_type_S2_f;
        msg_from_mshr_S3_f <= msg_from_mshr_S2_f;
        l2_load_data_subline_S3_f <= l2_load_data_subline_S2_f;
        state_mesi_S3_f <= state_mesi_S2;
        l2_miss_S3_f <= l2_miss_S2;
        
        mshr_smc_miss_S3_f <= mshr_smc_miss_S2_f;
        
        state_wr_en_S3_f <= state_wr_en_S2;
        mshr_wr_data_en_S3_f <= mshr_wr_data_en_S2;
        mshr_wr_state_en_S3_f <= mshr_wr_state_en_S2;
        mshr_state_in_S3_f <= mshr_state_in_S2;
        mshr_pending_index_S3_f <= mshr_pending_index_S2_f;
        special_addr_type_S3_f <= special_addr_type_S2_f;
        req_recycle_S3_f <= req_recycle_S2;
    end
end
reg stall_pre_S3;
reg stall_before_S3_f;
reg stall_before_S3_next;
reg req_recycle_S3;
reg req_recycle_cur_S3;
reg req_recycle_buf_S3_f;
reg req_recycle_buf_S3_next;
always @ *
begin
    stall_before_S3 = stall_before_S3_f;
    valid_S3 = valid_S3_f;
end
always @ *
begin
    req_recycle_cur_S3 = valid_S3 && (req_recycle_S3_f
     || (state_wr_en_S3_f
        && ((pipe2_valid_S1 && (pipe2_msg_type_S1 == 8'd12)
            && (addr_S3[39:6] == pipe2_addr_S1[39:6]))
        ||  (pipe2_valid_S2 && (pipe2_msg_type_S2 == 8'd12)
            && (addr_S3[39:6] == pipe2_addr_S2[39:6]))
        ||  (pipe2_valid_S3 && (pipe2_msg_type_S3 == 8'd12)
            && (addr_S3[39:6] == pipe2_addr_S3[39:6])))));
end
always @ *
begin
    if (!rst_n)
    begin
        req_recycle_buf_S3_next = 1'b0;
    end
    else
    begin
        if (!stall_S3)
        begin
            req_recycle_buf_S3_next = 1'b0;
        end
        else if (req_recycle_cur_S3)
        begin
            req_recycle_buf_S3_next = 1'b1;
        end
        else
        begin
            req_recycle_buf_S3_next = req_recycle_buf_S3_f;
        end
    end
end
always @ (posedge clk)
begin
    req_recycle_buf_S3_f <= req_recycle_buf_S3_next;
end
always @ *
begin
    req_recycle_S3 = req_recycle_cur_S3 | req_recycle_buf_S3_f;
end
always @ *
begin
    stall_pre_S3 = stall_S4;
    
end
always @ *
begin
    if (!rst_n)
    begin
        stall_before_S3_next = 0;
    end
    else
    begin
        stall_before_S3_next = stall_S3;
    end
end
always @ (posedge clk)
begin
    stall_before_S3_f <= stall_before_S3_next;
end
always @ *
begin
    stall_S3 = stall_pre_S3;
end
reg valid_S3_next;
always @ *
begin
    valid_S3_next = valid_S3 && !stall_S3;
end
reg valid_S4_f;
reg [3-1:0] data_size_S4_f;
reg [1-1:0] cache_type_S4_f;
reg msg_from_mshr_S4_f;
reg [2-1:0] l2_load_data_subline_S4_f;
reg [2-1:0] state_mesi_S4_f;
reg [1-1:0] l2_miss_S4_f;
reg mshr_smc_miss_S4_f;
reg state_wr_en_S4_f;
reg mshr_wr_data_en_S4_f;
reg mshr_wr_state_en_S4_f;
reg [2-1:0] mshr_state_in_S4_f;
reg [3-1:0] mshr_pending_index_S4_f;
reg special_addr_type_S4_f;
reg [64-1:0] dir_data_S4_f;
reg req_recycle_S4_f;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        valid_S4_f <= 1'b0;
        msg_type_S4_f <= 0;
        data_size_S4_f <= 0;
        cache_type_S4_f <= 0;
        msg_from_mshr_S4_f <= 0;
        l2_load_data_subline_S4_f <= 0;
        state_mesi_S4_f <= 0;
        l2_miss_S4_f <= 0;
        
        mshr_smc_miss_S4_f <= 0;
        
        state_wr_en_S4_f <= 0;
        mshr_wr_data_en_S4_f <= 0;
        mshr_wr_state_en_S4_f <= 0;
        mshr_state_in_S4_f <= 0;
        mshr_pending_index_S4_f <= 0;
        special_addr_type_S4_f <= 0;
        dir_data_S4_f <= 0;
        req_recycle_S4_f <= 0;
    end
    else if (!stall_S4)
    begin
        valid_S4_f <= valid_S3_next;
        msg_type_S4_f <= msg_type_S3_f;
        data_size_S4_f <= data_size_S3_f;
        cache_type_S4_f <= cache_type_S3_f;
        msg_from_mshr_S4_f <= msg_from_mshr_S3_f;
        l2_load_data_subline_S4_f <= l2_load_data_subline_S3_f;
        state_mesi_S4_f <= state_mesi_S3_f;
        l2_miss_S4_f <= l2_miss_S3_f;
        
        mshr_smc_miss_S4_f <= mshr_smc_miss_S3_f;
        
        state_wr_en_S4_f <= state_wr_en_S3_f;
        mshr_wr_data_en_S4_f <= mshr_wr_data_en_S3_f;
        mshr_wr_state_en_S4_f <= mshr_wr_state_en_S3_f;
        mshr_state_in_S4_f <= mshr_state_in_S3_f;
        mshr_pending_index_S4_f <= mshr_pending_index_S3_f;
        special_addr_type_S4_f <= special_addr_type_S3_f;
        dir_data_S4_f <= dir_data_S3;
        req_recycle_S4_f <= req_recycle_S3;
    end
end
reg stall_before_S4_f;
reg stall_before_S4_next;
reg dir_data_stall_S4;
reg state_wr_en_real_S4;
reg stall_inv_counter_S4;
reg msg_stall_S4;
reg load_store_mem_S4;
reg smc_stall_S4;
reg broadcast_stall_S4;
reg req_recycle_cur_S4;
reg req_recycle_buf_S4_f;
reg req_recycle_buf_S4_next;
reg [8-1:0] addr_type_S4;
reg [2-1:0] addr_op_S4;
reg msg0_send_valid_S4;
reg [8-1:0] msg0_send_type_S4;
reg msg1_send_valid_S4;
reg [8-1:0] msg1_send_type_S4;
reg smc_rd_diag_en_S4;
reg smc_rd_en_S4;
reg mshr_inv_flag_S4;
always @ *
begin
    valid_S4 = valid_S4_f;
    stall_before_S4 = stall_before_S4_f;
    msg_type_S4 = msg_type_S4_f;
    data_size_S4 = data_size_S4_f;
    cache_type_S4 = cache_type_S4_f;
    l2_miss_S4 = l2_miss_S4_f;
    special_addr_type_S4 = special_addr_type_S4_f;
    dir_data_S4 = dir_data_S4_f;
    msg_from_mshr_S4 = msg_from_mshr_S4_f;
end
always @ *
begin
    if (~special_addr_type_S4_f && req_recycle_S4)
    begin
        mshr_state_in_S4 = 2'd2;
    end
    else if(mshr_inv_flag_S4)
    begin
        mshr_state_in_S4 = 2'd0;
    end
    else
    begin
        mshr_state_in_S4 = mshr_state_in_S4_f;
    end
end
always @ *
begin
    req_recycle_cur_S4 = valid_S4 && (req_recycle_S4_f
     || (state_wr_en_S4_f
        && ((pipe2_valid_S1 && (pipe2_msg_type_S1 == 8'd12)
            && (addr_S4[39:6] == pipe2_addr_S1[39:6]))
        ||  (pipe2_valid_S2 && (pipe2_msg_type_S2 == 8'd12)
            && (addr_S4[39:6] == pipe2_addr_S2[39:6]))
        ||  (pipe2_valid_S3 && (pipe2_msg_type_S3 == 8'd12)
            && (addr_S4[39:6] == pipe2_addr_S3[39:6])))));
end
always @ *
begin
    if (!rst_n)
    begin
        req_recycle_buf_S4_next = 1'b0;
    end
    else
    begin
        if (!stall_S4)
        begin
            req_recycle_buf_S4_next = 1'b0;
        end
        else if (req_recycle_cur_S4)
        begin
            req_recycle_buf_S4_next = 1'b1;
        end
        else
        begin
            req_recycle_buf_S4_next = req_recycle_buf_S4_f;
        end
    end
end
always @ (posedge clk)
begin
    req_recycle_buf_S4_f <= req_recycle_buf_S4_next;
end
always @ *
begin
    req_recycle_S4 = req_recycle_cur_S4 | req_recycle_buf_S4_f;
end
reg smc_rd_diag_en_buf_S4_next;
reg smc_rd_en_buf_S4_next;
reg smc_rd_diag_en_buf_S4_f;
reg smc_rd_en_buf_S4_f;
always @ *
begin
    if (!rst_n)
    begin
        smc_rd_diag_en_buf_S4_next = 0;
        smc_rd_en_buf_S4_next = 0;
    end
    else if (!stall_smc_buf_S4)
    begin
        smc_rd_diag_en_buf_S4_next = smc_rd_diag_en_S4;
        smc_rd_en_buf_S4_next = smc_rd_en_S4;
    end
    else
    begin
        smc_rd_diag_en_buf_S4_next = smc_rd_diag_en_buf_S4_f;
        smc_rd_en_buf_S4_next = smc_rd_en_buf_S4_f;
    end
end
always @ (posedge clk)
begin
    smc_rd_diag_en_buf_S4_f <= smc_rd_diag_en_buf_S4_next;
    smc_rd_en_buf_S4_f <= smc_rd_en_buf_S4_next;
end
always @ *
begin
    smc_rd_diag_en_buf_S4 = smc_rd_diag_en_buf_S4_f;
    smc_rd_en_buf_S4 = smc_rd_en_buf_S4_f;
end
always @ *
begin
    if(valid_S4)
        begin
        if (~special_addr_type_S4_f && req_recycle_S4)
        begin
            mshr_wr_data_en_S4 = ~stall_S4;
            mshr_wr_state_en_S4 = ~stall_S4;
            mshr_inv_flag_S4 = 1'b0;
        end
        else if (load_store_mem_S4)
        begin
            mshr_wr_data_en_S4 = msg_send_valid_S4 && (msg_send_type_S4 == msg0_send_type_S4) && msg_send_ready_S4;
            mshr_wr_state_en_S4 = msg_send_valid_S4 && (msg_send_type_S4 == msg0_send_type_S4) && msg_send_ready_S4;
            mshr_inv_flag_S4 = 1'b0;
        end
        else if (msg_send_type_S4 == 8'd18)
        begin
            mshr_wr_data_en_S4 = ((msg_send_valid_S4 && msg_send_ready_S4 && (dir_sharer_counter_S4 == 1)) || (~stall_S4))
                              && mshr_wr_data_en_S4_f;
            mshr_wr_state_en_S4 = ((msg_send_valid_S4 && msg_send_ready_S4 && (dir_sharer_counter_S4 == 1)) || (~stall_S4))
                               && mshr_wr_state_en_S4_f;
            mshr_inv_flag_S4 = 1'b0;
        end
        else if ((msg_type_S4 == 8'd13) && l2_tag_hit_S4
              && (l2_way_state_mesi_S4 == 2'b10) && l2_way_state_subline_S4[addr_S4[5:4]]
              && req_from_owner_S4)
        begin
            mshr_wr_data_en_S4 = ~stall_S4;
            mshr_wr_state_en_S4 = ~stall_S4;
            mshr_inv_flag_S4 = 1'b0;
        end
        
        else if (csm_en && mshr_smc_miss_S4_f && (~mshr_wr_state_en_S4_f))
        begin
            mshr_wr_data_en_S4 = 1'b0;
            mshr_wr_state_en_S4 = ~stall_S4;
            mshr_inv_flag_S4 = 1'b1;
        end
        
        else
        begin
            mshr_wr_data_en_S4 = ~stall_S4 && mshr_wr_data_en_S4_f;
            mshr_wr_state_en_S4 = ~stall_S4 && mshr_wr_state_en_S4_f;
            mshr_inv_flag_S4 = 1'b0;
        end
    end
    else
    begin
        mshr_wr_data_en_S4 = 1'b0;
        mshr_wr_state_en_S4 = 1'b0;
        mshr_inv_flag_S4 = 1'b0;
    end
end
always @ *
begin
    if (valid_S4 && (!req_recycle_S4) && (msg_send_type_S4 == 8'd18)
     && (msg_send_valid_S4 && msg_send_ready_S4 && (dir_sharer_counter_S4 == 1) && stall_S4)
     && mshr_wr_data_en_S4_f)
    begin
        inv_fwd_pending_S4 = 1'b1;
    end
    else
    begin
        inv_fwd_pending_S4 = 1'b0;
    end
end
always @ *
begin
    addr_type_S4 = addr_S4[39:32];
    addr_op_S4 = addr_S4[31:30];
end
always @ *
begin
    if (!rst_n)
    begin
        stall_before_S4_next = 0;
    end
    else
    begin
        stall_before_S4_next = stall_S4;
    end
end
always @ (posedge clk)
begin
    stall_before_S4_f <= stall_before_S4_next;
end
reg [19-1:0] cs_S4;
always @ *
begin
    if (valid_S4)
    begin
        if (special_addr_type_S4_f)
        begin
            if (msg_type_S4_f == 8'd15)
            begin
                
                
                cs_S4 = {n,         y,          8'd28,  n,          8'd30};
            end
            else
            begin
                cs_S4 = {n,         y,          8'd29,  n,          8'd30};
            end
        end
        else if(req_recycle_S4)
        begin
            cs_S4 = {19{1'b0}};
        end
        else
        begin
            if (msg_type_S4_f == 8'd32)
            begin
                cs_S4 = {n,         y,          8'd33,    n,          8'd30};
            end
            else if (msg_type_S4_f == 8'd8)
            begin
                cs_S4 = {n,         n,          8'd30,    n,          8'd30};
            end
            else if (msg_type_S4_f == 8'd13)
            begin
                cs_S4 = {n,         n,          8'd30,    n,          8'd30};
            end
            else if (l2_evict_S4)
            begin
                begin
                    case (l2_way_state_mesi_S4)
                    2'b01, 2'b11:
                    begin
                        cs_S4 = {y,         y,          8'd18,    n,          8'd30};
                    end
                    2'b10:
                    begin
                        cs_S4 = {y,         y,          8'd17,    n,          8'd30};
                    end
                    2'b00:
                    begin
                        case (l2_way_state_vd_S4)
                        2'b10:
                        begin
                            if (msg_type_S4_f == 8'd34)
                            begin
                                cs_S4 = {n,         y,          8'd29,    n,          8'd30};
                            end
                            else if (msg_type_S4_f == 8'd14)
                            begin
                                
                                
                                
                                
                                    cs_S4 = {n,         y,          8'd19,    n,          8'd30};
                                
                            end
                            else
                            begin
                                cs_S4 = {n,         y,          8'd19,    n,          8'd30};
                            end
                        end
                        2'b11:
                        begin
                            if (msg_type_S4_f == 8'd34)
                            begin
                                cs_S4 = {n,         y,          8'd29,    y,          8'd20};
                            end
                            else if (msg_type_S4_f == 8'd14)
                            begin
                                
                                
                                
                                
                                    cs_S4 = {n,         y,          8'd19,    y,          8'd20};
                                
                            end
                            else
                            begin
                                cs_S4 = {n,         y,          8'd19,    y,          8'd20};
                            end
                        end
                        default:
                        begin
                            cs_S4 = {19{1'bx}};
                        end
                        endcase
                    end
                    default:
                    begin
                        cs_S4 = {19{1'bx}};
                    end
                    endcase
                end
            end
            else if (!l2_tag_hit_S4)
            begin
                begin
                    if (msg_type_S4_f == 8'd35 || msg_type_S4_f == 8'd34)
                    begin
                        cs_S4 = {n,         y,          8'd29,    n,          8'd30};
                    end
                    else if (msg_type_S4_f == 8'd15)
                    begin
                        if (msg_from_mshr_S4_f)
                        begin
                            
                            
                            cs_S4 = {n,          y,          8'd28,  n,          8'd30};
                        end
                        else
                        begin
                            cs_S4 = {n,          y,          8'd15,n,          8'd30};
                        end
                    end
                    else if (msg_type_S4_f == 8'd14)
                    begin
                        
                        
                        
                        
                            cs_S4 = {n,         y,          8'd19,    n,          8'd30};
                        
                    end
                    else
                    begin
                        cs_S4 = {n,         y,          8'd19,    n,          8'd30};
                    end
                end
            end
            else begin
            case (msg_type_S4_f)
                
                8'd35, 8'd34:
                begin
                   case (l2_way_state_mesi_S4)
                    2'b00:
                    begin
                        case (l2_way_state_vd_S4)
                        2'b10:
                        begin
                            cs_S4 = {n,         y,          8'd29,    n,          8'd30};
                        end
                        2'b11:
                        begin
                            cs_S4 = {n,         y,          8'd29,    y,          8'd20};
                        end
                        default:
                        begin
                            cs_S4 = {19{1'bx}};
                        end
                        endcase
                    end
                    2'b01, 2'b11:
                    begin
                        cs_S4 = {y,         y,          8'd18,    n,          8'd30};
                    end
                    2'b10:
                    begin
                        cs_S4 = {y,         y,          8'd17,   n,          8'd30};
                    end
                    default:
                    begin
                        cs_S4 = {19{1'bx}};
                    end
                    endcase
                end
                8'd15:
                begin
                   case (l2_way_state_mesi_S4)
                    2'b00:
                    begin
                        case (l2_way_state_vd_S4)
                        2'b10:
                        begin
                            cs_S4 = {n,         y,          8'd15,    n,          8'd30};
                        end
                        2'b11:
                        begin
                            cs_S4 = {n,         y,          8'd20,    n,          8'd30};
                        end
                        default:
                        begin
                            cs_S4 = {19{1'bx}};
                        end
                        endcase
                    end
                    2'b01, 2'b11:
                    begin
                        cs_S4 = {y,         y,          8'd18,    n,          8'd30};
                    end
                    2'b10:
                    begin
                        cs_S4 = {y,         y,          8'd17,   n,          8'd30};
                    end
                    default:
                    begin
                        cs_S4 = {19{1'bx}};
                    end
                    endcase
                end
                8'd14:
                begin
                   case (l2_way_state_mesi_S4)
                    2'b00:
                    begin
                        case (l2_way_state_vd_S4)
                        2'b10:
                        begin
                            cs_S4 = {n,         y,          8'd29,    n,          8'd30};
                        end
                        2'b11:
                        begin
                            cs_S4 = {n,         y,          8'd20,    n,          8'd30};
                        end
                        default:
                        begin
                            cs_S4 = {19{1'bx}};
                        end
                        endcase
                    end
                    2'b01, 2'b11:
                    begin
                        cs_S4 = {y,         y,          8'd18,    n,          8'd30};
                    end
                    2'b10:
                    begin
                        cs_S4 = {y,         y,          8'd17,   n,          8'd30};
                    end
                    default:
                    begin
                        cs_S4 = {19{1'bx}};
                    end
                    endcase
                end
                8'd31:
                begin
                    case (l2_way_state_mesi_S4)
                    2'b00:
                    begin
                        cs_S4 = {n,         y,          8'd29,    n,          8'd30};
                    end
                    2'b01, 2'b11:
                    begin
                        if (cache_type_S4_f == l2_way_state_cache_type_S4)
                        begin
                            cs_S4 = {n,         y,          8'd29,    n,          8'd30};
                        end
                        else
                        begin
                            cs_S4 = {y,         y,          8'd18,    n,          8'd30};
                        end
                    end
                    2'b10:
                    begin
                        if (req_from_owner_S4 && (cache_type_S4_f == l2_way_state_cache_type_S4))
                        begin
                            cs_S4 = {n,         y,          8'd29,    n,          8'd30};
                        end
                        else if (cache_type_S4_f != l2_way_state_cache_type_S4)
                        begin
                            cs_S4 = {y,         y,          8'd17,   n,          8'd30};
                        end
                        else
                        begin
                            cs_S4 = {y,         y,          8'd16,   n,          8'd30};
                        end
                    end
                    default:
                    begin
                        cs_S4 = {19{1'bx}};
                    end
                    endcase
                end
                8'd60:   
                begin
                    case (l2_way_state_mesi_S4)
                    2'b00:
                    begin
                        cs_S4 = {n,         y,          8'd29,    n,          8'd30};
                    end
                    2'b01:
                    begin
                        cs_S4 = {y,         y,          8'd18,    n,          8'd30};
                    end
                    2'b10:
                    begin
                        if (req_from_owner_S4 && (cache_type_S4_f == l2_way_state_cache_type_S4))
                        begin
                            cs_S4 = {n,         y,          8'd29,    n,          8'd30};
                        end
                        else
                        begin
                            cs_S4 = {y,         y,          8'd17,    n,          8'd30};
                        end
                    end
                    default:
                    begin
                        cs_S4 = {19{1'bx}};
                    end
                    endcase
                end
                8'd1:
                begin
                    cs_S4 = {n,         y,          8'd28,    n,          8'd30};
                end
                8'd2:
                begin
                    case (l2_way_state_mesi_S4)
                    2'b00:
                    begin
                        cs_S4 = {n,         y,          8'd29,    n,          8'd30};
                    end
                    2'b01, 2'b11:
                    begin
                        cs_S4 = {y,         y,          8'd18,    n,          8'd30};
                    end
                    2'b10:
                    begin
                        if (req_from_owner_S4 && (cache_type_S4_f == l2_way_state_cache_type_S4))
                        begin
                            cs_S4 = {n,         y,          8'd29,    n,          8'd30};
                        end
                        else
                        begin
                            cs_S4 = {y,         y,          8'd17,    n,          8'd30};
                        end
                    end
                    default:
                    begin
                        cs_S4 = {19{1'bx}};
                    end
                    endcase
                end
                8'd6, 8'd10,
                8'd44,
                8'd45,
                8'd46,
                8'd47,
                8'd48,
                8'd49,
                8'd50,
                8'd51:
                begin
                    case (l2_way_state_mesi_S4)
                    2'b00:
                    begin
                        cs_S4 = {n,         y,          8'd29,    n,          8'd30};
                    end
                    2'b01, 2'b11:
                    begin
                        cs_S4 = {y,         y,          8'd18,    n,          8'd30};
                    end
                    2'b10:
                    begin
                        cs_S4 = {y,         y,          8'd17,    n,          8'd30};
                    end
                    default:
                    begin
                        cs_S4 = {19{1'bx}};
                    end
                    endcase
                end
                8'd7, 8'd11,
                8'd52,
                8'd53,
                8'd54,
                8'd55,
                8'd56,
                8'd57,
                8'd58,
                8'd59:
                begin
                    case (l2_way_state_mesi_S4)
                    2'b00:
                    begin
                        cs_S4 = {n,         n,          8'd30,    n,          8'd30};
                    end
                    2'b01, 2'b11:
                    begin
                        cs_S4 = {y,         y,          8'd18,    n,          8'd30};
                    end
                    2'b10:
                    begin
                        cs_S4 = {y,         y,          8'd17,    n,          8'd30};
                    end
                    default:
                    begin
                        cs_S4 = {19{1'bx}};
                    end
                    endcase
                end
                default:
                begin
                    cs_S4 = {19{1'bx}};
                end
            endcase
            end
        end
    end
    else
    begin
        cs_S4 = {19{1'b0}};
    end
end
always @ *
begin
    msg0_send_valid_S4 = !(global_stall_S4 || stall_inv_counter_S4 || smc_stall_S4 || broadcast_stall_S4) && cs_S4[17];
    msg0_send_type_S4 = cs_S4[16:9];
    msg1_send_valid_S4 = !(global_stall_S4 || stall_inv_counter_S4|| smc_stall_S4 || broadcast_stall_S4) && cs_S4[8];
    msg1_send_type_S4 = cs_S4[7:0];
end
always @ *
begin
    load_store_mem_S4 = cs_S4[17] && cs_S4[8] &&
                       (msg0_send_type_S4 == 8'd19 || msg0_send_type_S4 == 8'd14)
                     &&(msg1_send_type_S4 == 8'd20);
end
localparam msg_state_0 = 1'b0;
localparam msg_state_1 = 1'b1;
reg msg_state_S4_f;
reg msg_state_S4_next;
always @ *
begin
    if (!rst_n)
    begin
        msg_state_S4_next = msg_state_0;
    end
    else if (msg0_send_valid_S4 && msg1_send_valid_S4 && valid_S4
    && !(dir_data_stall_S4 || smc_stall_S4 || (msg_send_valid_S4 && !msg_send_ready_S4) || global_stall_S4 || broadcast_stall_S4))
    begin
        if (msg_state_S4_f == msg_state_0)
        begin
            msg_state_S4_next = msg_state_1;
        end
        else
        begin
            if (l2_load_data_subline_S4_f == 2'd3)
            begin
                msg_state_S4_next = msg_state_0;
            end
            else
            begin
                msg_state_S4_next = msg_state_1;
            end
        end
    end
    else
    begin
        msg_state_S4_next = msg_state_S4_f;
    end
end
always @ (posedge clk)
begin
    msg_state_S4_f <= msg_state_S4_next;
end
always @ *
begin
    if (msg_state_S4_f == msg_state_0)
    begin
        msg_send_valid_S4 = msg0_send_valid_S4;
        msg_send_type_pre_S4 = msg0_send_type_S4;
    end
    else
    begin
        msg_send_valid_S4 = msg1_send_valid_S4;
        msg_send_type_pre_S4 = msg1_send_type_S4;
    end
end
always @ *
begin
    if (smc_miss_S4)
    begin
        msg_send_type_S4 = 8'd14;
    end
    else
    begin
        msg_send_type_S4 = msg_send_type_pre_S4;
    end
end
localparam smc_state_0 = 1'b0;
localparam smc_state_1 = 1'b1;
reg smc_state_S4_f;
reg smc_state_S4_next;
always @ *
begin
    if (!rst_n)
    begin
        smc_state_S4_next = smc_state_0;
    end
    else if (smc_rd_en_S4 && (~stall_smc_buf_S4))
    begin
        if (smc_state_S4_f == smc_state_0)
        begin
            smc_state_S4_next = smc_state_1;
        end
        else
        begin
            smc_state_S4_next = smc_state_0;
        end
    end
    else
    begin
        smc_state_S4_next = smc_state_S4_f;
    end
end
always @ (posedge clk)
begin
    smc_state_S4_f <= smc_state_S4_next;
end
always @ *
begin
    smc_stall_S4 = smc_rd_en_S4 && (smc_state_S4_f == smc_state_0);
end
reg [3-1:0] mshr_empty_index_buf_S4_f;
reg [3-1:0] mshr_empty_index_buf_S4_next;
reg [3-1:0] mshr_empty_index_sel_S4;
always @ *
begin
    if (stall_before_S4_f)
    begin
        mshr_empty_index_sel_S4 = mshr_empty_index_buf_S4_f;
    end
    else
    begin
        mshr_empty_index_sel_S4 = mshr_empty_index_S4;
    end
end
always @ *
begin
    if (!rst_n)
    begin
        mshr_empty_index_buf_S4_next = {3{1'b0}};
    end
    else if (stall_S4 && !stall_before_S4_f)
    begin
        mshr_empty_index_buf_S4_next = mshr_empty_index_S4;
    end
    else
    begin
        mshr_empty_index_buf_S4_next = mshr_empty_index_buf_S4_f;
    end
end
always @ (posedge clk)
begin
    mshr_empty_index_buf_S4_f <= mshr_empty_index_buf_S4_next;
end
always @ *
begin
    if (msg_send_valid_S4)
    begin
        case (msg_send_type_S4)
        8'd16, 8'd17, 8'd18:
        begin
            msg_send_mode_S4 = 3'd4;
            msg_send_length_S4 = 8'd2;
            msg_send_data_size_S4 = 3'b101;
            msg_send_cache_type_S4 = l2_way_state_cache_type_S4;
            msg_send_mshrid_S4 = mshr_wr_index_in_S4;
        end
        8'd28:
        begin
            msg_send_mode_S4 = 3'd1;
            msg_send_length_S4 = 8'd0;
            msg_send_data_size_S4 = 3'b000;
            msg_send_cache_type_S4 = cache_type_S4_f;
            msg_send_mshrid_S4 = mshrid_S4;
        end
        8'd29:
        begin
            
            if (special_addr_type_S4_f)
            begin
                msg_send_mode_S4 = 3'd3;
                msg_send_length_S4 = 8'd2;
                
                msg_send_cache_type_S4 = cache_type_S4_f;
                msg_send_mshrid_S4 = mshrid_S4;
            end
            else if (cache_type_S4_f == 1'b0)
            begin
                msg_send_mode_S4 = 3'd3;
                msg_send_length_S4 = 8'd2;
                
                msg_send_cache_type_S4 = cache_type_S4_f;
                msg_send_mshrid_S4 = mshrid_S4;
            end
            else
            begin
                
                msg_send_length_S4 = 8'd4;
                
                msg_send_cache_type_S4 = cache_type_S4_f;
                msg_send_mshrid_S4 = mshrid_S4;
                if (l2_load_data_subline_S4_f == 2'd0)
                begin
                    msg_send_mode_S4 = 3'd3;
                end
                else
                begin
                    msg_send_mode_S4 = 3'd7;
                end
            end
        end
        8'd19:
        begin
            msg_send_mode_S4 = 3'd4;
            msg_send_length_S4 = 8'd2;
            msg_send_data_size_S4 = data_size_S4_f;
            msg_send_cache_type_S4 = 1'b0;
            msg_send_mshrid_S4 = mshr_wr_index_in_S4;
        end
        8'd14:
        begin
            msg_send_mode_S4 = 3'd4;
            msg_send_length_S4 = 8'd2;
            msg_send_data_size_S4 = data_size_S4_f;
            if (smc_miss_S4)
            begin
                msg_send_data_size_S4 = 3'b101;
            end
            msg_send_cache_type_S4 = cache_type_S4_f;
            msg_send_mshrid_S4 = mshr_wr_index_in_S4;
        end
        8'd15:
        begin
            msg_send_mode_S4 = 3'd5;
            msg_send_length_S4 = 8'd3;
            msg_send_data_size_S4 = data_size_S4_f;
            msg_send_cache_type_S4 = cache_type_S4_f;
            msg_send_mshrid_S4 = mshr_wr_index_in_S4;
        end
        8'd33:
        begin
            msg_send_mode_S4 = 3'd2;
            msg_send_length_S4 = 8'd1;
            msg_send_data_size_S4 = data_size_S4_f;
            msg_send_cache_type_S4 = cache_type_S4_f;
            msg_send_mshrid_S4 = mshrid_S4;
        end
        8'd20:
        begin
            msg_send_length_S4 = 8'd10;
            msg_send_data_size_S4 = data_size_S4_f;
            msg_send_cache_type_S4 = 1'b0;
            msg_send_mshrid_S4 = mshr_wr_index_in_S4;
            if (l2_load_data_subline_S4_f == 2'd0)
            begin
                msg_send_mode_S4 = 3'd6;
            end
            else
            begin
                msg_send_mode_S4 = 3'd7;
            end
        end
        default:
        begin
            msg_send_mode_S4 = 3'd0;
            msg_send_length_S4 = 8'd0;
            msg_send_data_size_S4 = 3'b000;
            msg_send_cache_type_S4 = 1'b0;
            msg_send_mshrid_S4 = mshrid_S4;
        end
        endcase
    end
    else
    begin
        msg_send_mode_S4 = 3'd0;
        msg_send_length_S4 = 8'd0;
        msg_send_data_size_S4 = 3'b000;
        msg_send_cache_type_S4 = 1'b0;
        msg_send_mshrid_S4 = mshrid_S4;
    end
end
always @ *
begin
    msg_send_l2_miss_S4 = l2_miss_S4_f;
end
always @ *
begin
    if ((msg_send_type_S4 == 8'd33)
    || special_addr_type_S4_f
    || ((msg_type_S4_f == 8'd15) && !l2_tag_hit_S4))
    begin
        msg_send_subline_vector_S4 = {4{1'b0}};
    end
    else if (msg_send_type_S4 == 8'd18)
    begin
        msg_send_subline_vector_S4 = {4{1'b1}};
    end
    else
    begin
        msg_send_subline_vector_S4 = l2_way_state_subline_S4;
    end
end
always @ *
begin
    if ((msg_type_S4_f == 8'd2 || msg_type_S4_f == 8'd60) && msg_send_type_S4 == 8'd29)
    begin
        msg_send_mesi_S4 = 2'b11;
    end
    else if ((msg_send_type_S4 == 8'd33)
    || special_addr_type_S4_f
    || ((msg_type_S4_f == 8'd15) && !l2_tag_hit_S4))
    begin
        msg_send_mesi_S4 = 2'b00;
    end
    else
    begin
        if (state_mesi_S4_f == 2'b11)
        begin
            msg_send_mesi_S4 = 2'b01;
        end
        else
        begin
            msg_send_mesi_S4 = state_mesi_S4_f;
        end
    end
end
always @ *
begin
    l2_access_valid_S4 = valid_S4 && !stall_S4 && msg_send_valid_S4
                     && (msg_send_type_S4 == 8'd29 || msg_send_type_S4 == 8'd28);
end
always @ *
begin
    l2_miss_valid_S4 = l2_access_valid_S4 && msg_send_l2_miss_S4;
end
always @ *
begin
    msg_stall_S4 = msg0_send_valid_S4 && msg1_send_valid_S4
               && (msg_state_S4_f == msg_state_0);
end
reg [64-1:0] dir_data_buf_S4_f;
reg [64-1:0] dir_data_buf_S4_next;
reg [64-1:0] dir_data_trans_S4;
always @ *
begin
    if (stall_before_S4_f)
    begin
        dir_data_sel_S4 = dir_data_buf_S4_f;
    end
    else
    begin
        
        if(mshr_smc_miss_S4_f)
        begin
            
            dir_data_sel_S4 = (dir_data_S4 >> mshr_miss_lsid_S4) << mshr_miss_lsid_S4;
        end
        else
        
        begin
            dir_data_sel_S4 = dir_data_S4;
        end
    end
end
always @ *
begin
    if (!rst_n)
    begin
        dir_data_buf_S4_next = {64{1'b0}};
    end
    else if ((stall_S4 && !stall_before_S4_f) && (msg_send_type_pre_S4 == 8'd18) && (l2_way_state_mesi_S4 != 2'b11))
    begin
        if (msg_stall_S4 || smc_stall_S4 || (msg_send_valid_S4 && !msg_send_ready_S4)
         || global_stall_S4 || stall_inv_counter_S4 )
        begin
            if(mshr_smc_miss_S4_f)
            begin
                dir_data_buf_S4_next = (dir_data_S4 >> mshr_miss_lsid_S4) << mshr_miss_lsid_S4;
            end
            else
            begin
                dir_data_buf_S4_next = dir_data_S4;
            end
        end
        else
        begin
            dir_data_buf_S4_next = dir_data_trans_S4;
        end
    end
    else if (!((msg_send_valid_S4 && !msg_send_ready_S4) || global_stall_S4 || smc_stall_S4 || broadcast_stall_S4
             || stall_inv_counter_S4) && dir_data_stall_S4)
    begin
        dir_data_buf_S4_next = dir_data_trans_S4;
    end
    else
    begin
        dir_data_buf_S4_next = dir_data_buf_S4_f;
    end
end
always @ (posedge clk)
begin
    dir_data_buf_S4_f <= dir_data_buf_S4_next;
end
wire [64-1:0] dir_sharer_mask_S4;
wire nonzero_sharer_S4;
l2_priority_encoder_6 priority_encoder_6bits( 
    .data_in        (dir_data_sel_S4),
    .data_out       (dir_sharer_S4),
    .data_out_mask  (dir_sharer_mask_S4),
    .nonzero_out    (nonzero_sharer_S4)
);
reg [6-1:0] dir_sharer_counter_S4_f;
reg [6-1:0] dir_sharer_counter_S4_next;
always @ *
begin
    if (!rst_n)
    begin
        dir_sharer_counter_S4_next = 1;
    end
    else if (msg_send_valid_S4 && msg_send_ready_S4 && (msg_send_type_pre_S4 == 8'd18))
    begin
        if (dir_data_stall_S4)
        begin
            dir_sharer_counter_S4_next = dir_sharer_counter_S4_f + 1;
        end
        else
        begin
            dir_sharer_counter_S4_next = 1;
        end
    end
    else
    begin
        dir_sharer_counter_S4_next = dir_sharer_counter_S4_f;
    end
end
always @ (posedge clk)
begin
    dir_sharer_counter_S4_f <= dir_sharer_counter_S4_next;
end
always @ *
begin
    dir_sharer_counter_S4 = dir_sharer_counter_S4_f;
end
always @ *
begin
    dir_data_trans_S4 = dir_data_sel_S4 & (dir_sharer_mask_S4);
end
localparam broadcast_state_0 = 1'b0;
localparam broadcast_state_1 = 1'b1;
reg broadcast_state_S4_f;
reg broadcast_state_S4_next;
always @ *
begin
    if (!rst_n)
    begin
        broadcast_state_S4_next = broadcast_state_0;
    end
    else if (valid_S4 && (~stall_S4))
    begin
        broadcast_state_S4_next = broadcast_state_0;
    end
    else if (valid_S4 && (l2_way_state_mesi_S4 == 2'b11) && (msg_send_type_S4 == 8'd18)
         && (~(msg_stall_S4 || smc_stall_S4 || (msg_send_valid_S4 && !msg_send_ready_S4)
         || global_stall_S4 || stall_inv_counter_S4 || broadcast_stall_S4)))
    begin
        if (broadcast_state_S4_f == broadcast_state_0)
        begin
            broadcast_state_S4_next = broadcast_state_1;
        end
        else
        begin
            broadcast_state_S4_next = broadcast_state_S4_f;
        end
    end
    else
    begin
        broadcast_state_S4_next = broadcast_state_S4_f;
    end
end
always @ (posedge clk)
begin
    broadcast_state_S4_f <= broadcast_state_S4_next;
end
always @ *
begin
    broadcast_stall_S4 = (l2_way_state_mesi_S4 == 2'b11) && (msg_send_type_S4 == 8'd18)
                      && (broadcast_state_S4_f == broadcast_state_0) && (~broadcast_counter_avail_S4)
                      && (~(msg_from_mshr_S4_f && mshr_smc_miss_S4_f));
end
always @ *
begin
    broadcast_counter_op_val_S4 = valid_S4 && (~stall_smc_buf_S4) && (~smc_stall_S4) && (l2_way_state_mesi_S4 == 2'b11)
    && (msg_send_type_S4 == 8'd18) && (~((broadcast_state_S4_f == broadcast_state_1) && broadcast_counter_zero_S4));
end
always @ *
begin
    if (broadcast_counter_op_val_S4)
    begin
        broadcast_counter_op_S4 = 2'd2;
    end
    else
    begin
        broadcast_counter_op_S4 = 2'd0;
    end
end
always @ *
begin
    if (l2_way_state_mesi_S4 == 2'b11)
    begin
        dir_data_stall_S4 = (msg_send_type_S4 == 8'd18) && (~broadcast_counter_max_S4);
    end
    else
    begin
        dir_data_stall_S4 = (msg_send_type_S4 == 8'd18) && (| dir_data_trans_S4[64-1:0]);
    end
end
always @ *
begin
    state_wr_en_real_S4 = valid_S4 && !dir_data_stall_S4 &&  msg_send_valid_S4 && (msg_send_type_pre_S4 == 8'd18);
end
always @ *
begin
    if (load_store_mem_S4)
    begin
        state_wr_en_S4 = msg_send_valid_S4 && (msg_send_type_S4 == msg0_send_type_S4) && msg_send_ready_S4 && ~(req_recycle_S4 && ~special_addr_type_S4_f);
    end
    else
    begin
        state_wr_en_S4 = !stall_S4 && (state_wr_en_real_S4 || state_wr_en_S4_f) && ~(req_recycle_S4 && ~special_addr_type_S4_f);
    end
end
always @ *
begin
    smc_rd_en_S4 = valid_S4 &&
                ((special_addr_type_S4_f
                && (addr_S4[39:32] == 8'ha2)
                && (msg_type_S4 == 8'd14))
                || (csm_en
                && (((msg_send_type_pre_S4 == 8'd18) && (l2_way_state_mesi_S4 != 2'b11)))));
           
           
end
always @ *
begin
    smc_rd_diag_en_S4 =
                (special_addr_type_S4_f
                && (addr_S4[39:32] == 8'ha2)
                && (msg_type_S4 == 8'd14));
end
always @ *
begin
    smc_miss_S4 = smc_rd_en_S4  && ~smc_rd_diag_en_S4 && (~smc_hit_S4);
end
always @ *
begin
    if (msg_type_S4_f == 8'd6 && (msg_send_valid_S4 && msg_send_type_S4 == 8'd29)
    && valid_S4 && !stall_S4)
    begin
        cas_cmp_en_S4 = y;
    end
    else
    begin
        cas_cmp_en_S4 = n;
    end
end
always @ *
begin
    if ((msg_type_S4_f == 8'd6
        || msg_type_S4_f == 8'd10
        || msg_type_S4_f == 8'd44
        || msg_type_S4_f == 8'd45
        || msg_type_S4_f == 8'd46
        || msg_type_S4_f == 8'd47
        || msg_type_S4_f == 8'd48
        || msg_type_S4_f == 8'd49
        || msg_type_S4_f == 8'd50
        || msg_type_S4_f == 8'd51)
    && (msg_send_valid_S4 && msg_send_type_S4 == 8'd29)
    && valid_S4 && !stall_S4)
    begin
        atomic_read_data_en_S4 = y;
    end
    else
    begin
        atomic_read_data_en_S4 = n;
    end
end
always @ *
begin
    cas_cmp_data_size_S4 = data_size_S4_f;
end
always @ *
begin
    reg_rd_en_S4 = valid_S4  && (msg_type_S4 == 8'd14)
               && ((addr_type_S4 == 8'ha9)
                || (addr_type_S4 == 8'ha7)
                || (addr_type_S4 == 8'ha8)
                || (addr_type_S4 == 8'haa)
                || (addr_type_S4 == 8'hab));
end
always @ *
begin
    reg_rd_addr_type_S4 = addr_type_S4;
end
always @ *
begin
    if (state_wr_en_real_S4)
    begin
        state_wr_sel_S4 = 1'b1;
    end
    else
    begin
        state_wr_sel_S4 = 1'b0;
    end
end
always @ *
begin
    
    if (mshr_smc_miss_S4_f)
    begin
        mshr_wr_index_in_S4 = mshr_pending_index_S4_f;
    end
    else
    
    begin
        mshr_wr_index_in_S4 = mshr_empty_index_sel_S4;
    end
end
always @ *
begin
    mshr_inv_counter_rd_index_in_S4 = mshr_wr_index_in_S4;
end
always @ *
begin
    stall_inv_counter_S4 = valid_S4 && ((global_stall_S1 && (pipe2_msg_type_S1 == 8'd23))
                                     || (global_stall_S2 && (pipe2_msg_type_S2 == 8'd23)))
                       && (msg_send_type_pre_S4 == 8'd18);
                   
end
always @ *
begin
    stall_smc_buf_S4 = valid_S4 && (global_stall_S4
           || (msg_send_valid_S4 && !msg_send_ready_S4)
           || broadcast_stall_S4
           || stall_inv_counter_S4);
end
always @ *
begin
    stall_S4 = valid_S4 && (global_stall_S4 || msg_stall_S4 || dir_data_stall_S4
           || (msg_send_valid_S4 && !msg_send_ready_S4)
           || stall_inv_counter_S4
           || broadcast_stall_S4
           || smc_stall_S4);
end
endmodule
      
 
module l2_pipe1_dpath(
    input wire clk,
    input wire rst_n,
    
    input wire csm_en,
    
    input wire [22-1:0] smt_base_addr,
    
    
    input wire [40-1:0] cam_mshr_addr_S1,
    input wire [8-1:0] cam_mshr_mshrid_S1,
    input wire [2-1:0] cam_mshr_way_S1,
    input wire [14-1:0] cam_mshr_src_chipid_S1,
    input wire [8-1:0] cam_mshr_src_x_S1,
    input wire [8-1:0] cam_mshr_src_y_S1,
    input wire [4-1:0] cam_mshr_src_fbits_S1,
    input wire [10-1:0] cam_mshr_sdid_S1,
    input wire [6-1:0] cam_mshr_lsid_S1,
    input wire [6-1:0] cam_mshr_miss_lsid_S1,
    input wire cam_mshr_recycled_S1,
    
    input wire mshr_pending_S1,
    input wire [40-1:0] pending_mshr_addr_S1,
    input wire [8-1:0] pending_mshr_mshrid_S1,
    input wire [2-1:0] pending_mshr_way_S1,
    input wire [14-1:0] pending_mshr_src_chipid_S1,
    input wire [8-1:0] pending_mshr_src_x_S1,
    input wire [8-1:0] pending_mshr_src_y_S1,
    input wire [4-1:0] pending_mshr_src_fbits_S1,
    input wire [10-1:0] pending_mshr_sdid_S1,
    input wire [6-1:0] pending_mshr_lsid_S1,
    input wire [6-1:0] pending_mshr_miss_lsid_S1,
    input wire pending_mshr_recycled_S1,
 
    input wire dis_flush_S1,
    
    input wire [40-1:0] msg_addr_S1,
    input wire [8-1:0] msg_mshrid_S1,
    input wire [14-1:0] msg_src_chipid_S1,
    input wire [8-1:0] msg_src_x_S1,
    input wire [8-1:0] msg_src_y_S1,
    input wire [4-1:0] msg_src_fbits_S1,
    input wire [10-1:0] msg_sdid_S1,
    input wire [6-1:0] msg_lsid_S1,
    
    input wire [64-1:0] msg_data_S1,
    
    input wire valid_S1,
    input wire stall_S1,
    input wire msg_from_mshr_S1, 
    
 
    
    
    input wire [64-1:0] msg_data_S2,
   
    input wire [15*4+2+4-1:0] state_data_S2,
    
    
    input wire [104-1:0] tag_data_S2,
    
    input wire msg_from_mshr_S2,
    input wire special_addr_type_S2,
    input wire [8-1:0] msg_type_S2,
    input wire [3-1:0] data_size_S2,
    input wire [1-1:0] cache_type_S2,
    input wire [2-1:0] dir_op_S2,
    input wire state_owner_en_S2,
    input wire [2-1:0] state_owner_op_S2,
    input wire state_subline_en_S2,
    input wire [2-1:0] state_subline_op_S2,
    input wire state_di_en_S2,
    input wire state_vd_en_S2,
    input wire [2-1:0] state_vd_S2,
    input wire state_mesi_en_S2,
    input wire [2-1:0] state_mesi_S2,
    input wire state_lru_en_S2,
    input wire [1-1:0] state_lru_op_S2,
    input wire state_rb_en_S2,
    input wire l2_ifill_32B_S2,
    input wire [2-1:0] l2_load_data_subline_S2,
    input wire valid_S2,
    input wire stall_S2,
    input wire stall_before_S2,
    input wire state_load_sdid_S2, 
    input wire data_clk_en_S2,
    input wire stall_real_S2,
    input wire [4-1:0] amo_alu_op_S2,
    
    
    input wire [144-1:0] data_data_S3,
    input wire valid_S3,
    input wire stall_S3,
    input wire stall_before_S3, 
    
    
    input wire valid_S4,
    input wire stall_S4,
    input wire stall_before_S4, 
    input wire cas_cmp_en_S4,
    input wire atomic_read_data_en_S4,
    input wire [3-1:0] cas_cmp_data_size_S4,
    input wire [6-1:0] dir_sharer_S4,
    input wire [6-1:0] dir_sharer_counter_S4,
    input wire [6-1:0] mshr_inv_counter_out_S4,
    input wire [8-1:0] msg_send_type_S4,
    input wire [8-1:0] msg_send_length_S4,
    input wire [8-1:0] msg_send_type_pre_S4,
    input wire state_wr_sel_S4,
    input wire [8-1:0] msg_type_S4,
    input wire [3-1:0] data_size_S4,
    input wire [1-1:0] cache_type_S4,
    input wire [1-1:0] l2_miss_S4,
    
    input wire smc_miss_S4,
    
    input wire special_addr_type_S4,
    input wire [64-1:0] dir_data_sel_S4,
    input wire [64-1:0] dir_data_S4,
    
    input wire stall_smc_buf_S4,
    
    input wire msg_from_mshr_S4,
    input wire req_recycle_S4,
    input wire inv_fwd_pending_S4,
    
    
    input wire [14-1:0] broadcast_chipid_out_S4,
    input wire [8-1:0] broadcast_x_out_S4,
    input wire [8-1:0] broadcast_y_out_S4,
    
    
    
    input wire [30-1:0] smc_data_out_S4,
    input wire [4-1:0] smc_valid_out_S4,
    input wire [14-1:0] smc_tag_out_S4,
    
    
    input wire [14-1:0] my_nodeid_chipid_S4,
    input wire [8-1:0] my_nodeid_x_S4,
    input wire [8-1:0] my_nodeid_y_S4,
    input wire [64-1:0] reg_data_out_S4,
    
    
    
    output reg [40-1:0] addr_S1,
    output reg [8-1:0] mshr_addr_in_S1,
    output reg [8-1:0] tag_addr_S1,
    output reg [8-1:0] state_rd_addr_S1,
    output reg [64-1:0] reg_data_in_S1,
    output reg [104-1:0] tag_data_in_S1,
    output reg [104-1:0] tag_data_mask_in_S1,
    
   
 
    output reg [40-1:0] addr_S2,
    output reg l2_tag_hit_S2,
    output reg l2_evict_S2,
    output reg l2_wb_S2,
    output reg [2-1:0] l2_way_state_mesi_S2,
    output reg [2-1:0] l2_way_state_vd_S2,
    output reg [1-1:0] l2_way_state_cache_type_S2,
    output reg [4-1:0] l2_way_state_subline_S2,
    output reg req_from_owner_S2,
    output reg addr_l2_aligned_S2,
    output reg [6-1:0] lsid_S2,
    output reg [8+2-1:0] dir_addr_S2,
    output reg [64-1:0] dir_data_in_S2,
    output reg [64-1:0] dir_data_mask_in_S2,
    output reg [8+2+2-1:0] data_addr_S2,
    output reg [144-1:0] data_data_in_S2,
    output reg [144-1:0] data_data_mask_in_S2,
    
    output reg [16-1:0] smc_wr_addr_in_S2,
    output reg [128-1:0] smc_data_in_S2,
    
    
    output reg [40-1:0] addr_S3,
    
    output reg [40-1:0] addr_S4,
    output reg [8+2+2-1:0] data_addr_S4,
    output reg l2_tag_hit_S4,
    output reg l2_evict_S4,
    output reg [2-1:0] l2_way_state_mesi_S4,
    output reg [6-1:0] l2_way_state_owner_S4,
    output reg [2-1:0] l2_way_state_vd_S4,
    output reg [4-1:0] l2_way_state_subline_S4,
    output reg [1-1:0] l2_way_state_cache_type_S4,
    output reg [8-1:0] mshrid_S4,
    output reg req_from_owner_S4,
    output reg cas_cmp_S4,
    output reg [6-1:0] mshr_miss_lsid_S4,
    output reg [6-1:0] lsid_S4,
    output reg corr_error_S4,
    output reg uncorr_error_S4,
    output reg [40-1:0] msg_send_addr_S4,
    output reg [14-1:0] msg_send_dst_chipid_S4,
    output reg [8-1:0] msg_send_dst_x_S4,
    output reg [8-1:0] msg_send_dst_y_S4,
    output reg [4-1:0] msg_send_dst_fbits_S4,
    output reg [128-1:0] msg_send_data_S4,
    output reg [120+2-1:0] mshr_data_in_S4,
    output wire [120+2-1:0] mshr_data_mask_in_S4,
    
    output reg [16-1:0] smc_rd_addr_in_buf_S4,
    
    output reg [8-1:0] state_wr_addr_S4,
    output reg [15*4+2+4-1:0] state_data_in_S4,
    output reg [15*4+2+4-1:0] state_data_mask_in_S4
);
localparam y = 1'b1;
localparam n = 1'b0;
wire [128-1:0] data_data_ecc_S4;
reg [8-1:0] mshrid_S1;
reg [14-1:0] src_chipid_S1;
reg [8-1:0] src_x_S1;
reg [8-1:0] src_y_S1;
reg [4-1:0] src_fbits_S1;
reg [10-1:0] sdid_S1;
reg [6-1:0] lsid_S1;
reg [40-1:0] addr_trans_S1;
reg recycled_S1;
always @ *
begin
    if (msg_from_mshr_S1)
    begin
        addr_S1 = pending_mshr_addr_S1;
        mshrid_S1 = pending_mshr_mshrid_S1;
        src_chipid_S1 = pending_mshr_src_chipid_S1;
        src_x_S1 = pending_mshr_src_x_S1;
        src_y_S1 = pending_mshr_src_y_S1;
        src_fbits_S1 = pending_mshr_src_fbits_S1;
        sdid_S1 = pending_mshr_sdid_S1;
        lsid_S1 = pending_mshr_lsid_S1;
        recycled_S1 = pending_mshr_recycled_S1;
 
    end
    else
    begin
        addr_S1 = msg_addr_S1;
        mshrid_S1 = msg_mshrid_S1;
        src_chipid_S1 = msg_src_chipid_S1;
        src_x_S1 = msg_src_x_S1;   
        src_y_S1 = msg_src_y_S1;   
        src_fbits_S1 = msg_src_fbits_S1;
        sdid_S1 = msg_sdid_S1;
        lsid_S1 = msg_lsid_S1;
        recycled_S1 = 1'b0;
    end
end
always @ *
begin
    if (dis_flush_S1)
    begin
        
        addr_trans_S1 = {addr_S1[5:0],addr_S1[33:6],6'd0};
    end
    else
    begin
        addr_trans_S1 = addr_S1;
    end
end
always @ *
begin
    if (~msg_from_mshr_S1)
    begin
        mshr_addr_in_S1 = addr_trans_S1[6+8-1:6];
    end
    else 
    begin
        mshr_addr_in_S1 = {8{1'b0}};
    end
end
always @ *
begin
    tag_addr_S1 = addr_trans_S1[6+8-1:6];
end
always @ *
begin
    state_rd_addr_S1 = addr_trans_S1[6+8-1:6];
end
reg [128-1:0] atomic_read_data_S1_f;
reg [128-1:0] atomic_read_data_S1_next;
always @ *
begin
    if (!rst_n)
    begin
        atomic_read_data_S1_next = 0;
    end
    else if (atomic_read_data_en_S4)
    begin
        atomic_read_data_S1_next = data_data_ecc_S4;
    end
    else
    begin
        atomic_read_data_S1_next = atomic_read_data_S1_f;
    end
end
always @ (posedge clk)
begin
    atomic_read_data_S1_f <= atomic_read_data_S1_next;
end
always @ *
begin
    reg_data_in_S1 = msg_data_S1;
end
always @ *
begin
    tag_data_in_S1 = {4{msg_data_S1[26-1:0]}};
end
always @ *
begin
    tag_data_mask_in_S1 = {{(4-1)*26{1'b0}},{26{1'b1}}} 
                       << (addr_trans_S1[6+8+2-1:6+8] * 26);
end
reg [40-1:0] addr_S2_f;
reg [8-1:0] mshrid_S2_f;
reg [14-1:0] src_chipid_S2_f;
reg [8-1:0] src_x_S2_f;
reg [8-1:0] src_y_S2_f;
reg [4-1:0] src_fbits_S2_f;
reg [10-1:0] sdid_S2_f;
reg [6-1:0] lsid_S2_f;
reg [2-1:0] mshr_way_S2_f;
reg [6-1:0] mshr_miss_lsid_S2_f;
reg [128-1:0] atomic_read_data_S2_f;
reg recycled_S2_f;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        addr_S2_f <= 0; 
        mshrid_S2_f <= 0;
        src_chipid_S2_f <= 0;
        src_x_S2_f <= 0;
        src_y_S2_f <= 0;
        src_fbits_S2_f <= 0;
        sdid_S2_f <= 0;
        lsid_S2_f <= 0;
        mshr_way_S2_f <= 0;
        mshr_miss_lsid_S2_f <= 0;
        atomic_read_data_S2_f <= 0;
        recycled_S2_f <= 0;
    end
    else if (!stall_S2)
    begin
        addr_S2_f <= addr_trans_S1;
        mshrid_S2_f <= mshrid_S1;
        src_chipid_S2_f <= src_chipid_S1;
        src_x_S2_f <= src_x_S1;
        src_y_S2_f <= src_y_S1;
        src_fbits_S2_f <= src_fbits_S1;
        sdid_S2_f <= sdid_S1;
        lsid_S2_f <= lsid_S1;
        
        mshr_way_S2_f <= (mshr_pending_S1 == 1'b1) ? pending_mshr_way_S1 : cam_mshr_way_S1;
        mshr_miss_lsid_S2_f <= (mshr_pending_S1 == 1'b1) ? pending_mshr_miss_lsid_S1 : cam_mshr_miss_lsid_S1;
 
        atomic_read_data_S2_f <= atomic_read_data_S1_f;
        recycled_S2_f <= recycled_S1;
    end
end
reg [64-1:0] return_data_S2;
reg [2-1:0] l2_way_sel_S2;
reg [15*4+2+4-1:0] state_data_in_S2;
reg [15*4+2+4-1:0] state_data_mask_in_S2;
always @ *
begin
    addr_S2 = addr_S2_f;
    lsid_S2 = lsid_S2_f;
end
reg [104-1:0] tag_data_buf_S2_f;
reg [104-1:0] tag_data_buf_S2_next;
reg [104-1:0] tag_data_trans_S2;
always @ *
begin
    if (!rst_n)
    begin
        tag_data_buf_S2_next = 0;
    end
    else if (stall_S2 && !stall_before_S2)
    begin
        tag_data_buf_S2_next = tag_data_S2;
    end
    else
    begin
        tag_data_buf_S2_next = tag_data_buf_S2_f;
    end
end
always @ (posedge clk)
begin
    tag_data_buf_S2_f <= tag_data_buf_S2_next;
end
always @ *
begin
    if (stall_before_S2)
    begin
        tag_data_trans_S2 = tag_data_buf_S2_f;
    end
    else
    begin
        tag_data_trans_S2 = tag_data_S2;
    end
end
wire [6-1:0] flat_id_S2;
xy_to_flat_id flat_id_gen(
    .flat_id    (flat_id_S2),
    .x_coord    (src_x_S2_f),
    .y_coord    (src_y_S2_f)
);
reg [15*4+2+4-1:0] state_data_buf_S2_f;
reg [15*4+2+4-1:0] state_data_buf_S2_next;
reg [15*4+2+4-1:0] state_data_trans_S2;
always @ *
begin
    if (!rst_n)
    begin
        state_data_buf_S2_next = 0;
    end
    else if (stall_S2 && !stall_before_S2)
    begin
        state_data_buf_S2_next = state_data_S2;
    end
    else
    begin
        state_data_buf_S2_next = state_data_buf_S2_f;
    end
end
always @ (posedge clk)
begin
    state_data_buf_S2_f <= state_data_buf_S2_next;
end
always @ *
begin
    if (stall_before_S2)
    begin
        state_data_trans_S2 = state_data_buf_S2_f;
    end
    else
    begin
        state_data_trans_S2 = state_data_S2;
    end
end
wire [2-1:0] l2_hit_way_sel_S2;
reg [2-1:0] l2_evict_way_sel_S2;
reg [2-1:0] l2_rb_bits_S2;
reg [4-1:0] l2_lru_bits_S2;
always @ *
begin
    l2_rb_bits_S2 = state_data_trans_S2[15*4+2+4-1:15*4+4];
    l2_lru_bits_S2 = state_data_trans_S2[15*4+4-1:15*4];
end
reg [26 - 1:0] tag_data_way_S2 [3:0];
reg [3:0] tag_hit_way_S2;
reg [15 - 1:0] state_way_S2 [3:0];
always @ *
begin
    tag_data_way_S2[0] = tag_data_trans_S2[26 * 1 - 1: 26 * 0];
    tag_data_way_S2[1] = tag_data_trans_S2[26 * 2 - 1: 26 * 1];
    tag_data_way_S2[2] = tag_data_trans_S2[26 * 3 - 1: 26 * 2];
    tag_data_way_S2[3] = tag_data_trans_S2[26 * 4 - 1: 26 * 3];
end
always @ *
begin
    state_way_S2[0] = state_data_trans_S2[15 * 1 - 1: 
15 * 0];
    state_way_S2[1] = state_data_trans_S2[15 * 2 - 1: 
15 * 1];
    state_way_S2[2] = state_data_trans_S2[15 * 3 - 1: 
15 * 2];
    state_way_S2[3] = state_data_trans_S2[15 * 4 - 1: 
15 * 3];
end
always @ *
begin
    if ((addr_S2_f[39:6+8] == tag_data_way_S2[0]) && 
(state_way_S2[0][12:11] == 2'b10 || state_way_S2[0][12:11] == 2'b11 ))
    begin
        tag_hit_way_S2[0] = 1'b1;
    end
    else
    begin
        tag_hit_way_S2[0] = 1'b0;
    end
end
always @ *
begin
    if ((addr_S2_f[39:6+8] == tag_data_way_S2[1]) && 
(state_way_S2[1][12:11] == 2'b10 || state_way_S2[1][12:11] == 2'b11 ))
    begin
        tag_hit_way_S2[1] = 1'b1;
    end
    else
    begin
        tag_hit_way_S2[1] = 1'b0;
    end
end
always @ *
begin
    if ((addr_S2_f[39:6+8] == tag_data_way_S2[2]) && 
(state_way_S2[2][12:11] == 2'b10 || state_way_S2[2][12:11] == 2'b11 ))
    begin
        tag_hit_way_S2[2] = 1'b1;
    end
    else
    begin
        tag_hit_way_S2[2] = 1'b0;
    end
end
always @ *
begin
    if ((addr_S2_f[39:6+8] == tag_data_way_S2[3]) && 
(state_way_S2[3][12:11] == 2'b10 || state_way_S2[3][12:11] == 2'b11 ))
    begin
        tag_hit_way_S2[3] = 1'b1;
    end
    else
    begin
        tag_hit_way_S2[3] = 1'b0;
    end
end
wire l2_tag_cmp_hit_S2;
l2_priority_encoder_2 priority_encoder_tag_cmp_2bits( 
    .data_in        (tag_hit_way_S2),
    .data_out       (l2_hit_way_sel_S2),
    .data_out_mask  (),
    .nonzero_out    (l2_tag_cmp_hit_S2)
);
always @ *
begin
    if (special_addr_type_S2 || msg_type_S2 == 8'd34)
    begin
        l2_tag_hit_S2 = 1'b0;
    end
    else
    begin
        l2_tag_hit_S2 = l2_tag_cmp_hit_S2;
    end
end
 
always @ *
begin
     if (!state_way_S2[0][12:11]) 
        begin
            l2_evict_way_sel_S2 = 2'd0;
        end
     else if (!state_way_S2[1][12:11]) 
        begin
            l2_evict_way_sel_S2 = 2'd1;
        end
     else if (!state_way_S2[2][12:11]) 
        begin
            l2_evict_way_sel_S2 = 2'd2;
        end
     else if (!state_way_S2[3][12:11]) 
        begin
            l2_evict_way_sel_S2 = 2'd3;
        end
    else
    begin
    case (l2_rb_bits_S2)
    2'd0:
    begin
        if (!l2_lru_bits_S2[0])
        begin
            l2_evict_way_sel_S2 = 2'd0;
        end
        else if (!l2_lru_bits_S2[1])
        begin
            l2_evict_way_sel_S2 = 2'd1;
        end
        else if (!l2_lru_bits_S2[2])
        begin
            l2_evict_way_sel_S2 = 2'd2;
        end
        else
        begin
            l2_evict_way_sel_S2 = 2'd3;
        end
    end
    2'd1:
    begin
        if (!l2_lru_bits_S2[1])
        begin
            l2_evict_way_sel_S2 = 2'd1;
        end
        else if (!l2_lru_bits_S2[2])
        begin
            l2_evict_way_sel_S2 = 2'd2;
        end
        else if (!l2_lru_bits_S2[3])
        begin
            l2_evict_way_sel_S2 = 2'd3;
        end
        else
        begin
            l2_evict_way_sel_S2 = 2'd0;
        end
    end
    2'd2:
    begin
        if (!l2_lru_bits_S2[2])
        begin
            l2_evict_way_sel_S2 = 2'd2;
        end
        else if (!l2_lru_bits_S2[3])
        begin
            l2_evict_way_sel_S2 = 2'd3;
        end
        else if (!l2_lru_bits_S2[0])
        begin
            l2_evict_way_sel_S2 = 2'd0;
        end
        else
        begin
            l2_evict_way_sel_S2 = 2'd1;
        end
    end
    2'd3:
    begin
        if (!l2_lru_bits_S2[3])
        begin
            l2_evict_way_sel_S2 = 2'd3;
        end
        else if (!l2_lru_bits_S2[0])
        begin
            l2_evict_way_sel_S2 = 2'd0;
        end
        else if (!l2_lru_bits_S2[1])
        begin
            l2_evict_way_sel_S2 = 2'd1;
        end
        else
        begin
            l2_evict_way_sel_S2 = 2'd2;
        end
    end
    default:
    begin
        l2_evict_way_sel_S2 = 2'd0;
    end
    endcase
    end
end
always @ *
begin
    if (special_addr_type_S2 || msg_type_S2 == 8'd34)
    begin
        l2_way_sel_S2 = addr_S2[6+8+2-1:6+8];
    end
    else if (l2_tag_hit_S2)
    begin
        l2_way_sel_S2 = l2_hit_way_sel_S2;
    end
    else   
    begin
        l2_way_sel_S2 = l2_evict_way_sel_S2;
    end
end
always @ *
begin
    if (special_addr_type_S2 
     || msg_type_S2 == 8'd13
     || msg_type_S2 == 8'd15)
    begin
        l2_evict_S2 = 1'b0;
    end
    else if (!l2_tag_hit_S2 && (state_way_S2[l2_way_sel_S2][12:11] == 2'b10 || 
        state_way_S2[l2_way_sel_S2][12:11] == 2'b11))
    begin
        l2_evict_S2 = 1'b1;
    end
    else
    begin
        l2_evict_S2 = 1'b0;
    end
end
always @ *
begin
    if (special_addr_type_S2
     || msg_type_S2 == 8'd13)
    begin
        l2_wb_S2 = 1'b0;
    end
    else if (((!l2_tag_hit_S2 && (msg_type_S2 != 8'd15))
           || (msg_type_S2 == 8'd14 || msg_type_S2 == 8'd35)
           || (l2_tag_hit_S2 && msg_type_S2 == 8'd15))
    && (state_way_S2[l2_way_sel_S2][14:13] == 2'b00)
    && (state_way_S2[l2_way_sel_S2][12:11] == 2'b11))
    begin
        l2_wb_S2 = 1'b1;
    end
    else
    begin
        l2_wb_S2 = 1'b0;
    end
end
reg [6-1:0] l2_way_state_owner_S2;
always @ *
begin
    l2_way_state_mesi_S2 = state_way_S2[l2_way_sel_S2][14:13];
    l2_way_state_vd_S2 = state_way_S2[l2_way_sel_S2][12:11];
    l2_way_state_subline_S2 = state_way_S2[l2_way_sel_S2][9:6];
    l2_way_state_cache_type_S2 = state_way_S2[l2_way_sel_S2][10];
    l2_way_state_owner_S2 = state_way_S2[l2_way_sel_S2][5:0];
end
always @ *
begin
    
    if (csm_en)
    begin
        req_from_owner_S2 = (l2_way_state_owner_S2 == lsid_S2_f) && (lsid_S2_f != 6'd63);
    end
    else
    
    begin
        req_from_owner_S2 = (l2_way_state_owner_S2 == flat_id_S2);
    end
end
always @ *
begin
    dir_addr_S2 = {addr_S2_f[6+8-1:6],l2_way_sel_S2}; 
end
always @ *
begin
    if (l2_wb_S2)
    begin
        data_addr_S2 = {addr_S2_f[6+8-1:6],l2_way_sel_S2, l2_load_data_subline_S2};
    end
    else if (l2_ifill_32B_S2)
    begin
        data_addr_S2 = {addr_S2_f[6+8-1:6],l2_way_sel_S2, 
                        addr_S2_f[5], l2_load_data_subline_S2[0]};
    end
    else
    begin
        data_addr_S2 = {addr_S2_f[6+8-1:6],l2_way_sel_S2, addr_S2_f[5:4]};
    end
end
reg [40-1:0] evict_addr_S2;
always @ *
begin
    evict_addr_S2 = {tag_data_way_S2[l2_way_sel_S2], addr_S2_f[6+8-1:6], {6{1'b0}}}; 
end
always @ *
begin
    addr_l2_aligned_S2 = (addr_S2_f[6-1:0] == {6{1'b0}}); 
end
always @ *
begin
    if (special_addr_type_S2)
    begin  
        if (addr_S2[39:32] == 8'ha4)
        begin
            return_data_S2 = {{(64 - 26){1'b0}}, tag_data_way_S2[l2_way_sel_S2]};
        end
        else if (addr_S2[39:32] == 8'ha6)
        begin
        
            if (addr_S2[31:30] == {2{1'b0}})
            begin
                return_data_S2 = {{(64 - 15*4){1'b0}}, state_data_trans_S2[15*4-1:0]};
            end
            else
            begin
                return_data_S2 = {{(64 - 2 - 4){1'b0}}, l2_rb_bits_S2, l2_lru_bits_S2};
            end
        end
        else
        begin
            return_data_S2 = {64{1'b0}};
        end 
    end
    else
    begin
        return_data_S2 = {64{1'b0}};
    end
end
always @ *
begin
    if (special_addr_type_S2)
    begin  
        dir_data_in_S2 = msg_data_S2;  
    end
    else
    begin
        
        
        if (csm_en && (dir_op_S2 == 2'd1))
        begin
            dir_data_in_S2 = {sdid_S2_f, src_chipid_S2_f, src_y_S2_f,src_x_S2_f};  
        end
        else        
        
        begin
            dir_data_in_S2 = {64{1'b1}}; 
        end 
    end
end
always @ *
begin
    if (special_addr_type_S2)
    begin  
        dir_data_mask_in_S2 = {64{1'b1}};
    end
    else
    begin
        
        if (csm_en)
        begin
            if (dir_op_S2 == 2'd1)
            begin
                dir_data_mask_in_S2 = {64{1'b1}};
            end
            else
            begin
                dir_data_mask_in_S2 = {{(64-1){1'b0}},1'b1} << lsid_S2_f;
            end
        end
        else    
        
        begin
            dir_data_mask_in_S2 = {{(64-1){1'b0}},1'b1} << flat_id_S2;
        end
    end 
end
reg [128-1:0] msg_data_mask_in_S2;
reg [128-1:0] data_data_merge_S2;
wire [8-1:0] data_data_parity1_S2;
wire [8-1:0] data_data_parity2_S2;
wire [128-1:0] amo_result_S2;
always @ *
begin
    if (data_size_S2 == 3'b001)
    begin
        msg_data_mask_in_S2 = {{8{1'b1}}, {(128-8){1'b0}}};
        msg_data_mask_in_S2 = msg_data_mask_in_S2 >> (8*addr_S2_f[3:0]);
    end
    else if (data_size_S2 == 3'b010)
    begin
        msg_data_mask_in_S2 = {{16{1'b1}}, {(128-16){1'b0}}};
        msg_data_mask_in_S2 = msg_data_mask_in_S2 >> (16*addr_S2_f[3:1]);
    end
    else if (data_size_S2 == 3'b011)
    begin
        msg_data_mask_in_S2 = {{32{1'b1}}, {(128-32){1'b0}}};
        msg_data_mask_in_S2 = msg_data_mask_in_S2 >> (32*addr_S2_f[3:2]);
    end
    else
    begin   
        msg_data_mask_in_S2 = {128{1'b1}}; 
    end
    msg_data_mask_in_S2 = {msg_data_mask_in_S2[63:0], msg_data_mask_in_S2[127:64]};
end
l2_amo_alu l2_amo_alu (
    .amo_alu_op     (amo_alu_op_S2),
    .address        (addr_S2_f),
    .data_size      (data_size_S2),
    .memory_operand (atomic_read_data_S2_f),
    .cpu_operand    ({msg_data_S2, msg_data_S2}),
    .amo_result     (amo_result_S2)
);
always @ *
begin
    data_data_merge_S2 = ({msg_data_S2, msg_data_S2} & msg_data_mask_in_S2)
                       | (atomic_read_data_S2_f & ~msg_data_mask_in_S2); 
    if (amo_alu_op_S2 != 4'd0)
    begin
        data_data_merge_S2 = amo_result_S2;
    end
end
l2_data_pgen data_pgen1( 
    .din            (data_data_merge_S2[64-1:0]),
    .parity         (data_data_parity1_S2)
);
l2_data_pgen data_pgen2( 
    .din            (data_data_merge_S2[128-1:64]),
    .parity         (data_data_parity2_S2)
);
always @ *
begin
    if (special_addr_type_S2)
    begin
        data_data_in_S2 = {msg_data_S2[8-1:0], msg_data_S2,
                           msg_data_S2[8-1:0], msg_data_S2};
    end
    else
    begin
        data_data_in_S2 = {data_data_parity2_S2, data_data_merge_S2[127:64], data_data_parity1_S2, data_data_merge_S2[63:0]}; 
    end
end
always @ *
begin
    if (special_addr_type_S2)
    begin
        if (addr_S2_f[31:30] == {2{1'b0}})
        begin
            data_data_mask_in_S2 = {{(144-72){1'b0}},
                                    {8{1'b0}}, {64{1'b1}}};
        end
        else
        begin
            data_data_mask_in_S2 = {{(144-72){1'b0}},
                                    {8{1'b1}}, {64{1'b0}}};
        end
        data_data_mask_in_S2 = data_data_mask_in_S2 << (72*addr_S2_f[3]);
    end
    else if (data_size_S2 == 3'b001 || data_size_S2 == 3'b010
    ||  data_size_S2 == 3'b011 || data_size_S2 == 3'b100
    )
    begin
        data_data_mask_in_S2 = {{(144-72){1'b0}},{72{1'b1}}};
        data_data_mask_in_S2 = data_data_mask_in_S2 << (72*addr_S2_f[3]);
    end
    else
    begin   
        data_data_mask_in_S2 = {144{1'b1}}; 
    end
end
reg [6-1:0] state_owner_S2;
reg [4-1:0] state_subline_S2;
reg [2-1:0] state_rb_S2;
reg [4-1:0] state_lru_S2;
always @ *
begin
    state_owner_S2 = l2_way_state_owner_S2; 
    if (state_owner_op_S2 == 2'd1)
    begin
        
        if (csm_en)
        begin
            if (state_load_sdid_S2)
            begin
                state_owner_S2 = sdid_S2_f[5:0];
            end
            else
            begin
                state_owner_S2 = lsid_S2_f; 
            end
        end
        else
        
        begin
            state_owner_S2 = flat_id_S2; 
        end
    end
    else if (state_owner_op_S2 == 2'd2)
    begin
        state_owner_S2 = l2_way_state_owner_S2 + 1; 
    end
    else if (state_owner_op_S2 == 2'd3)
    begin
        state_owner_S2 = l2_way_state_owner_S2 - 1; 
    end
    else if (state_owner_op_S2 == 2'd0)
    begin
        state_owner_S2 = 0; 
    end
end
reg [4-1:0] addr_subline_S2;
always @ *
begin
    if (cache_type_S2 == 1'b0)
    begin
        
        addr_subline_S2= {{(4-1){1'b0}},1'b1} << addr_S2_f[5:4];
    end
    else
    begin
        addr_subline_S2= {{(4-2){1'b0}},2'b11} << (2*addr_S2_f[5]);
        
    end
end
always @ *
begin
    if (state_load_sdid_S2)
    begin
        state_subline_S2 = sdid_S2_f[9:6];
    end
    else if (state_subline_op_S2 == 2'd2)
    begin
        state_subline_S2 = l2_way_state_subline_S2 | addr_subline_S2;
    end
    else if (state_subline_op_S2 == 2'd3)
    begin
        state_subline_S2 = l2_way_state_subline_S2 & (~addr_subline_S2);
    end
    else if (state_subline_op_S2 == 2'd0)
    begin
        state_subline_S2 = {4{1'b0}};
    end
    else
    begin
        state_subline_S2 = {4{1'bx}};
    end
end
always @ *
begin
    state_rb_S2 = l2_rb_bits_S2 + 1; 
end
always @ *
begin
    if (state_lru_en_S2)
    begin
        if (state_lru_op_S2 == 1'b0)
        begin
            state_lru_S2 = l2_lru_bits_S2 & (~({{(4-1){1'b0}},1'b1} << l2_way_sel_S2));
        end
        else
        begin
            state_lru_S2 = l2_lru_bits_S2 | ({{(4-1){1'b0}},1'b1} << l2_way_sel_S2);
            
            if (state_lru_S2 == {4{1'b1}})
            begin
                state_lru_S2 = {4{1'b0}};
            end
        end
    end
    else
    begin
        state_lru_S2 = l2_lru_bits_S2; 
    end
end
always @ *
begin
    if (special_addr_type_S2)
    begin   
        state_data_in_S2 = {msg_data_S2[2+4-1:0], msg_data_S2[15*4-1:0]};
    end
    else
    begin
        state_data_in_S2 = {state_rb_S2, state_lru_S2, 
        {4{state_mesi_S2, state_vd_S2, cache_type_S2, state_subline_S2, state_owner_S2}}};
    end
end
reg [15*4-1:0] state_way_data_mask_in_S2;
always @ *
begin
    state_way_data_mask_in_S2 = {{(4-1)*15{1'b0}},
                                {{2{state_mesi_en_S2}}, 
                                 {2{state_vd_en_S2}}, 
                                 {1{state_di_en_S2}}, 
                                 {4{state_subline_en_S2}}, 
                                 {6{state_owner_en_S2}}}} 
    << (l2_way_sel_S2 * 15); 
end
always @ *
begin
    if (special_addr_type_S2)
    begin
        if (addr_S2_f[31:30] == {2{1'b0}})
        begin
            state_data_mask_in_S2 = {{(2+4){1'b0}}, {15*4{1'b1}}};
        end
        else
        begin
            state_data_mask_in_S2 = {{(2+4){1'b1}}, {15*4{1'b0}}};
        end
    end
    else
    begin
        state_data_mask_in_S2 = {{2{state_rb_en_S2}}, 
                                {4{state_lru_en_S2}},
                                state_way_data_mask_in_S2}; 
    end
end
reg [64-1:0] msg_data_S2_next;
always @ *
begin
    if (special_addr_type_S2)
    begin
        msg_data_S2_next = return_data_S2;
    end
    else
    begin
        msg_data_S2_next = msg_data_S2;
    end
end
always @ *
begin
    smc_wr_addr_in_S2 = addr_S2[16+3:4];
end
always @ *
begin
    smc_data_in_S2 = {msg_data_S2, msg_data_S2};
end
reg [40-1:0] addr_S3_f;
reg [8-1:0] mshrid_S3_f;
reg [14-1:0] src_chipid_S3_f;
reg [8-1:0] src_x_S3_f;
reg [8-1:0] src_y_S3_f;
reg [4-1:0] src_fbits_S3_f;
reg [10-1:0] sdid_S3_f;
reg [6-1:0] lsid_S3_f;
reg [6-1:0] mshr_miss_lsid_S3_f;
reg [40-1:0] evict_addr_S3_f;
reg l2_tag_hit_S3_f;
reg l2_evict_S3_f;
reg [2-1:0] l2_way_sel_S3_f;
reg [6-1:0] l2_way_state_owner_S3_f;
reg [2-1:0] l2_way_state_mesi_S3_f;
reg [2-1:0] l2_way_state_vd_S3_f;
reg [4-1:0] l2_way_state_subline_S3_f;
reg [1-1:0] l2_way_state_cache_type_S3_f;
reg [64-1:0] msg_data_S3_f;
reg req_from_owner_S3_f;
reg [15*4+2+4-1:0] state_data_in_S3_f;
reg [15*4+2+4-1:0] state_data_mask_in_S3_f;
reg [8+2+2-1:0] data_addr_S3_f;
reg recycled_S3_f;
reg data_clk_en_S3_f; 
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        addr_S3_f <= 0;
        mshrid_S3_f <= 0;
        src_chipid_S3_f <= 0;
        src_x_S3_f <= 0;
        src_y_S3_f <= 0;
        src_fbits_S3_f <= 0;
        sdid_S3_f <= 0;
        lsid_S3_f <= 0;
        mshr_miss_lsid_S3_f <= 0;
        evict_addr_S3_f <= 0;
        l2_tag_hit_S3_f <= 0;
        l2_evict_S3_f <= 0;
        l2_way_sel_S3_f <= 0;
        l2_way_state_owner_S3_f <= 0;
        l2_way_state_mesi_S3_f <= 0;
        l2_way_state_vd_S3_f <= 0;
        l2_way_state_subline_S3_f <= 0;
        l2_way_state_cache_type_S3_f <= 0;
        msg_data_S3_f <= 0;
        req_from_owner_S3_f <= 0; 
        state_data_in_S3_f <= 0;
        state_data_mask_in_S3_f <= 0;
        data_addr_S3_f <= 0;
        recycled_S3_f <= 0;
        data_clk_en_S3_f <= 0;
    end
    else if (!stall_S3)
    begin
        addr_S3_f <= addr_S2;
        mshrid_S3_f <= mshrid_S2_f;
        src_chipid_S3_f <= src_chipid_S2_f;
        src_x_S3_f <= src_x_S2_f;
        src_y_S3_f <= src_y_S2_f;
        src_fbits_S3_f <= src_fbits_S2_f;
        sdid_S3_f <= sdid_S2_f;
        lsid_S3_f <= lsid_S2_f;
        mshr_miss_lsid_S3_f <= mshr_miss_lsid_S2_f;
        evict_addr_S3_f <= evict_addr_S2;
        l2_tag_hit_S3_f <= l2_tag_hit_S2;
        l2_evict_S3_f <= l2_evict_S2;
        l2_way_sel_S3_f <= l2_way_sel_S2;
        l2_way_state_owner_S3_f <= l2_way_state_owner_S2;
        l2_way_state_mesi_S3_f <= l2_way_state_mesi_S2;
        l2_way_state_vd_S3_f <= l2_way_state_vd_S2;
        l2_way_state_subline_S3_f <= l2_way_state_subline_S2;
        l2_way_state_cache_type_S3_f <= l2_way_state_cache_type_S2;
        msg_data_S3_f <= msg_data_S2_next;
        req_from_owner_S3_f <= req_from_owner_S2; 
        state_data_in_S3_f <= state_data_in_S2;
        state_data_mask_in_S3_f <= state_data_mask_in_S2;
        data_addr_S3_f <= data_addr_S2;
        recycled_S3_f <= recycled_S2_f;
    end
    data_clk_en_S3_f <= (data_clk_en_S2 && valid_S2 && !stall_real_S2); 
end
always @ *
begin
    addr_S3 = addr_S3_f;
end
reg [40-1:0] addr_S4_f;
reg [8-1:0] mshrid_S4_f;
reg [14-1:0] src_chipid_S4_f;
reg [8-1:0] src_x_S4_f;
reg [8-1:0] src_y_S4_f;
reg [4-1:0] src_fbits_S4_f;
reg [10-1:0] sdid_S4_f;
reg [6-1:0] lsid_S4_f;
reg [6-1:0] mshr_miss_lsid_S4_f;
reg [40-1:0] evict_addr_S4_f;
reg l2_tag_hit_S4_f;
reg l2_evict_S4_f;
reg [2-1:0] l2_way_sel_S4_f;
reg [6-1:0] l2_way_state_owner_S4_f;
reg [2-1:0] l2_way_state_mesi_S4_f;
reg [2-1:0] l2_way_state_vd_S4_f;
reg [4-1:0] l2_way_state_subline_S4_f;
reg [1-1:0] l2_way_state_cache_type_S4_f;
reg [64-1:0] msg_data_S4_f;
reg req_from_owner_S4_f;
reg [15*4+2+4-1:0] state_data_in_S4_f;
reg [15*4+2+4-1:0] state_data_mask_in_S4_f;
reg [144-1:0] data_data_S4_f;
reg [8+2+2-1:0] data_addr_S4_f;
reg recycled_S4_f;
reg data_stalled_skid_buffer_en_S3_f;
reg [144-1:0] data_stalled_skid_buffer_S3_f;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        addr_S4_f <= 0;
        mshrid_S4_f <= 0;
        src_chipid_S4_f <= 0;
        src_x_S4_f <= 0;
        src_y_S4_f <= 0;
        src_fbits_S4_f <= 0;
        sdid_S4_f <= 0;
        lsid_S4_f <= 0;
        mshr_miss_lsid_S4_f <= 0;
        evict_addr_S4_f <= 0;
        l2_tag_hit_S4_f <= 0;
        l2_evict_S4_f <= 0;
        l2_way_sel_S4_f <= 0;
        l2_way_state_owner_S4_f <= 0;
        l2_way_state_mesi_S4_f <= 0;
        l2_way_state_vd_S4_f <= 0;
        l2_way_state_subline_S4_f <= 0;
        l2_way_state_cache_type_S4_f <= 0;
        msg_data_S4_f <= 0;
        req_from_owner_S4_f <= 0; 
        state_data_in_S4_f <= 0;
        state_data_mask_in_S4_f <= 0;
        data_data_S4_f <= 0;
        data_addr_S4_f <= 0;
        recycled_S4_f <= 0;
    end
    else if (!stall_S4)
    begin
        addr_S4_f <= addr_S3_f;
        mshrid_S4_f <= mshrid_S3_f;
        src_chipid_S4_f <= src_chipid_S3_f;
        src_x_S4_f <= src_x_S3_f;
        src_y_S4_f <= src_y_S3_f;
        src_fbits_S4_f <= src_fbits_S3_f;
        sdid_S4_f <= sdid_S3_f;
        lsid_S4_f <= lsid_S3_f;
        mshr_miss_lsid_S4_f <= mshr_miss_lsid_S3_f;
        evict_addr_S4_f <= evict_addr_S3_f;
        l2_tag_hit_S4_f <= l2_tag_hit_S3_f;
        l2_evict_S4_f <= l2_evict_S3_f;
        l2_way_sel_S4_f <= l2_way_sel_S3_f;
        l2_way_state_owner_S4_f <= l2_way_state_owner_S3_f;
        l2_way_state_mesi_S4_f <= l2_way_state_mesi_S3_f;
        l2_way_state_vd_S4_f <= l2_way_state_vd_S3_f;
        l2_way_state_subline_S4_f <= l2_way_state_subline_S3_f;
        l2_way_state_cache_type_S4_f <= l2_way_state_cache_type_S3_f;
        msg_data_S4_f <= msg_data_S3_f;
        req_from_owner_S4_f <= req_from_owner_S3_f; 
        state_data_in_S4_f <= state_data_in_S3_f;
        state_data_mask_in_S4_f <= state_data_mask_in_S3_f;
        data_data_S4_f <= data_data_S3;
        data_addr_S4_f <= data_addr_S3_f;
        recycled_S4_f <= recycled_S3_f;
        if (data_stalled_skid_buffer_en_S3_f) begin
            data_data_S4_f <= data_stalled_skid_buffer_S3_f;
        end
    end
end
wire data_stalled_skid_buffer_en_S3 = data_clk_en_S3_f && valid_S3 && stall_S3;
wire data_stalled_skid_buffer_consume_S3 = valid_S3 && !stall_S3;
always @ (posedge clk) begin
    if (data_stalled_skid_buffer_en_S3) begin
        data_stalled_skid_buffer_S3_f <= data_data_S3;
        data_stalled_skid_buffer_en_S3_f <= 1'b1;
    end
    if (data_stalled_skid_buffer_consume_S3) begin
        data_stalled_skid_buffer_en_S3_f <= 1'b0;
    end
end
 
reg [15*4+2+4-1:0] state_data_in_real_S4;
reg [15*4+2+4-1:0] state_data_mask_in_real_S4;
reg [16-1:0] smc_rd_addr_in_S4;
reg [144-1:0] data_data_S4;
reg [10-1:0] sdid_S4;
always @ *
begin
    addr_S4 = addr_S4_f;
    mshrid_S4 = mshrid_S4_f;
    l2_evict_S4 = l2_evict_S4_f;
    l2_tag_hit_S4 = l2_tag_hit_S4_f;
    l2_way_state_mesi_S4 = l2_way_state_mesi_S4_f;
    l2_way_state_owner_S4 = l2_way_state_owner_S4_f;
    l2_way_state_vd_S4 = l2_way_state_vd_S4_f;
    l2_way_state_subline_S4 = l2_way_state_subline_S4_f; 
    l2_way_state_cache_type_S4 = l2_way_state_cache_type_S4_f;
    mshr_miss_lsid_S4 = mshr_miss_lsid_S4_f;
    lsid_S4 = lsid_S4_f;
    data_data_S4 = data_data_S4_f;
    data_addr_S4 = data_addr_S4_f;
end
always @ *
begin
    
    if (csm_en && (!msg_from_mshr_S4 || recycled_S4_f) && l2_evict_S4)
    begin
        if (l2_way_state_mesi_S4 == 2'b10)
        begin
            sdid_S4 = dir_data_S4[14+8+8+10-1:14+8+8]; 
        end
        else if (l2_way_state_mesi_S4 == 2'b01 || l2_way_state_mesi_S4 == 2'b11)
        begin
            sdid_S4 = {l2_way_state_subline_S4, l2_way_state_owner_S4};
        end
        else
        begin
            sdid_S4 = sdid_S4_f;
        end
    end
    else
    
    begin
        sdid_S4 = sdid_S4_f;
    end
end
always @ *
begin
    
    if (csm_en && (msg_type_S4 == 8'd13) && l2_tag_hit_S4
     && (l2_way_state_mesi_S4 == 2'b10) && l2_way_state_subline_S4[addr_S4[5:4]])
    begin
        req_from_owner_S4 = (src_chipid_S4_f == dir_data_S4[29:16])
                         && (src_x_S4_f == dir_data_S4[7:0])
                         && (src_y_S4_f == dir_data_S4[15:8]);
    end
    else
    
    begin
        req_from_owner_S4 = req_from_owner_S4_f;
    end
end
reg [16-1:0] smc_rd_addr_in_buf_S4_next;
reg [16-1:0] smc_rd_addr_in_buf_S4_f;
always @ *
begin
    if (!rst_n)
    begin
        smc_rd_addr_in_buf_S4_next = 0;
    end
    else if (!stall_smc_buf_S4)
    begin
        smc_rd_addr_in_buf_S4_next = smc_rd_addr_in_S4;
    end
    else 
    begin
        smc_rd_addr_in_buf_S4_next = smc_rd_addr_in_buf_S4_f;
    end
end
always @ (posedge clk)
begin
    smc_rd_addr_in_buf_S4_f <= smc_rd_addr_in_buf_S4_next;
end
always @ *
begin
    smc_rd_addr_in_buf_S4 = smc_rd_addr_in_buf_S4_f;
end
always @ *
begin
    state_wr_addr_S4 = addr_S4_f[6+8-1:6]; 
end
always @ *
begin
    
    
    
    
    if(!msg_from_mshr_S4 || recycled_S4_f)
    begin
        
        if (smc_miss_S4)
        begin
            state_data_in_real_S4 = {{2{1'b0}}, {4{1'b0}}, 
            {4{{2{1'b0}}, {2{1'b0}}, {1{1'b0}}, {4{1'b0}}, 
            (dir_sharer_counter_S4 - mshr_inv_counter_out_S4 - 6'b1)}}};
        end
        else
        
        begin
            state_data_in_real_S4 = {{2{1'b0}}, {4{1'b0}}, 
            {4{{2{1'b0}}, {2{1'b0}}, {1{1'b0}}, {4{1'b0}}, 
            (dir_sharer_counter_S4 - mshr_inv_counter_out_S4)}}};
        end
    end
    else
    begin
        
        if (smc_miss_S4)
        begin
            state_data_in_real_S4 = {{2{1'b0}}, {4{1'b0}}, 
            {4{{2{1'b0}}, {2{1'b0}}, {1{1'b0}}, {4{1'b0}}, 
            (dir_sharer_counter_S4 + l2_way_state_owner_S4_f - mshr_inv_counter_out_S4 - 6'b1)}}};
        end
        else
        
        begin
            state_data_in_real_S4 = {{2{1'b0}}, {4{1'b0}}, 
            {4{{2{1'b0}}, {2{1'b0}}, {1{1'b0}}, {4{1'b0}}, 
            (dir_sharer_counter_S4 + l2_way_state_owner_S4_f - mshr_inv_counter_out_S4)}}};
        end
    end
end
reg [4*15-1:0] state_way_data_mask_in_S4;
always @ *
begin
    state_way_data_mask_in_S4 = {{(4-1)*15{1'b0}},
                                {{2{1'b0}}, 
                                 {2{1'b0}}, 
                                 {1{1'b0}}, 
                                 {4{1'b0}}, 
                                 {6{state_wr_sel_S4}}}} 
    << (l2_way_sel_S4_f * 15); 
end
always @ *
begin
    state_data_mask_in_real_S4 = {{2{1'b0}}, 
                                 {4{1'b0}},
                                 state_way_data_mask_in_S4}; 
end
always @ *
begin
    state_data_mask_in_S4 = state_data_mask_in_S4_f | state_data_mask_in_real_S4;
end
always @ *
begin
    state_data_in_S4 = (state_data_in_S4_f & state_data_mask_in_S4_f) | 
                       (state_data_in_real_S4 & state_data_mask_in_real_S4);
end
reg [144-1:0] data_data_buf_S4_f;
reg [144-1:0] data_data_buf_S4_next;
reg [144-1:0] data_data_trans_S4;
reg [128-1:0] data_data_shift_S4;
wire corr_error1_S4, corr_error2_S4;
wire uncorr_error1_S4, uncorr_error2_S4;
always @ *
begin
    if (!rst_n)
    begin
        data_data_buf_S4_next = 0;
    end
    else if (stall_S4 && !stall_before_S4)
    begin
        data_data_buf_S4_next = data_data_S4;
    end
    else
    begin
        data_data_buf_S4_next = data_data_buf_S4_f;
    end
end
always @ (posedge clk)
begin
    data_data_buf_S4_f <= data_data_buf_S4_next;
end
always @ *
begin
    if (stall_before_S4)
    begin
        data_data_trans_S4 = data_data_buf_S4_f;
    end
    else
    begin
        data_data_trans_S4 = data_data_S4;
    end
end
l2_data_ecc data_ecc1 ( 
    .din                (data_data_trans_S4[63:0]),
    .parity             (data_data_trans_S4[71:64]),        
    .dout               (data_data_ecc_S4[63:0]),
    .corr_error         (corr_error1_S4),
    .uncorr_error       (uncorr_error1_S4)
);
l2_data_ecc data_ecc2 ( 
    .din                (data_data_trans_S4[135:72]),
    .parity             (data_data_trans_S4[143:136]),        
    .dout               (data_data_ecc_S4[127:64]),
    .corr_error         (corr_error2_S4),
    .uncorr_error       (uncorr_error2_S4)
);
always @ *
begin
    corr_error_S4 = corr_error1_S4 | corr_error2_S4; 
    uncorr_error_S4 = uncorr_error1_S4 | uncorr_error2_S4; 
end
always @ *
begin
    case (cas_cmp_data_size_S4)
    3'b011:  
    begin
        data_data_shift_S4 = {data_data_ecc_S4[63:0],data_data_ecc_S4[127:64]} << 32*addr_S4_f[3:2];
    end
    3'b100:
    begin
        data_data_shift_S4 = {data_data_ecc_S4[63:0], data_data_ecc_S4[127:64]} << 64*addr_S4_f[3];
    end
    default:
    begin
        data_data_shift_S4 = {data_data_ecc_S4[63:0], data_data_ecc_S4[127:64]};
    end
    endcase
end
always @ *
begin
    if (cas_cmp_en_S4)
    begin
    case (cas_cmp_data_size_S4)
        3'b011:  
        begin
            if (data_data_shift_S4[127:96] == msg_data_S4_f[31:0])
            begin
                cas_cmp_S4 = y;
            end
            else
            begin
                cas_cmp_S4 = n;
            end
        end
        3'b100:
        begin
            if (data_data_shift_S4[127:64] == msg_data_S4_f[63:0])
            begin
                cas_cmp_S4 = y;
            end
            else
            begin
                cas_cmp_S4 = n;
            end
        end
        default:
        begin
            cas_cmp_S4 = n;
        end
    endcase
    end
    else
    begin
        cas_cmp_S4 = n;
    end
end
always @ *
begin
    if (l2_evict_S4 
    && (msg_send_type_S4 == 8'd20
    ||  msg_send_type_S4 == 8'd18
    ||  msg_send_type_S4 == 8'd17))
    begin
        msg_send_addr_S4 = evict_addr_S4_f;
    end
    else if (msg_send_type_S4 == 8'd17
         ||  msg_send_type_S4 == 8'd18
         ||  msg_send_type_S4 == 8'd16)
    begin
        msg_send_addr_S4 = {addr_S4_f[39:6+8], addr_S4_f[6+8-1:6], {6{1'b0}}}; 
    end
    else if (msg_send_type_S4 == 8'd14)
    begin
        
        if (csm_en)
        begin 
            if (smc_miss_S4)
            begin 
                msg_send_addr_S4 = {smt_base_addr, smc_rd_addr_in_S4[15:2], 4'd0};
            end
            else
            begin
                msg_send_addr_S4 = addr_S4_f;
            end
        end
        else
        
        begin
            msg_send_addr_S4 = addr_S4_f;
        end
    end
    else    
    begin
        msg_send_addr_S4 = addr_S4_f;
    end
end
wire [(8-1) : 0] owner_x_S4; 
wire [(8-1) : 0] owner_y_S4; 
wire [(8-1) : 0] sharer_x_S4; 
wire [(8-1) : 0] sharer_y_S4; 
flat_id_to_xy owner_xy_gen(
    .flat_id            (l2_way_state_owner_S4_f),
    .x_coord            (owner_x_S4),
    .y_coord            (owner_y_S4)
);
flat_id_to_xy sharer_xy_gen(
    .flat_id            (dir_sharer_S4),
    .x_coord            (sharer_x_S4),
    .y_coord            (sharer_y_S4)
);
always @ *
begin
    case (msg_send_type_S4)
    8'd16, 8'd17: 
    begin
        
        if (csm_en)
        begin
            msg_send_dst_chipid_S4 = dir_data_S4[29:16];
            msg_send_dst_x_S4 = dir_data_S4[7:0];
            msg_send_dst_y_S4 = dir_data_S4[15:8];
        end
        else    
        
        begin
      
            msg_send_dst_chipid_S4 = my_nodeid_chipid_S4;
      
            msg_send_dst_x_S4 = owner_x_S4; 
            msg_send_dst_y_S4 = owner_y_S4;
        end
        msg_send_dst_fbits_S4 = 4'd0;
    end
    8'd18:
    begin
        
        if (csm_en)
        begin
            if (l2_way_state_mesi_S4_f == 2'b11)
            begin
                msg_send_dst_chipid_S4 = broadcast_chipid_out_S4;
                msg_send_dst_x_S4 = broadcast_x_out_S4;
                msg_send_dst_y_S4 = broadcast_y_out_S4;
            end
            else
            begin
                msg_send_dst_chipid_S4 = smc_data_out_S4[29:16];
                msg_send_dst_x_S4 = smc_data_out_S4[7:0];
                msg_send_dst_y_S4 = smc_data_out_S4[15:8];
            end
        end
        else
        
        begin
            msg_send_dst_chipid_S4 = my_nodeid_chipid_S4;
            msg_send_dst_x_S4 = sharer_x_S4; 
            msg_send_dst_y_S4 = sharer_y_S4;
        end
        msg_send_dst_fbits_S4 = 4'd0;
    end
    8'd28, 8'd29:
    begin
        msg_send_dst_chipid_S4 = src_chipid_S4_f;
        msg_send_dst_x_S4 = src_x_S4_f; 
        msg_send_dst_y_S4 = src_y_S4_f;
        msg_send_dst_fbits_S4 = 4'd0;
    end
    8'd19, 8'd14, 8'd15, 8'd20:
    begin
        msg_send_dst_chipid_S4 = {1'b1, my_nodeid_chipid_S4[12:0]};
        msg_send_dst_x_S4 = 0; 
        msg_send_dst_y_S4 = 0;
        msg_send_dst_fbits_S4 = 4'd2;
    end
    8'd33:
    begin
        msg_send_dst_chipid_S4 = my_nodeid_chipid_S4;
        msg_send_dst_x_S4 = my_nodeid_x_S4; 
        msg_send_dst_y_S4 = my_nodeid_y_S4;
        msg_send_dst_fbits_S4 = 4'd0;
    end
    default:
    begin
        msg_send_dst_chipid_S4 = my_nodeid_chipid_S4;
        msg_send_dst_x_S4 = my_nodeid_x_S4; 
        msg_send_dst_y_S4 = my_nodeid_y_S4;
        msg_send_dst_fbits_S4 = 4'd0;
    end
    endcase
end
always @ *
begin
    if (special_addr_type_S4)
    begin  
        if (addr_S4[39:32] == 8'ha0)
        begin
            if (addr_S4[31:30] == {2{1'b0}})
            begin
                if (addr_S4[3] == 0)
                begin
                    msg_send_data_S4 = {2{data_data_trans_S4[63:0]}}; 
                end
                else
                begin
                    msg_send_data_S4 = {2{data_data_trans_S4[135:72]}}; 
                end
            end
            else
            begin
                if (addr_S4[3] == 0)
                begin
                    msg_send_data_S4 = {2{56'b0, data_data_trans_S4[71:64]}}; 
                end
                else
                begin
                    msg_send_data_S4 = {2{56'b0, data_data_trans_S4[143:136]}}; 
                end
            end
        end
        else if (addr_S4[39:32] == 8'ha1)
        begin
            msg_send_data_S4 = {2{dir_data_sel_S4}}; 
        end
        
        else if (addr_S4[39:32] == 8'ha2)
        begin
            case (addr_S4[31:30])
            2'd0:
            begin
                msg_send_data_S4 = {2{{(64-30){1'b0}}, smc_data_out_S4}}; 
            end
            2'd1:
            begin
                msg_send_data_S4 = {2{{(64-4){1'b0}}, smc_valid_out_S4}}; 
            end
            2'd2: 
            begin
                msg_send_data_S4 = {2{{(64-14){1'b0}}, smc_tag_out_S4}}; 
            end
            default:
            begin
                msg_send_data_S4 = {128{1'b0}}; 
            end
            endcase
        end
        
        else if (addr_S4[39:32] == 8'ha9 
              || addr_S4[39:32] == 8'ha7
              || addr_S4[39:32] == 8'ha8
              || addr_S4[39:32] == 8'haa
              || addr_S4[39:32] == 8'hab)
        begin
            msg_send_data_S4 = {2{reg_data_out_S4}}; 
        end
        else
        begin
            msg_send_data_S4 = {2{msg_data_S4_f}}; 
        end 
    end
    else if ((msg_type_S4 == 8'd34 || msg_type_S4 == 8'd35) 
         &&  (msg_send_type_S4 == 8'd29))
    begin
        msg_send_data_S4 = {128{1'b0}}; 
    end  
    else if (msg_send_type_S4 == 8'd15 || (msg_send_type_S4 == 8'd33))
    begin
        msg_send_data_S4 = {2{msg_data_S4_f}}; 
    end
    else    
    begin
        msg_send_data_S4 = data_data_ecc_S4;
    end
end
always @ *
begin
    if (special_addr_type_S4 && (addr_S4[39:32] == 8'ha2))
    begin
        smc_rd_addr_in_S4 = addr_S4[16+3:4];
    end
    else if (msg_send_type_pre_S4 == 8'd18)
    begin
        smc_rd_addr_in_S4 = {sdid_S4, dir_sharer_S4};
    end
    else
    begin
        smc_rd_addr_in_S4 = {sdid_S4, l2_way_state_owner_S4_f};
    end
end
always @ *
begin
    mshr_data_in_S4 = {inv_fwd_pending_S4,
                       (req_recycle_S4 && (!msg_from_mshr_S4 || recycled_S4_f)),
                       smc_miss_S4,
                       smc_rd_addr_in_S4[5:0],
                       lsid_S4_f, 
                       sdid_S4,
                       src_fbits_S4_f,
                       src_y_S4_f,
                       src_x_S4_f,
                       src_chipid_S4_f,
                       l2_miss_S4,
                       msg_type_S4,
                       data_size_S4,
                       cache_type_S4,
                       mshrid_S4_f,
                       l2_way_sel_S4_f,
                       addr_S4_f};
end
assign mshr_data_mask_in_S4 = {120+2{1'b1}}; 
endmodule
      
 
module l2_pipe2_buf_in(
    input wire clk,
    input wire rst_n,
    input wire valid_in,
    input wire [64-1:0] data_in,
    output reg ready_in,
    output reg msg_header_valid_out,
    output reg [192-1:0] msg_header_out,
    input wire msg_header_ready_out,
    output reg msg_data_valid_out,
    output reg [128-1:0] msg_data_out,
    input wire msg_data_ready_out
);
localparam msg_data_state_0F = 4'd0;
localparam msg_data_state_1F = 4'd1; 
localparam msg_data_state_2F = 4'd2;
localparam msg_data_state_4F = 4'd3;
localparam msg_data_state_8F = 4'd4;
localparam msg_state_header0 = 4'd0;
localparam msg_state_header1 = 4'd1;
localparam msg_state_header2 = 4'd2;
localparam msg_state_data0 = 4'd3;
localparam msg_state_data1 = 4'd4;
localparam msg_state_data2 = 4'd5;
localparam msg_state_data3 = 4'd6;
localparam msg_state_data4 = 4'd7;
localparam msg_state_data5 = 4'd8;
localparam msg_state_data6 = 4'd9;
localparam msg_state_data7 = 4'd10;
reg [4-1:0] msg_state_f;
reg [4-1:0] msg_state_next;
reg [4-1:0] msg_data_state_f;
reg [4-1:0] msg_data_state_next;
always @ *
begin
    if (!rst_n)
    begin
        msg_data_state_next = msg_data_state_0F;
    end
    else if((msg_state_f == msg_state_header0) && valid_in)
    begin
        if (data_in[29:22] == 8'd8)
        begin
            msg_data_state_next = msg_data_state_8F;
        end
        else if (data_in[29:22] == 8'd0)
        begin
            msg_data_state_next = msg_data_state_0F;
        end
        else    
        begin
            msg_data_state_next = msg_data_state_2F;
        end
    end
    else
    begin
        msg_data_state_next = msg_data_state_f;
    end
end
always @ (posedge clk)
begin
    msg_data_state_f <= msg_data_state_next;
end
always @ *
begin
    if (!rst_n)
    begin
        msg_state_next = msg_state_header0;
    end
    else if (valid_in && ready_in)
    begin
        if ((msg_state_f == msg_state_header0) && (data_in[21:14] != 8'd12))
        begin
            if (data_in[29:22] == 8'd0)
            begin
                msg_state_next = msg_state_header0;
            end
            else
            begin
                msg_state_next = msg_state_data0;
            end
        end
        else if ((msg_state_f == msg_state_data1) && (msg_data_state_f == msg_data_state_2F))
        begin
            msg_state_next = msg_state_header0;
        end
        else
        begin
            if (msg_state_f == msg_state_data7)
            begin
                msg_state_next = msg_state_header0;
            end
            else
            begin
                msg_state_next = msg_state_f + 4'd1;
            end
        end
    end
    else
    begin
        msg_state_next = msg_state_f;
    end 
end
always @ (posedge clk)
begin
    msg_state_f <= msg_state_next;
end
localparam msg_mux_header = 1'b0;
localparam msg_mux_data = 1'b1;
reg msg_mux_sel;
always @ *
begin
    if ((msg_state_f == msg_state_header0)
    ||  (msg_state_f == msg_state_header1)
    ||  (msg_state_f == msg_state_header2))
    begin
        msg_mux_sel = msg_mux_header;
    end
    else
        msg_mux_sel = msg_mux_data;
end
reg msg_header_valid_in;
reg [64-1:0] msg_header_in;
reg msg_header_ready_in;
reg msg_data_valid_in;
reg [64-1:0] msg_data_in;
reg msg_data_ready_in;
always @ *
begin
    if (msg_mux_sel == msg_mux_header)
    begin
        msg_header_valid_in = valid_in;
        msg_header_in = data_in;
    end
    else
    begin
        msg_header_valid_in = 0;
        msg_header_in = 0;
    end
end
always @ *
begin
    if (msg_mux_sel == msg_mux_data)
    begin
        msg_data_valid_in = valid_in;
        msg_data_in = data_in;
    end
    else
    begin
        msg_data_valid_in = 0;
        msg_data_in = 0;
    end
end
always @ *
begin
    if (msg_mux_sel == msg_mux_data)
    begin
        ready_in = msg_data_ready_in; 
    end
    else
    begin
        ready_in = msg_header_ready_in;
    end
end
reg [64-1:0] header_buf_mem_f [4-1:0];
reg header_buf_empty;
reg header_buf_full;
reg [2:0] header_buf_counter_f;
reg [2:0] header_buf_counter_next;
reg [2-1:0] header_rd_ptr_f;
reg [2-1:0] header_rd_ptr_next;
reg [2-1:0] header_rd_ptr_plus1;
reg [2-1:0] header_rd_ptr_plus2;
reg [2-1:0] header_wr_ptr_f;
reg [2-1:0] header_wr_ptr_next;
always @ *
begin
    header_buf_empty = (header_buf_counter_f == 0);
    header_buf_full = (header_buf_counter_f ==  4);
end
reg [1:0] msg_header_flits;
always @ *
begin
    msg_header_flits = 1;
    if (header_buf_mem_f[header_rd_ptr_f][21:14] == 8'd12)
    begin
        msg_header_flits = 3;
    end
    else
    begin
        msg_header_flits = 1;
    end
end
always @ *
begin
   if (!rst_n)
    begin
        header_buf_counter_next = 0;
    end
    else if ((msg_header_valid_in && msg_header_ready_in) && (msg_header_valid_out && msg_header_ready_out))
    begin
        header_buf_counter_next = header_buf_counter_f + 1 - msg_header_flits;
    end
    else if (msg_header_valid_in && msg_header_ready_in)
    begin 
        header_buf_counter_next = header_buf_counter_f + 1;
    end
    else if (msg_header_valid_out && msg_header_ready_out)
    begin 
        header_buf_counter_next = header_buf_counter_f - msg_header_flits;
    end
    else
    begin
        header_buf_counter_next = header_buf_counter_f;
    end
end
always @ (posedge clk)
begin
    header_buf_counter_f <= header_buf_counter_next;
end
always @ *
begin
    if (!rst_n)
    begin   
        header_rd_ptr_next = 0;
    end
    else if (msg_header_valid_out && msg_header_ready_out)
    begin
        header_rd_ptr_next = header_rd_ptr_f + msg_header_flits;
    end
    else
    begin
        header_rd_ptr_next = header_rd_ptr_f;
    end
end
always @ (posedge clk)
begin
    header_rd_ptr_f <= header_rd_ptr_next;
end
always @ *
begin
    if (!rst_n)
    begin   
        header_wr_ptr_next = 0;
    end
    else if (msg_header_valid_in && msg_header_ready_in)
    begin
        header_wr_ptr_next = header_wr_ptr_f + 1;
    end
    else
    begin
        header_wr_ptr_next = header_wr_ptr_f;
    end
end
always @ (posedge clk)
begin
    header_wr_ptr_f <= header_wr_ptr_next;
end
always @ *
begin
    header_rd_ptr_plus1 = header_rd_ptr_f + 1;
    header_rd_ptr_plus2 = header_rd_ptr_f + 2;
end
always @ *
begin
   msg_header_ready_in = !header_buf_full;
end
always @ *
begin
    msg_header_valid_out = (!header_buf_empty) && (header_buf_counter_f >= msg_header_flits);
end
always @ *
begin
    if (msg_header_flits == 3)
    begin
        msg_header_out = {header_buf_mem_f[header_rd_ptr_plus2], 
                          header_buf_mem_f[header_rd_ptr_plus1], 
                          header_buf_mem_f[header_rd_ptr_f]};
    end
    else
    begin
        msg_header_out = {{(2*64){1'b0}},header_buf_mem_f[header_rd_ptr_f]}; 
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin   
        header_buf_mem_f[0] <= 0;
        header_buf_mem_f[1] <= 0;
        header_buf_mem_f[2] <= 0;
        header_buf_mem_f[3] <= 0;
    end
    else if (msg_header_valid_in && msg_header_ready_in)
    begin
        header_buf_mem_f[header_wr_ptr_f] <= msg_header_in;
    end
    else
    begin 
        header_buf_mem_f[header_wr_ptr_f] <= header_buf_mem_f[header_wr_ptr_f];
    end
end
reg [64-1:0] data_buf_mem_f [16-1:0];
reg data_buf_empty;
reg data_buf_full;
reg [4:0] data_buf_counter_f;
reg [4:0] data_buf_counter_next;
reg [4-1:0] data_rd_ptr_f;
reg [4-1:0] data_rd_ptr_next;
reg [4-1:0] data_rd_ptr_plus1;
reg [4-1:0] data_wr_ptr_f;
reg [4-1:0] data_wr_ptr_next;
reg [4-1:0] data_wr_ptr_plus1;
always @ *
begin
    data_buf_empty = (data_buf_counter_f == 0);
    data_buf_full = (data_buf_counter_f ==  16);
end
always @ *
begin
    if ((msg_data_valid_in && msg_data_ready_in) && (msg_data_valid_out && msg_data_ready_out))
    begin
        data_buf_counter_next = data_buf_counter_f + 1 - 2;
    end
    else if (msg_data_valid_in && msg_data_ready_in)
    begin 
        data_buf_counter_next = data_buf_counter_f + 1;
    end
    else if (msg_data_valid_out && msg_data_ready_out)
    begin 
        data_buf_counter_next = data_buf_counter_f - 2;
    end
    else
    begin
        data_buf_counter_next = data_buf_counter_f;
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
        data_buf_counter_f <= 0;
    else
        data_buf_counter_f <= data_buf_counter_next;
end
always @ *
begin
    if (!rst_n)
    begin   
        data_rd_ptr_next = 0;
    end
    else if (msg_data_valid_out && msg_data_ready_out)
    begin
        data_rd_ptr_next = data_rd_ptr_f + 2;
    end
    else
    begin
        data_rd_ptr_next = data_rd_ptr_f;
    end
end
always @ (posedge clk)
begin
    data_rd_ptr_f <= data_rd_ptr_next;
end
always @ *
begin
    if (!rst_n)
    begin   
        data_wr_ptr_next = 0;
    end
    else if (msg_data_valid_in && msg_data_ready_in)
    begin
        data_wr_ptr_next = data_wr_ptr_f + 1;
    end
    else
    begin
        data_wr_ptr_next = data_wr_ptr_f;
    end
end
always @ (posedge clk)
begin
    data_wr_ptr_f <= data_wr_ptr_next;
end
always @ *
begin
    data_rd_ptr_plus1 = data_rd_ptr_f + 1;
end
always @ *
begin
   msg_data_ready_in = !data_buf_full;
end
always @ *
begin
    msg_data_valid_out = (data_buf_counter_f >= 2);
    msg_data_out = {data_buf_mem_f[data_rd_ptr_plus1], data_buf_mem_f[data_rd_ptr_f]}; 
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin   
        data_buf_mem_f[0] <= 0;
        data_buf_mem_f[1] <= 0;
        data_buf_mem_f[2] <= 0;
        data_buf_mem_f[3] <= 0;
        data_buf_mem_f[4] <= 0;
        data_buf_mem_f[5] <= 0;
        data_buf_mem_f[6] <= 0;
        data_buf_mem_f[7] <= 0;
        data_buf_mem_f[8] <= 0;
        data_buf_mem_f[9] <= 0;
        data_buf_mem_f[10] <= 0;
        data_buf_mem_f[11] <= 0;
        data_buf_mem_f[12] <= 0;
        data_buf_mem_f[13] <= 0;
        data_buf_mem_f[14] <= 0;
        data_buf_mem_f[15] <= 0;
    end
    else if (msg_data_valid_in && msg_data_ready_in)
    begin
        data_buf_mem_f[data_wr_ptr_f] <= msg_data_in;
    end
    else
    begin 
        data_buf_mem_f[data_wr_ptr_f] <=  data_buf_mem_f[data_wr_ptr_f];
    end
end
endmodule
      
 
module l2_pipe2_ctrl(
    input wire clk,
    input wire rst_n,
    
    input wire csm_en,
    
    
 
    input wire msg_header_valid_S1,
    input wire [8-1:0] msg_type_S1,
    input wire [8-1:0] msg_length_S1,
    input wire [3-1:0] msg_data_size_S1,
    input wire [1-1:0] msg_cache_type_S1,
    input wire [1-1:0] msg_last_subline_S1,
    input wire [2-1:0] msg_mesi_S1,
    
    input wire [8-1:0] mshr_msg_type_S1,
    input wire [1-1:0] mshr_l2_miss_S1,
    input wire [3-1:0] mshr_data_size_S1,
    input wire [1-1:0] mshr_cache_type_S1, 
    
    input wire mshr_smc_miss_S1,
    
    input wire [2-1:0] mshr_state_out_S1,
    input wire mshr_inv_fwd_pending_S1,
    input wire [40-1:0] addr_S1,
    input wire is_same_address_S1,
    
   
 
    input wire l2_tag_hit_S2,
    input wire [2-1:0] l2_way_sel_S2,
    input wire l2_wb_S2,
    input wire [6-1:0] l2_way_state_owner_S2,
    input wire [2-1:0] l2_way_state_mesi_S2,
    input wire [2-1:0] l2_way_state_vd_S2,
    input wire [4-1:0] l2_way_state_subline_S2,
    input wire [1-1:0] l2_way_state_cache_type_S2,
    input wire addr_l2_aligned_S2,
    input wire subline_valid_S2,
    input wire [6-1:0] lsid_S2,
    
    input wire broadcast_counter_zero_S2,
    input wire broadcast_counter_max_S2,
    input wire [14-1:0] broadcast_chipid_out_S2,
    input wire [8-1:0] broadcast_x_out_S2,
    input wire [8-1:0] broadcast_y_out_S2,
    
    input wire msg_data_valid_S2,
    
    input wire [40-1:0] addr_S2,
    
    input wire [40-1:0] addr_S3,
    
    output reg valid_S1,  
    output reg stall_S1,
    output reg active_S1, 
    output reg msg_from_mshr_S1, 
 
    output reg mshr_rd_en_S1,
    
    output reg msg_header_ready_S1,
    output reg tag_clk_en_S1,
    output reg tag_rdw_en_S1,
    output reg state_rd_en_S1,
    
    output reg valid_S2,    
    output reg stall_S2,  
    output reg stall_before_S2,
    output reg active_S2, 
    output reg msg_from_mshr_S2,
    output reg [8-1:0] msg_type_S2,
    output reg [3-1:0] data_size_S2,
    output reg [1-1:0] cache_type_S2,
    output reg dir_clk_en_S2,
    output reg dir_rdw_en_S2,
    output reg dir_clr_en_S2,
    output reg data_clk_en_S2,
    output wire data_rdw_en_S2,
    
    output reg [2-1:0] broadcast_counter_op_S2,
    output reg broadcast_counter_op_val_S2,
    
    output reg state_owner_en_S2,
    output reg [2-1:0] state_owner_op_S2,
    output reg state_subline_en_S2,
    output reg [2-1:0] state_subline_op_S2,
    output reg state_di_en_S2,
    output reg state_vd_en_S2,
    output reg [2-1:0] state_vd_S2,
    output reg state_mesi_en_S2,
    output reg [2-1:0] state_mesi_S2,
    output reg state_lru_en_S2,
    output reg [1-1:0] state_lru_op_S2,
    output wire state_rb_en_S2,
    output reg l2_load_64B_S2, 
    output reg l2_load_32B_S2, 
    output reg [2-1:0] l2_load_data_subline_S2,
    output reg msg_data_ready_S2,
    
    output reg smc_wr_en_S2,
    
    
    output reg valid_S3,    
    output wire stall_S3,  
    output reg active_S3, 
    output reg [8-1:0] msg_type_S3,
    output reg mshr_wr_state_en_S3,
    output wire mshr_wr_data_en_S3,
    output reg [2-1:0] mshr_state_in_S3,
    output reg mshr_inc_counter_en_S3,
    output reg state_wr_en_S3
);
localparam y = 1'b1;
localparam n = 1'b0;
localparam rd = 1'b1;
localparam wr = 1'b0;
reg stall_pre_S1;
reg [3-1:0] data_size_S1;
reg [1-1:0] cache_type_S1;
reg smc_miss_S1;
reg inv_fwd_pending_S1;
reg stall_hazard_S1;
always @ *
begin
    stall_hazard_S1 = (valid_S2 && (addr_S1[6+8-1:6] == addr_S2[6+8-1:6])) ||
                      (valid_S3 && (addr_S1[6+8-1:6] == addr_S3[6+8-1:6]));
end
always @ *
begin
    valid_S1 = msg_header_valid_S1;
end
always @ *
begin
    stall_pre_S1 = stall_S2; 
end
always @ *
begin
    mshr_rd_en_S1 = valid_S1 && (msg_type_S1 != 8'd12) && (msg_type_S1 != 8'd25);
end
always @ *
begin
    msg_from_mshr_S1 = mshr_rd_en_S1
                    && (mshr_state_out_S1 != 2'd0); 
end
always @ *
begin
    if (msg_from_mshr_S1)
    begin
        data_size_S1 = mshr_data_size_S1;
    end
    else
    begin
        data_size_S1 = msg_data_size_S1;
    end
end
always @ *
begin
    if (msg_from_mshr_S1)
    begin
        cache_type_S1 = mshr_cache_type_S1;
    end
    else
    begin
        cache_type_S1 = msg_cache_type_S1;
    end
end
always @ *
begin
    if (msg_from_mshr_S1)
    begin
        inv_fwd_pending_S1 = mshr_inv_fwd_pending_S1;
    end
    else
    begin
        inv_fwd_pending_S1 = 1'b0;
    end
end
reg [3-1:0] cs_S1;
always @ *
begin
    cs_S1 = {3{1'bx}};
    if (valid_S1)
    begin
        case (msg_type_S1)
        8'd23:
        begin
            
            cs_S1 = {n,              rd,           y};
        end
        8'd21, 8'd22:
        begin
            cs_S1 = {n,              rd,         y};
        end
        8'd24, 8'd26:
        begin
            
            if (smc_miss_S1)
            begin
                cs_S1 = {n,              rd,           n};
            end
            else
            
            begin
                cs_S1 = {y,              wr,         n};
            end
        end
        8'd25, 8'd27:
        begin
            cs_S1 = {n,              rd,         n};
        end
        8'd12:
        begin
            cs_S1 = {y,              rd,          y};
        end
        default:
        begin
            cs_S1 = {3{1'bx}};
        end
        endcase
    end
    else
    begin
        cs_S1 = {3{1'b0}};
    end
end
always @ *
begin
    stall_S1 = valid_S1 && (stall_pre_S1 || stall_hazard_S1);
end
always @ *
begin
    msg_header_ready_S1 = !stall_S1; 
end
always @ *
begin
    tag_clk_en_S1 = valid_S1 && !stall_S1 && cs_S1[2];
end
always @ *
begin
    tag_rdw_en_S1 = valid_S1 && !stall_S1 && cs_S1[1];
end
always @ *
begin
    state_rd_en_S1 =  valid_S1 && !stall_S1 && cs_S1[0];
end
always @ *
begin
    if (msg_from_mshr_S1)
    begin
        smc_miss_S1 = mshr_smc_miss_S1;
    end
    else
    begin
        smc_miss_S1 = 0;
    end
end
reg valid_next_S1;
always @ *
begin
    valid_next_S1 = valid_S1 && !stall_S1;
end
always @ *
begin
    active_S1 = valid_S1;
end
reg valid_S2_f;
reg [8-1:0] msg_length_S2_f;
reg [1-1:0] msg_last_subline_S2_f;
reg [3-1:0] data_size_S2_f;
reg [1-1:0] cache_type_S2_f;
reg msg_from_mshr_S2_f;
reg [2-1:0] msg_mesi_S2_f;
reg smc_miss_S2_f;
reg [8-1:0] msg_type_S2_f;
reg inv_fwd_pending_S2_f;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        valid_S2_f <= 1'b0;
        msg_type_S2_f <= 0;
        msg_length_S2_f <= 0;
        msg_last_subline_S2_f <= 0;
        data_size_S2_f <= 0;  
        cache_type_S2_f <= 0; 
        msg_from_mshr_S2_f <= 1'b0;
        msg_mesi_S2_f <= 0;
        
        smc_miss_S2_f <= 0;
        
        inv_fwd_pending_S2_f <= 0;
    end
    else if (!stall_S2)
    begin
        valid_S2_f <= valid_next_S1;
        msg_type_S2_f <= msg_type_S1;
        msg_length_S2_f <= msg_length_S1;
        msg_last_subline_S2_f <= msg_last_subline_S1;
        data_size_S2_f <= data_size_S1;
        cache_type_S2_f <= cache_type_S1;
        msg_from_mshr_S2_f <= msg_from_mshr_S1;
        msg_mesi_S2_f <= msg_mesi_S1;
        
        smc_miss_S2_f <= smc_miss_S1;
        
        inv_fwd_pending_S2_f <= inv_fwd_pending_S1;
    end
end
reg stall_real_S2;
reg stall_load_S2;
reg stall_before_S2_f;
reg stall_before_S2_next;
reg state_wr_en_S2;
reg mshr_wr_state_en_S2;
reg [2-1:0] mshr_state_in_S2;
always @ *
begin
    valid_S2 = valid_S2_f;
    msg_type_S2 = msg_type_S2_f;
    msg_from_mshr_S2 = msg_from_mshr_S2_f;
    data_size_S2 = data_size_S2_f;
    cache_type_S2 = cache_type_S2_f;
    stall_before_S2 = stall_before_S2_f;
end
always @ *
begin
    if (!rst_n)
    begin
        stall_before_S2_next = 0;
    end
    else
    begin
        stall_before_S2_next = stall_S2;
    end
end
always @ (posedge clk)
begin
    stall_before_S2_f <= stall_before_S2_next;
end
reg is_last_subline_S2;
always @ *
begin
    is_last_subline_S2 = msg_last_subline_S2_f;
end
reg [19-1:0] cs_S2;
always @ *
begin
    if (valid_S2)
    begin
    case (msg_type_S2_f)
        8'd21:
        begin
            case (l2_way_state_mesi_S2)
            2'b10:
            begin
                if (is_last_subline_S2)
                begin
                    
                    if (csm_en)
                    begin
                        if (lsid_S2 == 6'd63)
                        begin
                            if (subline_valid_S2)   
                            begin
                                if (msg_length_S2_f != 0)
                                begin
                                    
                                    
                                    cs_S2 = {y,     y,         wr,         y,        y,         2'd0,     n,           2'd0,    n, 
                                    
                                    
                                             y,      2'b11,  y,      2'b11,      n,      1'b0};  
                                end     
                                else
                                begin       
                                    cs_S2 = {n,     y,         wr,         y,        y,         2'd0,     n,           2'd0,    n, 
                                             y,      2'b11,  y,      2'b11,      n,      1'b0};  
                                end
                            end
                            else
                            begin
                                cs_S2 = {n,     n,         wr,         n,       y,         2'd0,     n,           2'd0,    n, 
                                         y,      2'b11,  y,      2'b11,      n,      1'b0};    
                            end
                        end
                        else
                        begin
                            if (subline_valid_S2)   
                            begin
                                if (msg_length_S2_f != 0)
                                begin
                                    
                                    
                                    cs_S2 = {y,     y,         wr,         n,        y,         2'd1,     y,           2'd1,    n, 
                                    
                                    
                                             y,      2'b11,  y,      2'b01,      n,      1'b0};  
                                end     
                                else
                                begin       
                                    cs_S2 = {n,     y,         wr,         n,        y,         2'd1,     y,           2'd1,    n, 
                                             y,      2'b11,  y,      2'b01,      n,      1'b0};  
                                end
                            end
                            else
                            begin
                                cs_S2 = {n,     y,         wr,         n,       y,         2'd1,     y,           2'd1,    n, 
                                         y,      2'b11,  y,      2'b01,      n,      1'b0};    
                            end
                        end
                    end
                    else
                    
                    begin
                        if (subline_valid_S2)   
                        begin
                            if (msg_length_S2_f != 0)
                            begin
                                
                                
                                cs_S2 = {y,     y,         wr,         n,        y,         2'd0,     n,           2'd0,    n, 
                                
                                
                                         y,      2'b11,  y,      2'b01,      n,      1'b0};  
                            end     
                            else
                            begin       
                                cs_S2 = {n,     y,         wr,         n,        y,         2'd0,     n,           2'd0,    n, 
                                         y,      2'b11,  y,      2'b01,      n,      1'b0};  
                            end
                        end
                        else
                        begin
                            cs_S2 = {n,     y,         wr,         n,       y,         2'd0,     n,           2'd0,    n, 
                                     y,      2'b11,  y,      2'b01,      n,      1'b0};    
                        end
                    end
                end
                else
                begin
                    if (subline_valid_S2)   
                    begin
                        if (msg_length_S2_f != 0)
                        begin
                            cs_S2 = {y,     n,         rd,         n,       n,         2'd0,     n,           2'd0,    n,       
                                     n,      2'b01,  n,      2'b00,  n,      1'b0};
                        end
                        else
                        begin
                            cs_S2 = {n,     n,         rd,         n,       n,         2'd0,     n,           2'd0,    n,       
                                     n,      2'b01,  n,      2'b00,  n,      1'b0};
                        end
                    end
                    else
                    begin
                        cs_S2 = {n,     n,         rd,         n,       n,         2'd0,     n,           2'd0,    n,       
                                 n,      2'b01,  n,      2'b00,  n,      1'b0};
                    end
                end  
            end
            2'b00:
            begin
                cs_S2 = {n,     n,         rd,         n,       n,         2'd0,      n,           2'd0,    n,       
                         n,      2'b01,  n,      2'b00,  n,      1'b0};
            end
            default:
            begin
                cs_S2 = {19{1'bx}};
            end
            endcase
        end
        8'd22:
        begin
            case (l2_way_state_mesi_S2)
            2'b10:
            begin
                if (is_last_subline_S2)
                begin
                    if (subline_valid_S2)   
                    begin
                        if (msg_length_S2_f != 0)
                        begin
                            cs_S2 = {y,     y,         wr,         y,       y,         2'd0,     y,           2'd0,    n, 
                                     y,      2'b11,  y,      2'b00,      n,      1'b0};  
                        end
                        else
                        begin
                            cs_S2 = {n,     y,         wr,         y,       y,         2'd0,     y,           2'd0,    n, 
                                     y,      2'b11,  y,      2'b00,      n,      1'b0};  
                        end
                        
                    end
                    else
                    begin
                        cs_S2 = {n,     y,         wr,         y,       y,         2'd0,     y,           2'd0,    n, 
                                 y,      2'b11,  y,      2'b00,      n,      1'b0};  
                    end  
                end
                else
                begin
                    if (subline_valid_S2)   
                    begin
                        if (msg_length_S2_f != 0)
                        begin
                            cs_S2 = {y,     n,         rd,         n,       n,         2'd0,     n,           2'd0,    n,       
                                     n,      2'b01,  n,      2'b00,  n,      1'b0};
                        end
                        else
                        begin
                            cs_S2 = {n,     n,         rd,         n,       n,         2'd0,     n,           2'd0,    n,       
                                     n,      2'b01,  n,      2'b00,  n,      1'b0};
                        end
                    end
                    else
                    begin
                        cs_S2 = {n,     n,         rd,         n,       n,         2'd0,     n,           2'd0,    n,       
                                 n,      2'b01,  n,      2'b00,  n,      1'b0};
                    end 
                end 
            end
            2'b00:
            begin
                cs_S2 = {n,     n,         rd,         n,       n,         2'd0,     n,           2'd0,    n,       
                         n,      2'b01,  n,      2'b00,  n,      1'b0};
            end
            default:
            begin
                cs_S2 = {19{1'bx}};
            end
            endcase
        end
        8'd23:
        begin
            if (is_last_subline_S2)
            begin
                
                if (l2_way_state_mesi_S2 == 2'b11)
                begin   
                    if (broadcast_counter_max_S2)
                    begin
                        cs_S2 = {n,     n,         rd,         n,       y,         2'd0,     y,           2'd0,    n, 
                                 n,      2'b01,  y,      2'b00,      n,      1'b0};    
                    end
                    else
                    begin
                        cs_S2 = {n,     n,         rd,         n,       y,         2'd3,     n,           2'd0,    n, 
                                 n,      2'b01,  n,      2'b00, n,      1'b0};    
                    end
                end
                else 
                
                begin
                    
                    if ((l2_way_state_owner_S2 == 1) && (~smc_miss_S2_f) && (~inv_fwd_pending_S2_f))
                    
                    
                    begin
                        cs_S2 = {n,     n,         rd,         n,       y,         2'd0,     y,           2'd0,    n, 
                                 n,      2'b01,  y,      2'b00,      n,      1'b0};    
                    end
                    else
                    begin
                        cs_S2 = {n,     n,         rd,         n,       y,         2'd3,     n,           2'd0,    n, 
                                 n,      2'b01,  n,      2'b00, n,      1'b0};    
                    end
                end
            end
            else
            begin
                cs_S2 = {n,     n,         rd,         n,       n,         2'd0,     n,           2'd0,    n,       
                         n,      2'b01,  n,      2'b00,  n,      1'b0};
            end  
        end
        8'd24:
        begin
            cs_S2 = {y,     y,         wr,         y,       n,         2'd0,     y,           2'd0,    n,       
                     y,      2'b10,  n,      2'b00,  n,      1'b0};
        end
        8'd26:
        begin
            
            if (smc_miss_S2_f)
            begin
                cs_S2 = {n,     n,         rd,         n,       n,         2'd0,     n,           2'd0,    n,       
                         n,      2'b10,  n,      2'b00,  n,      1'b0};
            end
            else
            
            begin
                cs_S2 = {y,     n,         rd,         n,       n,         2'd0,     n,           2'd0,    n,       
                         y,      2'b10,  n,      2'b00,  n,      1'b0};
            end
        end
        8'd25, 8'd27:
        begin
            cs_S2 = {n,     n,         rd,         n,       n,         2'd0,     n,           2'd0,    n,       
                     n,      2'b01,  n,      2'b00,  n,      1'b0};
        end
        8'd12:
        begin
            begin
            
            if (l2_way_state_subline_S2 == ({{(4-1){1'b0}}, 1'b1} << addr_S2[5:4]))
            begin
                cs_S2 = {y,     y,         wr,         y,       n,         2'd0,     y,        2'd3,    n,       
                         y,     2'b11,  y,      2'b00,     n,      1'b0};
            end
            else
            begin
                cs_S2 = {y,     n,         rd,         n,       n,         2'd0,     y,        2'd3,    n,       
                         n,      2'b01,  n,      2'b00,     n,      1'b0};
            end
            end
         end
        default:
        begin
            cs_S2 = {19{1'bx}};
        end
    endcase
    end
    else    
    begin
        cs_S2 = {19{1'b0}};
    end
end
always @ *
begin
    broadcast_counter_op_val_S2 = !stall_S2 && valid_S2 && is_last_subline_S2 
                               && (msg_type_S2_f == 8'd23) && (l2_way_state_mesi_S2 == 2'b11);
end
always @ *
begin
    if (broadcast_counter_max_S2)
    begin
        broadcast_counter_op_S2 = 2'd0;
    end
    else
    begin
        broadcast_counter_op_S2 = 2'd2;
    end
end
always @ *
begin
    dir_clk_en_S2 = !stall_S2 && cs_S2[17];
end
always @ *
begin
    dir_rdw_en_S2 = cs_S2[16];
end
always @ *
begin
    dir_clr_en_S2 = cs_S2[15];
end
always @ *
begin
    data_clk_en_S2 = !stall_real_S2 && cs_S2[18];
end
assign data_rdw_en_S2 = wr;
always @ *
begin
    if (msg_type_S2_f == 8'd12 || msg_type_S2_f == 8'd25)
    begin
        mshr_wr_state_en_S2 = n;
        mshr_state_in_S2 = 2'd0;
    end
    else if (msg_type_S2_f == 8'd23 
          || msg_type_S2_f == 8'd21
          || msg_type_S2_f == 8'd22)
    begin
        if (is_last_subline_S2)
        begin
             
            if (msg_type_S2_f == 8'd23 
            && ((l2_way_state_owner_S2 != 1) || smc_miss_S2_f || inv_fwd_pending_S2_f))
            
            
            begin
                mshr_wr_state_en_S2 = n;
                mshr_state_in_S2 = 2'd0;
            end
            else
            begin
                mshr_wr_state_en_S2 = !stall_S2;
                mshr_state_in_S2 = 2'd2;
            end
        end
        else
        begin
            mshr_wr_state_en_S2 = n;
            mshr_state_in_S2 = 2'd0;
        end
    end
    else
    begin
        mshr_wr_state_en_S2 = !stall_S2;
        mshr_state_in_S2 = 2'd2;
    end
end
always @ *
begin
    state_owner_en_S2 = !stall_S2 && cs_S2[14];
end
always @ *
begin
    state_owner_op_S2 = cs_S2[13:12];
end
always @ *
begin
    state_subline_en_S2 = !stall_S2 && cs_S2[11];
end
always @ *
begin
    state_subline_op_S2 = cs_S2[10:9];
end
always @ *
begin
    state_di_en_S2 = cs_S2[8];
end
always @ *
begin
    state_vd_en_S2 = !stall_S2 && cs_S2[7];
end
always @ *
begin
    state_vd_S2 = cs_S2[6:5];
end
always @ *
begin
    state_mesi_en_S2 = !stall_S2 && cs_S2[4];
end
always @ *
begin
    state_mesi_S2 = cs_S2[3:2];
end
always @ *
begin
    state_lru_en_S2 = !stall_S2 && cs_S2[1];
end
always @ *
begin
    state_lru_op_S2 = cs_S2[0];
end
always @ *
begin
    state_wr_en_S2 = !stall_S2 && (state_owner_en_S2 || state_subline_en_S2 || state_vd_en_S2
                  ||  state_di_en_S2 || state_mesi_en_S2 || state_lru_en_S2 || state_rb_en_S2);
end
always @ *
begin
    msg_data_ready_S2 = !stall_real_S2 && (data_clk_en_S2 || smc_wr_en_S2);
end
always @ *
begin
    smc_wr_en_S2 = valid_S2 && smc_miss_S2_f && (msg_type_S2_f == 8'd26);
end
assign state_rb_en_S2 = n;
always @ *
begin
    if (msg_type_S2_f == 8'd24)
    begin
        l2_load_64B_S2 = y;
        l2_load_32B_S2 = n;
    end
    else    
    begin
        l2_load_64B_S2 = n;
        l2_load_32B_S2 = n;
    end
end
reg [2-1:0] l2_load_data_subline_S2_f;
reg [2-1:0] l2_load_data_subline_S2_next;
always @ *
begin
    if (!rst_n)
    begin
        l2_load_data_subline_S2_next = 2'd0;
    end
    else if (valid_S2 && !stall_real_S2 && l2_load_64B_S2)
    begin
        l2_load_data_subline_S2_next = l2_load_data_subline_S2_f + 1;
    end
    else
    begin
        l2_load_data_subline_S2_next = l2_load_data_subline_S2_f;
    end
end
always @ (posedge clk)
begin
    l2_load_data_subline_S2_f <= l2_load_data_subline_S2_next;
end
always @ *
begin
    if (l2_load_64B_S2)
    begin
        stall_load_S2 = (l2_load_data_subline_S2_f != 2'd3);
    end
    else
    begin
        stall_load_S2 = n;
    end
end
always @ *
begin
    l2_load_data_subline_S2 = l2_load_data_subline_S2_f;
end
always @ *
begin
    stall_real_S2 = valid_S2 && ((cs_S2[18] || smc_wr_en_S2) && !msg_data_valid_S2);
end
always @ *
begin
    stall_S2 = valid_S2 && (stall_real_S2 || stall_load_S2);
end
always @ *
begin
    active_S2 = valid_S2;
end
reg valid_next_S2;
always @ *
begin
    valid_next_S2 = valid_S2 && !stall_S2;
end
reg valid_S3_f;
reg state_wr_en_S3_f;
reg mshr_wr_state_en_S3_f;
reg [2-1:0] mshr_state_in_S3_f;
reg smc_miss_S3_f;
reg msg_from_mshr_S3_f;
reg [8-1:0] msg_type_S3_f;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        valid_S3_f <= 1'b0;
        state_wr_en_S3_f <= 1'b0;
        mshr_wr_state_en_S3_f <= 0;
        mshr_state_in_S3_f <= 0;
        
        smc_miss_S3_f <= 0;
        
        msg_from_mshr_S3_f <= 0;
        msg_type_S3_f <= 0;
    end
    else if (!stall_S3)
    begin
        valid_S3_f <= valid_next_S2;
        state_wr_en_S3_f <= state_wr_en_S2;
        mshr_wr_state_en_S3_f <= mshr_wr_state_en_S2;
        mshr_state_in_S3_f <= mshr_state_in_S2;
        
        smc_miss_S3_f <= smc_miss_S2_f;
        
        msg_from_mshr_S3_f <= msg_from_mshr_S2_f;
        msg_type_S3_f <= msg_type_S2_f;
    end
end
always @ *
begin
    valid_S3 = valid_S3_f;
    state_wr_en_S3 = !stall_S3 && valid_S3 && state_wr_en_S3_f;
    mshr_wr_state_en_S3 = !stall_S3 && valid_S3 && mshr_wr_state_en_S3_f;
    mshr_state_in_S3 = mshr_state_in_S3_f;
    msg_type_S3 = msg_type_S3_f;
end
assign mshr_wr_data_en_S3 = 1'b0;
always @ *
begin
    mshr_inc_counter_en_S3 = valid_S3 && (msg_type_S3_f == 8'd23);
end
always @ *
begin
    active_S3 = valid_S3;
end
assign stall_S3 = 1'b0;
endmodule
      
 
module l2_pipe2_dpath(
    input wire clk,
    input wire rst_n,
    
    input wire [40-1:0] mshr_addr_S1,
    input wire [8-1:0] mshr_mshrid_S1,
    input wire [2-1:0] mshr_way_S1,
    input wire [14-1:0] mshr_src_chipid_S1,
    input wire [8-1:0] mshr_src_x_S1,
    input wire [8-1:0] mshr_src_y_S1,
    input wire [4-1:0] mshr_src_fbits_S1,
    input wire [10-1:0] mshr_sdid_S1,
    input wire [6-1:0] mshr_lsid_S1,
    input wire [6-1:0] mshr_miss_lsid_S1,
    input wire [40-1:0] msg_addr_S1,
    input wire [8-1:0] msg_type_S1,
    input wire [2-1:0] msg_subline_id_S1,
    input wire [8-1:0] msg_mshrid_S1,
    input wire [14-1:0] msg_src_chipid_S1,
    input wire [8-1:0] msg_src_x_S1,
    input wire [8-1:0] msg_src_y_S1,
    input wire [4-1:0] msg_src_fbits_S1,
    input wire [10-1:0] msg_sdid_S1,
    input wire [6-1:0] msg_lsid_S1,
    input wire valid_S1,
    input wire stall_S1,
    input wire msg_from_mshr_S1, 
    
    
    input wire [15*4+2+4-1:0] state_data_S2,
    input wire [104-1:0] tag_data_S2,
    input wire [128-1:0] msg_data_S2,
    input wire msg_from_mshr_S2,
    input wire [8-1:0] msg_type_S2,
   
    input wire [3-1:0] data_size_S2,
    input wire [1-1:0] cache_type_S2,
    input wire state_owner_en_S2,
    input wire [2-1:0] state_owner_op_S2,
    input wire state_subline_en_S2,
    input wire [2-1:0] state_subline_op_S2,
    input wire state_di_en_S2,
    input wire state_vd_en_S2,
    input wire [2-1:0] state_vd_S2,
    input wire state_mesi_en_S2,
    input wire [2-1:0] state_mesi_S2,
    input wire state_lru_en_S2,
    input wire [1-1:0] state_lru_op_S2,
    input wire state_rb_en_S2,
    input wire dir_clr_en_S2,
   
    input wire l2_load_64B_S2, 
    input wire l2_load_32B_S2, 
    input wire [2-1:0] l2_load_data_subline_S2,
 
    input wire valid_S2,
    input wire stall_S2,
    input wire stall_before_S2,
    
    input wire valid_S3,
    input wire stall_S3,
    
    
    
    output reg [40-1:0] addr_S1,
    output reg [3-1:0] mshr_rd_index_S1,
    output reg [8-1:0] tag_addr_S1,
    output reg [8-1:0] state_rd_addr_S1,
    
    output reg [104-1:0] tag_data_in_S1,
    output reg [104-1:0] tag_data_mask_in_S1,
    output reg is_same_address_S1,
    
   
 
    output reg [40-1:0] addr_S2,
    output reg l2_tag_hit_S2,
    output reg [2-1:0] l2_way_sel_S2,
    output reg l2_wb_S2,
    output reg [6-1:0] l2_way_state_owner_S2,
    output reg [2-1:0] l2_way_state_mesi_S2,
    output reg [2-1:0] l2_way_state_vd_S2,
    output reg [4-1:0] l2_way_state_subline_S2,
    output reg [1-1:0] l2_way_state_cache_type_S2,
    output reg addr_l2_aligned_S2,
    output reg subline_valid_S2, 
    output reg [6-1:0] lsid_S2,
    output reg [8+2-1:0] dir_addr_S2,
    output reg [64-1:0] dir_data_in_S2,
    output wire [64-1:0] dir_data_mask_in_S2,
    output reg [8+2+2-1:0] data_addr_S2,
    output reg [144-1:0] data_data_in_S2,
    output wire [144-1:0] data_data_mask_in_S2,
    
    output reg [16-1:0] smc_wr_addr_in_S2,
    output reg [128-1:0] smc_data_in_S2,
    
    
    output reg [40-1:0] addr_S3,
    output reg [3-1:0] mshr_wr_index_S3,
    output wire [120+2-1:0] mshr_data_in_S3,
    output wire [120+2-1:0] mshr_data_mask_in_S3,
    output reg [8-1:0] state_wr_addr_S3,
    output reg [15*4+2+4-1:0] state_data_in_S3,
    output reg [15*4+2+4-1:0] state_data_mask_in_S3
);
reg [8-1:0] mshrid_S1;
reg [14-1:0] src_chipid_S1;
reg [8-1:0] src_x_S1;
reg [8-1:0] src_y_S1;
reg [4-1:0] src_fbits_S1;
reg [10-1:0] sdid_S1;
reg [6-1:0] lsid_S1;
always @ *
begin
    if (msg_from_mshr_S1)
    begin
        addr_S1 = {mshr_addr_S1[39:6+8], mshr_addr_S1[6+8-1:6],
                         msg_subline_id_S1, mshr_addr_S1[3:0]};
 
        src_chipid_S1 = mshr_src_chipid_S1;
        src_x_S1 = mshr_src_x_S1;   
        src_y_S1 = mshr_src_y_S1;   
        src_fbits_S1 = mshr_src_fbits_S1;
        sdid_S1 = mshr_sdid_S1;
        lsid_S1 = mshr_lsid_S1;
    end
    else
    begin
        addr_S1 = msg_addr_S1;
        src_chipid_S1 = msg_src_chipid_S1;
        src_x_S1 = msg_src_x_S1;   
        src_y_S1 = msg_src_y_S1;   
        src_fbits_S1 = msg_src_fbits_S1;
        sdid_S1 = msg_sdid_S1;
        lsid_S1 = msg_lsid_S1;
    end
end
always @ *
begin
    is_same_address_S1 = (mshr_addr_S1 == msg_addr_S1);
end
always @ *
begin
    mshrid_S1 = msg_mshrid_S1;
end
always @ *
begin
    mshr_rd_index_S1 = msg_mshrid_S1;
end
always @ *
begin
    tag_addr_S1 = addr_S1[6+8-1:6];
end
always @ *
begin
    state_rd_addr_S1 = addr_S1[6+8-1:6];
end
always @ *
begin
    tag_data_in_S1 = {4{addr_S1[39:6+8]}};
end
always @ *
begin
    tag_data_mask_in_S1 = {{(4-1)*26{1'b0}},{26{1'b1}}} 
                       << (mshr_way_S1 * 26);
end
reg [40-1:0] addr_S2_f;
reg [8-1:0] mshrid_S2_f;
reg [14-1:0] src_chipid_S2_f;
reg [8-1:0] src_x_S2_f;
reg [8-1:0] src_y_S2_f;
reg [4-1:0] src_fbits_S2_f;
reg [10-1:0] sdid_S2_f;
reg [6-1:0] lsid_S2_f;
reg [2-1:0] mshr_way_S2_f;
reg [2-1:0] msg_subline_id_S2_f;
reg [6-1:0] mshr_miss_lsid_S2_f;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        addr_S2_f <= 0; 
        mshrid_S2_f <= 0;
        src_chipid_S2_f <= 0;
        src_x_S2_f <= 0;
        src_y_S2_f <= 0;
        src_fbits_S2_f <= 0;
        sdid_S2_f <= 0;
        lsid_S2_f <= 0;
        mshr_way_S2_f <= 0;
        msg_subline_id_S2_f <= 0;
        mshr_miss_lsid_S2_f <= 0;
    end
    else if (!stall_S2)
    begin
        addr_S2_f <= addr_S1;
        mshrid_S2_f <= mshrid_S1;
        src_chipid_S2_f <= src_chipid_S1;
        src_x_S2_f <= src_x_S1;
        src_y_S2_f <= src_y_S1;
        src_fbits_S2_f <= src_fbits_S1;
        sdid_S2_f <= sdid_S1;
        lsid_S2_f <= lsid_S1;
        mshr_way_S2_f <= mshr_way_S1;
        msg_subline_id_S2_f <= msg_subline_id_S1;
        mshr_miss_lsid_S2_f <= mshr_miss_lsid_S1;
    end
end
reg [15*4+2+4-1:0] state_data_in_S2;
reg [15*4+2+4-1:0] state_data_mask_in_S2;
always @ *
begin
    addr_S2 = addr_S2_f;
    lsid_S2 = lsid_S2_f;
end
reg [104-1:0] tag_data_buf_S2_f;
reg [104-1:0] tag_data_buf_S2_next;
reg [104-1:0] tag_data_trans_S2;
always @ *
begin
    if (!rst_n)
    begin
        tag_data_buf_S2_next = 0;
    end
    else if (stall_S2 && !stall_before_S2)
    begin
        tag_data_buf_S2_next = tag_data_S2;
    end
    else
    begin
        tag_data_buf_S2_next = tag_data_buf_S2_f;
    end
end
always @ (posedge clk)
begin
    tag_data_buf_S2_f <= tag_data_buf_S2_next;
end
always @ *
begin
    if (stall_before_S2)
    begin
        tag_data_trans_S2 = tag_data_buf_S2_f;
    end
    else
    begin
        tag_data_trans_S2 = tag_data_S2;
    end
end
reg [104-1:0] state_data_buf_S2_f;
reg [104-1:0] state_data_buf_S2_next;
reg [104-1:0] state_data_trans_S2;
always @ *
begin
    if (!rst_n)
    begin
        state_data_buf_S2_next = 0;
    end
    else if (stall_S2 && !stall_before_S2)
    begin
        state_data_buf_S2_next = state_data_S2;
    end
    else
    begin
        state_data_buf_S2_next = state_data_buf_S2_f;
    end
end
always @ (posedge clk)
begin
    state_data_buf_S2_f <= state_data_buf_S2_next;
end
always @ *
begin
    if (stall_before_S2)
    begin
        state_data_trans_S2 = state_data_buf_S2_f;
    end
    else
    begin
        state_data_trans_S2 = state_data_S2;
    end
end
reg [2-1:0] l2_hit_way_sel_S2;
reg [2-1:0] l2_rb_bits_S2;
reg [4-1:0] l2_lru_bits_S2;
always @ *
begin
    l2_rb_bits_S2 = state_data_trans_S2[15*4+2+4-1:15*4+4];
    l2_lru_bits_S2 = state_data_trans_S2[15*4+4-1:15*4];
end
reg [26 - 1:0] tag_data_way_S2 [3:0];
reg [3:0] tag_hit_way_S2;
reg [15 - 1:0] state_way_S2 [3:0];
always @ *
begin
    tag_data_way_S2[0] = tag_data_trans_S2[26 * 1 - 1: 26 * 0];
    tag_data_way_S2[1] = tag_data_trans_S2[26 * 2 - 1: 26 * 1];
    tag_data_way_S2[2] = tag_data_trans_S2[26 * 3 - 1: 26 * 2];
    tag_data_way_S2[3] = tag_data_trans_S2[26 * 4 - 1: 26 * 3];
end
always @ *
begin
    state_way_S2[0] = state_data_trans_S2[15 * 1 - 1: 
15 * 0];
    state_way_S2[1] = state_data_trans_S2[15 * 2 - 1: 
15 * 1];
    state_way_S2[2] = state_data_trans_S2[15 * 3 - 1: 
15 * 2];
    state_way_S2[3] = state_data_trans_S2[15 * 4 - 1: 
15 * 3];
end
always @ *
begin
    if ((addr_S2_f[39:6+8] == tag_data_way_S2[0]) && 
(state_way_S2[0][12:11] == 2'b10 || state_way_S2[0][12:11] == 2'b11 ))
    begin
        tag_hit_way_S2[0] = 1'b1;
    end
    else
    begin
        tag_hit_way_S2[0] = 1'b0;
    end
end
always @ *
begin
    if ((addr_S2_f[39:6+8] == tag_data_way_S2[1]) && 
(state_way_S2[1][12:11] == 2'b10 || state_way_S2[1][12:11] == 2'b11 ))
    begin
        tag_hit_way_S2[1] = 1'b1;
    end
    else
    begin
        tag_hit_way_S2[1] = 1'b0;
    end
end
always @ *
begin
    if ((addr_S2_f[39:6+8] == tag_data_way_S2[2]) && 
(state_way_S2[2][12:11] == 2'b10 || state_way_S2[2][12:11] == 2'b11 ))
    begin
        tag_hit_way_S2[2] = 1'b1;
    end
    else
    begin
        tag_hit_way_S2[2] = 1'b0;
    end
end
always @ *
begin
    if ((addr_S2_f[39:6+8] == tag_data_way_S2[3]) && 
(state_way_S2[3][12:11] == 2'b10 || state_way_S2[3][12:11] == 2'b11 ))
    begin
        tag_hit_way_S2[3] = 1'b1;
    end
    else
    begin
        tag_hit_way_S2[3] = 1'b0;
    end
end
always @ *
begin
    if (msg_from_mshr_S2)
    begin
        l2_tag_hit_S2 = tag_hit_way_S2[mshr_way_S2_f];
    end
    else
        l2_tag_hit_S2 = tag_hit_way_S2[0] || tag_hit_way_S2[1] || tag_hit_way_S2[2] || tag_hit_way_S2[3];
end
always @ *
begin
    l2_hit_way_sel_S2 = {2{1'bx}};
    if (tag_hit_way_S2[0])
    begin
        l2_hit_way_sel_S2 = 2'd0;
    end
    if (tag_hit_way_S2[1])
    begin
        l2_hit_way_sel_S2 = 2'd1;
    end
    if (tag_hit_way_S2[2])
    begin
        l2_hit_way_sel_S2 = 2'd2;
    end
    if (tag_hit_way_S2[3])
    begin
        l2_hit_way_sel_S2 = 2'd3;
    end
end
always @ *
begin
    if(valid_S2)
    begin
        if (msg_from_mshr_S2)
        begin
            l2_way_sel_S2 = mshr_way_S2_f;
        end
        else
        begin
            l2_way_sel_S2 = l2_hit_way_sel_S2;
        end
    end
    else
    begin
        l2_way_sel_S2 = 0;
    end
end
always @ *
begin
    if (!l2_tag_hit_S2 && (state_way_S2[l2_way_sel_S2][12:11] == 2'b11))
    begin
        l2_wb_S2 = 1'b1;
    end
    else
    begin
        l2_wb_S2 = 1'b0;
    end
end
always @ *
begin
    l2_way_state_mesi_S2 = state_way_S2[l2_way_sel_S2][14:13];
    l2_way_state_vd_S2 = state_way_S2[l2_way_sel_S2][12:11];
    l2_way_state_subline_S2 = state_way_S2[l2_way_sel_S2][9:6];
    l2_way_state_cache_type_S2 = state_way_S2[l2_way_sel_S2][10];
    l2_way_state_owner_S2 = state_way_S2[l2_way_sel_S2][5:0];
end
always @ *
begin
    dir_addr_S2 = {addr_S2_f[6+8-1:6],l2_way_sel_S2}; 
end
always @ *
begin
    if (l2_load_64B_S2)
    begin
        data_addr_S2 = {addr_S2_f[6+8-1:6],l2_way_sel_S2, l2_load_data_subline_S2};
    end
    else
    begin
        data_addr_S2 = {addr_S2_f[6+8-1:6],l2_way_sel_S2, addr_S2_f[5:4]};
    end
end
always @ *
begin
    addr_l2_aligned_S2 = (addr_S2_f[6-1:0] == {6{1'b0}}); 
end
assign dir_data_mask_in_S2 = {64{1'b1}};
always @ *
begin
    if (dir_clr_en_S2)
    begin
        dir_data_in_S2 = {(64){1'b0}}; 
    end
    else
    begin
        dir_data_in_S2 = {{(64-1){1'b0}},1'b1} << l2_way_state_owner_S2; 
    end
end
wire [8-1:0] msg_data_parity1_S2;
wire [8-1:0] msg_data_parity2_S2;
l2_data_pgen data_pgen1( 
    .din            (msg_data_S2[64-1:0]),
    .parity         (msg_data_parity1_S2)
);
l2_data_pgen data_pgen2( 
    .din            (msg_data_S2[128-1:64]),
    .parity         (msg_data_parity2_S2)
);
always @ *
begin
    data_data_in_S2 = {msg_data_parity2_S2, msg_data_S2[127:64], msg_data_parity1_S2, msg_data_S2[63:0]}; 
end
assign data_data_mask_in_S2 = {144{1'b1}}; 
reg [6-1:0] state_owner_S2;
reg [4-1:0] state_subline_S2;
reg [2-1:0] state_rb_S2;
reg [4-1:0] state_lru_S2;
always @ *
begin
    state_owner_S2 = l2_way_state_owner_S2; 
    if (state_owner_op_S2 == 2'd1)
    begin
        state_owner_S2 = sdid_S2_f[5:0]; 
    end
    else if (state_owner_op_S2 == 2'd2)
    begin
        state_owner_S2 = l2_way_state_owner_S2 + 1; 
    end
    else if (state_owner_op_S2 == 2'd3)
    begin
        state_owner_S2 = l2_way_state_owner_S2 - 1; 
    end
    else if (state_owner_op_S2 == 2'd0)
    begin
        state_owner_S2 = 0; 
    end
end
reg [4-1:0] addr_subline_S2;
always @ *
begin
    if (cache_type_S2 == 1'b0)
    begin
        
        addr_subline_S2= {{(4-1){1'b0}},1'b1} << addr_S2_f[5:4];
    end
    else
    begin
        
        addr_subline_S2= {{(4-2){1'b0}},2'b11} << (2*addr_S2_f[5]);
    end
end
always @ *
begin
    if (state_subline_op_S2 == 2'd1)
    begin
        state_subline_S2 = sdid_S2_f[9:6];
    end
    else if (state_subline_op_S2 == 2'd2)
    begin
        state_subline_S2 = l2_way_state_subline_S2 | addr_subline_S2;
    end
    else if (state_subline_op_S2 == 2'd3)
    begin
        state_subline_S2 = l2_way_state_subline_S2 & (~addr_subline_S2);
    end
    else if (state_subline_op_S2 == 2'd0)
    begin
        state_subline_S2 = {4{1'b0}};
    end
    else
    begin
        state_subline_S2 = {4{1'bx}};
    end
end
always @ *
begin
    state_rb_S2 = l2_rb_bits_S2 + 1; 
end
always @ *
begin
    if (state_lru_en_S2)
    begin
        if (state_lru_op_S2 == 1'b0)
        begin
            state_lru_S2 = l2_lru_bits_S2 & (~({{(4-1){1'b0}},1'b1} << l2_way_sel_S2));
        end
        else
        begin
            state_lru_S2 = l2_lru_bits_S2 | ({{(4-1){1'b0}},1'b1} << l2_way_sel_S2);
            if (state_lru_S2 == {4{1'b1}})
            begin
                state_lru_S2 = {4{1'b0}};
            end
        end
    end
    else
    begin
        state_lru_S2 = l2_lru_bits_S2; 
    end
end
always @ *
begin
    subline_valid_S2 = l2_way_state_subline_S2[msg_subline_id_S2_f]; 
end
always @ *
begin
    state_data_in_S2 = {state_rb_S2, state_lru_S2, 
    {4{state_mesi_S2, state_vd_S2, cache_type_S2, state_subline_S2, state_owner_S2}}};
end
reg [4*15-1:0] state_way_data_mask_in_S2;
always @ *
begin
    state_way_data_mask_in_S2 = {{(4-1)*15{1'b0}},
                                {{2{state_mesi_en_S2}}, 
                                 {2{state_vd_en_S2}}, 
                                 {1{state_di_en_S2}}, 
                                 {4{state_subline_en_S2}}, 
                                 {6{state_owner_en_S2}}}} 
    << (l2_way_sel_S2 * 15); 
end
always @ *
begin
    state_data_mask_in_S2 = {{2{state_rb_en_S2}}, 
                             {4{state_lru_en_S2}},
                              state_way_data_mask_in_S2}; 
end
always @ *
begin
    smc_wr_addr_in_S2 = {sdid_S2_f, mshr_miss_lsid_S2_f}; 
end
always @ *
begin
    smc_data_in_S2 = msg_data_S2; 
end
reg [40-1:0] addr_S3_f;
reg [15*4+2+4-1:0] state_data_in_S3_f;
reg [15*4+2+4-1:0] state_data_mask_in_S3_f;
reg [8-1:0] mshrid_S3_f;
reg [6-1:0] mshr_miss_lsid_S3_f;
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        addr_S3_f <= 0; 
        state_data_in_S3_f <= 0;
        state_data_mask_in_S3_f <= 0;
        mshrid_S3_f <= 0;
        mshr_miss_lsid_S3_f <= 0;
    end
    else if (!stall_S3)
    begin
        addr_S3_f <= addr_S2_f;
        state_data_in_S3_f <= state_data_in_S2;
        state_data_mask_in_S3_f <= state_data_mask_in_S2;
        mshrid_S3_f <= mshrid_S2_f;
        mshr_miss_lsid_S3_f <= mshr_miss_lsid_S2_f;
    end
end
always @ *
begin
    state_data_in_S3 = state_data_in_S3_f;
    state_data_mask_in_S3 = state_data_mask_in_S3_f;
    addr_S3 = addr_S3_f;
end
always @ *
begin
    state_wr_addr_S3 = addr_S3_f[6+8-1:6]; 
end
always @ *
begin
    mshr_wr_index_S3 = mshrid_S3_f; 
end
assign mshr_data_in_S3 = {120+2{1'b0}}; 
assign mshr_data_mask_in_S3 = {1'b1, {(120+2-1){1'b0}}}; 
endmodule
      
 
module l2_priority_encoder_1(
    input wire [1:0] data_in,
    output wire [0:0] data_out,
    output wire [1:0] data_out_mask,
    output wire nonzero_out
);
assign data_out = data_in[0] ? 1'b0 : 1'b1;
assign data_out_mask = data_in[0] ? 2'b10 : 2'b01;
assign nonzero_out = | (data_in[1:0]);
endmodule
module l2_priority_encoder_2(
    input wire [3:0] data_in,
    output wire [1:0] data_out,
    output wire [3:0] data_out_mask,
    output wire nonzero_out
);
wire [0:0] data_low;
wire [0:0] data_high;
wire [1:0] data_low_mask;
wire [1:0] data_high_mask;
wire nonzero_low;
wire nonzero_high;
l2_priority_encoder_1 encoder_high_1 (.data_in(data_in[3:2]), .data_out(data_high), .data_out_mask(data_high_mask), .nonzero_out(nonzero_high));
l2_priority_encoder_1 encoder_low_1(.data_in(data_in[1:0]), .data_out(data_low), .data_out_mask(data_low_mask), .nonzero_out(nonzero_low));
assign data_out = nonzero_low ? {1'b0, data_low} : {1'b1, data_high};
assign data_out_mask = nonzero_low ? {{2{1'b1}}, data_low_mask} : {data_high_mask,{2{1'b1}}};
assign nonzero_out = nonzero_low | nonzero_high;
endmodule
module l2_priority_encoder_3(
    input wire [7:0] data_in,
    output wire [2:0] data_out,
    output wire [7:0] data_out_mask,
    output wire nonzero_out
);
wire [1:0] data_low;
wire [1:0] data_high;
wire [3:0] data_low_mask;
wire [3:0] data_high_mask;
wire nonzero_low;
wire nonzero_high;
l2_priority_encoder_2 encoder_high_2 (.data_in(data_in[7:4]), .data_out(data_high), .data_out_mask(data_high_mask), .nonzero_out(nonzero_high));
l2_priority_encoder_2 encoder_low_2(.data_in(data_in[3:0]), .data_out(data_low), .data_out_mask(data_low_mask), .nonzero_out(nonzero_low));
assign data_out = nonzero_low ? {1'b0, data_low} : {1'b1, data_high};
assign data_out_mask = nonzero_low ? {{4{1'b1}}, data_low_mask} : {data_high_mask,{4{1'b1}}};
assign nonzero_out = nonzero_low | nonzero_high;
endmodule
module l2_priority_encoder_4(
    input wire [15:0] data_in,
    output wire [3:0] data_out,
    output wire [15:0] data_out_mask,
    output wire nonzero_out
);
wire [2:0] data_low;
wire [2:0] data_high;
wire [7:0] data_low_mask;
wire [7:0] data_high_mask;
wire nonzero_low;
wire nonzero_high;
l2_priority_encoder_3 encoder_high_3 (.data_in(data_in[15:8]), .data_out(data_high), .data_out_mask(data_high_mask), .nonzero_out(nonzero_high));
l2_priority_encoder_3 encoder_low_3(.data_in(data_in[7:0]), .data_out(data_low), .data_out_mask(data_low_mask), .nonzero_out(nonzero_low));
assign data_out = nonzero_low ? {1'b0, data_low} : {1'b1, data_high};
assign data_out_mask = nonzero_low ? {{8{1'b1}}, data_low_mask} : {data_high_mask,{8{1'b1}}};
assign nonzero_out = nonzero_low | nonzero_high;
endmodule
module l2_priority_encoder_5(
    input wire [31:0] data_in,
    output wire [4:0] data_out,
    output wire [31:0] data_out_mask,
    output wire nonzero_out
);
wire [3:0] data_low;
wire [3:0] data_high;
wire [15:0] data_low_mask;
wire [15:0] data_high_mask;
wire nonzero_low;
wire nonzero_high;
l2_priority_encoder_4 encoder_high_4 (.data_in(data_in[31:16]), .data_out(data_high), .data_out_mask(data_high_mask), .nonzero_out(nonzero_high));
l2_priority_encoder_4 encoder_low_4(.data_in(data_in[15:0]), .data_out(data_low), .data_out_mask(data_low_mask), .nonzero_out(nonzero_low));
assign data_out = nonzero_low ? {1'b0, data_low} : {1'b1, data_high};
assign data_out_mask = nonzero_low ? {{16{1'b1}}, data_low_mask} : {data_high_mask,{16{1'b1}}};
assign nonzero_out = nonzero_low | nonzero_high;
endmodule
module l2_priority_encoder_6(
    input wire [63:0] data_in,
    output wire [5:0] data_out,
    output wire [63:0] data_out_mask,
    output wire nonzero_out
);
wire [4:0] data_low;
wire [4:0] data_high;
wire [31:0] data_low_mask;
wire [31:0] data_high_mask;
wire nonzero_low;
wire nonzero_high;
l2_priority_encoder_5 encoder_high_5 (.data_in(data_in[63:32]), .data_out(data_high), .data_out_mask(data_high_mask), .nonzero_out(nonzero_high));
l2_priority_encoder_5 encoder_low_5(.data_in(data_in[31:0]), .data_out(data_low), .data_out_mask(data_low_mask), .nonzero_out(nonzero_low));
assign data_out = nonzero_low ? {1'b0, data_low} : {1'b1, data_high};
assign data_out_mask = nonzero_low ? {{32{1'b1}}, data_low_mask} : {data_high_mask,{32{1'b1}}};
assign nonzero_out = nonzero_low | nonzero_high;
endmodule
      
 
module l2_smc(
    input wire clk,
    input wire rst_n,
    
    input wire rd_en,
    
    input wire wr_en,
    
    input wire rd_diag_en,
    
    input wire wr_diag_en,
    
    input wire flush_en,
    input wire [2-1:0] addr_op,
    
    input wire [16-1:0] rd_addr_in,
    input wire [16-1:0] wr_addr_in,
    
    input wire [128-1:0] data_in,
    output reg hit,
    
    
    output reg [30-1:0] data_out,
    output reg [4-1:0] valid_out,
    output reg [14-1:0] tag_out
);
reg [16-1:0] entry_used_f;
reg [16-1:0] entry_used_next;
reg [16-1:0] entry_used_and_mask;
reg [16-1:0] entry_used_or_mask;
reg [16-1:0] entry_locked_f;
reg [16-1:0] entry_locked_next;
reg [16-1:0] entry_locked_and_mask;
reg [16-1:0] entry_locked_or_mask;
reg [138-1:0] data_mem_f [16-1:0];
reg [14-1:0] smc_tag [16-1:0];
reg [4-1:0] smc_valid [16-1:0];
reg [120-1:0] smc_data [16-1:0];
reg [10-1:0] smc_sdid [16-1:0];
reg [14-1:0] rd_tag_in;
reg [14-1:0] wr_tag_in;
reg [4-1:0] rd_index_in;
reg [4-1:0] wr_index_in;
reg [2-1:0] rd_offset_in;
reg [2-1:0] wr_offset_in;
reg [10-1:0] wr_sdid_in;
reg [4-1:0] smc_valid_in;
reg [120-1:0] smc_data_in;
reg [4-1:0] hit_index;
reg [4-1:0] replace_index;
reg wr_hit;
reg [4-1:0] wr_hit_index;
reg [4-1:0] wr_index;
always @ *
begin
    smc_tag[0] = data_mem_f[0][137:124];
    smc_tag[1] = data_mem_f[1][137:124];
    smc_tag[2] = data_mem_f[2][137:124];
    smc_tag[3] = data_mem_f[3][137:124];
    smc_tag[4] = data_mem_f[4][137:124];
    smc_tag[5] = data_mem_f[5][137:124];
    smc_tag[6] = data_mem_f[6][137:124];
    smc_tag[7] = data_mem_f[7][137:124];
    smc_tag[8] = data_mem_f[8][137:124];
    smc_tag[9] = data_mem_f[9][137:124];
    smc_tag[10] = data_mem_f[10][137:124];
    smc_tag[11] = data_mem_f[11][137:124];
    smc_tag[12] = data_mem_f[12][137:124];
    smc_tag[13] = data_mem_f[13][137:124];
    smc_tag[14] = data_mem_f[14][137:124];
    smc_tag[15] = data_mem_f[15][137:124];
end
always @ *
begin
    smc_valid[0] = data_mem_f[0][123:120];
    smc_valid[1] = data_mem_f[1][123:120];
    smc_valid[2] = data_mem_f[2][123:120];
    smc_valid[3] = data_mem_f[3][123:120];
    smc_valid[4] = data_mem_f[4][123:120];
    smc_valid[5] = data_mem_f[5][123:120];
    smc_valid[6] = data_mem_f[6][123:120];
    smc_valid[7] = data_mem_f[7][123:120];
    smc_valid[8] = data_mem_f[8][123:120];
    smc_valid[9] = data_mem_f[9][123:120];
    smc_valid[10] = data_mem_f[10][123:120];
    smc_valid[11] = data_mem_f[11][123:120];
    smc_valid[12] = data_mem_f[12][123:120];
    smc_valid[13] = data_mem_f[13][123:120];
    smc_valid[14] = data_mem_f[14][123:120];
    smc_valid[15] = data_mem_f[15][123:120];
end
always @ *
begin
    smc_data[0] = data_mem_f[0][119:0];
    smc_data[1] = data_mem_f[1][119:0];
    smc_data[2] = data_mem_f[2][119:0];
    smc_data[3] = data_mem_f[3][119:0];
    smc_data[4] = data_mem_f[4][119:0];
    smc_data[5] = data_mem_f[5][119:0];
    smc_data[6] = data_mem_f[6][119:0];
    smc_data[7] = data_mem_f[7][119:0];
    smc_data[8] = data_mem_f[8][119:0];
    smc_data[9] = data_mem_f[9][119:0];
    smc_data[10] = data_mem_f[10][119:0];
    smc_data[11] = data_mem_f[11][119:0];
    smc_data[12] = data_mem_f[12][119:0];
    smc_data[13] = data_mem_f[13][119:0];
    smc_data[14] = data_mem_f[14][119:0];
    smc_data[15] = data_mem_f[15][119:0];
end
always @ *
begin
    smc_sdid[0] = data_mem_f[0][137:128];
    smc_sdid[1] = data_mem_f[1][137:128];
    smc_sdid[2] = data_mem_f[2][137:128];
    smc_sdid[3] = data_mem_f[3][137:128];
    smc_sdid[4] = data_mem_f[4][137:128];
    smc_sdid[5] = data_mem_f[5][137:128];
    smc_sdid[6] = data_mem_f[6][137:128];
    smc_sdid[7] = data_mem_f[7][137:128];
    smc_sdid[8] = data_mem_f[8][137:128];
    smc_sdid[9] = data_mem_f[9][137:128];
    smc_sdid[10] = data_mem_f[10][137:128];
    smc_sdid[11] = data_mem_f[11][137:128];
    smc_sdid[12] = data_mem_f[12][137:128];
    smc_sdid[13] = data_mem_f[13][137:128];
    smc_sdid[14] = data_mem_f[14][137:128];
    smc_sdid[15] = data_mem_f[15][137:128];
end
always @ *
begin
    rd_tag_in = rd_addr_in[15:2];
    rd_offset_in = rd_addr_in[1:0];
    rd_index_in = rd_addr_in[5:2];
end
always @ *
begin
    wr_tag_in = wr_addr_in[15:2];
    wr_offset_in = wr_addr_in[1:0];
    wr_index_in = wr_addr_in[5:2];
    wr_sdid_in = wr_addr_in[15:6];
end
always @ *
begin
    smc_valid_in = { data_in[127], data_in[95], data_in[63], data_in[31] };
    smc_data_in = { data_in[125:96], data_in[93:64], data_in[61:32], data_in[29:0] };
end
wire [4-1:0] tag_hit_index;
wire tag_hit;
reg [15:0] smc_tag_cmp;
always @ *
begin
    smc_tag_cmp[0] = (smc_tag[0] == rd_tag_in) && smc_valid[0][rd_offset_in];
    smc_tag_cmp[1] = (smc_tag[1] == rd_tag_in) && smc_valid[1][rd_offset_in];
    smc_tag_cmp[2] = (smc_tag[2] == rd_tag_in) && smc_valid[2][rd_offset_in];
    smc_tag_cmp[3] = (smc_tag[3] == rd_tag_in) && smc_valid[3][rd_offset_in];
    smc_tag_cmp[4] = (smc_tag[4] == rd_tag_in) && smc_valid[4][rd_offset_in];
    smc_tag_cmp[5] = (smc_tag[5] == rd_tag_in) && smc_valid[5][rd_offset_in];
    smc_tag_cmp[6] = (smc_tag[6] == rd_tag_in) && smc_valid[6][rd_offset_in];
    smc_tag_cmp[7] = (smc_tag[7] == rd_tag_in) && smc_valid[7][rd_offset_in];
    smc_tag_cmp[8] = (smc_tag[8] == rd_tag_in) && smc_valid[8][rd_offset_in];
    smc_tag_cmp[9] = (smc_tag[9] == rd_tag_in) && smc_valid[9][rd_offset_in];
    smc_tag_cmp[10] = (smc_tag[10] == rd_tag_in) && smc_valid[10][rd_offset_in];
    smc_tag_cmp[11] = (smc_tag[11] == rd_tag_in) && smc_valid[11][rd_offset_in];
    smc_tag_cmp[12] = (smc_tag[12] == rd_tag_in) && smc_valid[12][rd_offset_in];
    smc_tag_cmp[13] = (smc_tag[13] == rd_tag_in) && smc_valid[13][rd_offset_in];
    smc_tag_cmp[14] = (smc_tag[14] == rd_tag_in) && smc_valid[14][rd_offset_in];
    smc_tag_cmp[15] = (smc_tag[15] == rd_tag_in) && smc_valid[15][rd_offset_in];
end
l2_priority_encoder_4 priority_encoder_cmp_4bits( 
    .data_in        (smc_tag_cmp),
    .data_out       (tag_hit_index),
    .data_out_mask  (),
    .nonzero_out    (tag_hit)
);
always @ *
begin
    if (rd_en && rd_diag_en)
    begin
        hit = 1'b0;
        hit_index = rd_index_in;
    end
    else
    begin
        if(rd_en)
        begin
            hit = tag_hit;
            hit_index = tag_hit_index;
        end
        else
        begin
            hit = 1'b0;
            hit_index = 0;
        end
    end
end
wire [4-1:0] tag_wr_hit_index;
wire tag_wr_hit;
reg [15:0] smc_tag_wr_cmp;
always @ *
begin
    smc_tag_wr_cmp[0] = (smc_tag[0] == wr_tag_in) && (smc_valid[0] != 0);
    smc_tag_wr_cmp[1] = (smc_tag[1] == wr_tag_in) && (smc_valid[1] != 0);
    smc_tag_wr_cmp[2] = (smc_tag[2] == wr_tag_in) && (smc_valid[2] != 0);
    smc_tag_wr_cmp[3] = (smc_tag[3] == wr_tag_in) && (smc_valid[3] != 0);
    smc_tag_wr_cmp[4] = (smc_tag[4] == wr_tag_in) && (smc_valid[4] != 0);
    smc_tag_wr_cmp[5] = (smc_tag[5] == wr_tag_in) && (smc_valid[5] != 0);
    smc_tag_wr_cmp[6] = (smc_tag[6] == wr_tag_in) && (smc_valid[6] != 0);
    smc_tag_wr_cmp[7] = (smc_tag[7] == wr_tag_in) && (smc_valid[7] != 0);
    smc_tag_wr_cmp[8] = (smc_tag[8] == wr_tag_in) && (smc_valid[8] != 0);
    smc_tag_wr_cmp[9] = (smc_tag[9] == wr_tag_in) && (smc_valid[9] != 0);
    smc_tag_wr_cmp[10] = (smc_tag[10] == wr_tag_in) && (smc_valid[10] != 0);
    smc_tag_wr_cmp[11] = (smc_tag[11] == wr_tag_in) && (smc_valid[11] != 0);
    smc_tag_wr_cmp[12] = (smc_tag[12] == wr_tag_in) && (smc_valid[12] != 0);
    smc_tag_wr_cmp[13] = (smc_tag[13] == wr_tag_in) && (smc_valid[13] != 0);
    smc_tag_wr_cmp[14] = (smc_tag[14] == wr_tag_in) && (smc_valid[14] != 0);
    smc_tag_wr_cmp[15] = (smc_tag[15] == wr_tag_in) && (smc_valid[15] != 0);
end
l2_priority_encoder_4 priority_encoder_wr_cmp_4bits( 
    .data_in        (smc_tag_wr_cmp),
    .data_out       (tag_wr_hit_index),
    .data_out_mask  (),
    .nonzero_out    (tag_wr_hit)
);
always @ *
begin
    if(wr_en || (flush_en && (addr_op == 2'd1)))
    begin
        wr_hit = tag_wr_hit;
        wr_hit_index = tag_wr_hit_index;
    end
    else
    begin
        wr_hit = 1'b0;
        wr_hit_index = 0;
    end
end
always @ *
begin
    data_out = smc_data[hit_index]>>(rd_offset_in * 30);
    valid_out = smc_valid[hit_index];
    tag_out = smc_tag[hit_index];
end
always @ *
begin
    entry_locked_and_mask = {16{1'b1}};
    entry_locked_or_mask = {16{1'b0}};
    if (!rst_n)
    begin
        entry_locked_and_mask = {16{1'b0}};
    end
    else if (wr_en && ~wr_diag_en)
    begin
        if(smc_valid_in)
        begin
            entry_locked_or_mask[wr_index] = 1'b1;
        end
        else
        begin
            entry_locked_and_mask[wr_index] = 1'b0;
        end
        if (rd_en && ~rd_diag_en && hit && (wr_index != hit_index) && entry_locked_f[hit_index])
        begin
            entry_locked_and_mask[hit_index] = 1'b0;
        end 
    end
    else if (rd_en && ~rd_diag_en && hit && entry_locked_f[hit_index])
    begin
        entry_locked_and_mask[hit_index] = 1'b0;
    end
end
always @ *
begin
    entry_locked_next = (entry_locked_f & entry_locked_and_mask) | entry_locked_or_mask;
end
always @ (posedge clk)
begin
    entry_locked_f <= entry_locked_next;
end
always @ *
begin
    entry_used_and_mask = {16{1'b1}};
    entry_used_or_mask = {16{1'b0}};
    if (!rst_n)
    begin
        entry_used_and_mask = {16{1'b0}};
    end
    else if (wr_en && ~wr_diag_en)
    begin
        if(smc_valid_in)
        begin
            entry_used_or_mask[wr_index] = 1'b1;
        end
        else
        begin
            entry_used_and_mask[wr_index] = 1'b0;
        end
        if (rd_en && ~rd_diag_en && hit && (wr_index != hit_index))
        begin
            entry_used_or_mask[hit_index] = 1'b1;
        end 
    end
    else if (rd_en && ~rd_diag_en && hit)
    begin
        entry_used_or_mask[hit_index] = 1'b1;
    end
end
always @ *
begin
    entry_used_next = (entry_used_f & entry_used_and_mask) | entry_used_or_mask;
    if (entry_used_next == {16{1'b1}})
    begin
        entry_used_next = {16{1'b0}};
    end
end
always @ (posedge clk)
begin
    entry_used_f <= entry_used_next;
end
wire [4-1:0] entry_replace_index;
wire replace_hit;
reg [15:0] replace_cmp;
always @ *
begin
    replace_cmp[0] = (~entry_used_f[0] && ~entry_locked_f[0]);
    replace_cmp[1] = (~entry_used_f[1] && ~entry_locked_f[1]);
    replace_cmp[2] = (~entry_used_f[2] && ~entry_locked_f[2]);
    replace_cmp[3] = (~entry_used_f[3] && ~entry_locked_f[3]);
    replace_cmp[4] = (~entry_used_f[4] && ~entry_locked_f[4]);
    replace_cmp[5] = (~entry_used_f[5] && ~entry_locked_f[5]);
    replace_cmp[6] = (~entry_used_f[6] && ~entry_locked_f[6]);
    replace_cmp[7] = (~entry_used_f[7] && ~entry_locked_f[7]);
    replace_cmp[8] = (~entry_used_f[8] && ~entry_locked_f[8]);
    replace_cmp[9] = (~entry_used_f[9] && ~entry_locked_f[9]);
    replace_cmp[10] = (~entry_used_f[10] && ~entry_locked_f[10]);
    replace_cmp[11] = (~entry_used_f[11] && ~entry_locked_f[11]);
    replace_cmp[12] = (~entry_used_f[12] && ~entry_locked_f[12]);
    replace_cmp[13] = (~entry_used_f[13] && ~entry_locked_f[13]);
    replace_cmp[14] = (~entry_used_f[14] && ~entry_locked_f[14]);
    replace_cmp[15] = (~entry_used_f[15] && ~entry_locked_f[15]);
end
l2_priority_encoder_4 priority_encoder_replace_cmp_4bits( 
    .data_in        (replace_cmp),
    .data_out       (entry_replace_index),
    .data_out_mask  (),
    .nonzero_out    (replace_hit)
);
always @ *
begin
    if (replace_hit)
    begin
        replace_index = entry_replace_index;
    end
    else
    begin
        replace_index = {4{1'b0}};
    end
end
always @ *
begin
    if (wr_en && wr_diag_en)
    begin
        wr_index = wr_index_in;
    end
    else if ((flush_en || wr_en) && wr_hit)
    begin
        wr_index = wr_hit_index;
    end
    else
    begin
        wr_index = replace_index;
    end
end
always @ (posedge clk)
begin
    if (!rst_n)
    begin
        data_mem_f[0] <= {138{1'b0}};
        data_mem_f[1] <= {138{1'b0}};
        data_mem_f[2] <= {138{1'b0}};
        data_mem_f[3] <= {138{1'b0}};
        data_mem_f[4] <= {138{1'b0}};
        data_mem_f[5] <= {138{1'b0}};
        data_mem_f[6] <= {138{1'b0}};
        data_mem_f[7] <= {138{1'b0}};
        data_mem_f[8] <= {138{1'b0}};
        data_mem_f[9] <= {138{1'b0}};
        data_mem_f[10] <= {138{1'b0}};
        data_mem_f[11] <= {138{1'b0}};
        data_mem_f[12] <= {138{1'b0}};
        data_mem_f[13] <= {138{1'b0}};
        data_mem_f[14] <= {138{1'b0}};
        data_mem_f[15] <= {138{1'b0}};
    end
    else if (flush_en)
    begin
        case (addr_op)
        2'd0:
        begin
            data_mem_f[0][123:120] <= {4{1'b0}};
            data_mem_f[1][123:120] <= {4{1'b0}};
            data_mem_f[2][123:120] <= {4{1'b0}};
            data_mem_f[3][123:120] <= {4{1'b0}};
            data_mem_f[4][123:120] <= {4{1'b0}};
            data_mem_f[5][123:120] <= {4{1'b0}};
            data_mem_f[6][123:120] <= {4{1'b0}};
            data_mem_f[7][123:120] <= {4{1'b0}};
            data_mem_f[8][123:120] <= {4{1'b0}};
            data_mem_f[9][123:120] <= {4{1'b0}};
            data_mem_f[10][123:120] <= {4{1'b0}};
            data_mem_f[11][123:120] <= {4{1'b0}};
            data_mem_f[12][123:120] <= {4{1'b0}};
            data_mem_f[13][123:120] <= {4{1'b0}};
            data_mem_f[14][123:120] <= {4{1'b0}};
            data_mem_f[15][123:120] <= {4{1'b0}};
        end
        2'd1:
        begin
            if (wr_hit)
            begin
                data_mem_f[wr_index][120+wr_offset_in] <= 1'b0;
                
            end
        end
        2'd2:
        begin
            if ((smc_sdid[0] == wr_sdid_in) && (smc_valid[0] != 0))
                data_mem_f[0][123:120] <= {4{1'b0}};
            if ((smc_sdid[1] == wr_sdid_in) && (smc_valid[1] != 0))
                data_mem_f[1][123:120] <= {4{1'b0}};
            if ((smc_sdid[2] == wr_sdid_in) && (smc_valid[2] != 0))
                data_mem_f[2][123:120] <= {4{1'b0}};
            if ((smc_sdid[3] == wr_sdid_in) && (smc_valid[3] != 0))
                data_mem_f[3][123:120] <= {4{1'b0}};
            if ((smc_sdid[4] == wr_sdid_in) && (smc_valid[4] != 0))
                data_mem_f[4][123:120] <= {4{1'b0}};
            if ((smc_sdid[5] == wr_sdid_in) && (smc_valid[5] != 0))
                data_mem_f[5][123:120] <= {4{1'b0}};
            if ((smc_sdid[6] == wr_sdid_in) && (smc_valid[6] != 0))
                data_mem_f[6][123:120] <= {4{1'b0}};
            if ((smc_sdid[7] == wr_sdid_in) && (smc_valid[7] != 0))
                data_mem_f[7][123:120] <= {4{1'b0}};
            if ((smc_sdid[8] == wr_sdid_in) && (smc_valid[8] != 0))
                data_mem_f[8][123:120] <= {4{1'b0}};
            if ((smc_sdid[9] == wr_sdid_in) && (smc_valid[9] != 0))
                data_mem_f[9][123:120] <= {4{1'b0}};
            if ((smc_sdid[10] == wr_sdid_in) && (smc_valid[10] != 0))
                data_mem_f[10][123:120] <= {4{1'b0}};
            if ((smc_sdid[11] == wr_sdid_in) && (smc_valid[11] != 0))
                data_mem_f[11][123:120] <= {4{1'b0}};
            if ((smc_sdid[12] == wr_sdid_in) && (smc_valid[12] != 0))
                data_mem_f[12][123:120] <= {4{1'b0}};
            if ((smc_sdid[13] == wr_sdid_in) && (smc_valid[13] != 0))
                data_mem_f[13][123:120] <= {4{1'b0}};
            if ((smc_sdid[14] == wr_sdid_in) && (smc_valid[14] != 0))
                data_mem_f[14][123:120] <= {4{1'b0}};
            if ((smc_sdid[15] == wr_sdid_in) && (smc_valid[15] != 0))
                data_mem_f[15][123:120] <= {4{1'b0}};
        end
        default:
        begin
            data_mem_f[wr_index] <= data_mem_f[wr_index];
        end
        endcase
    end
    else if (wr_en)
    begin
        if (wr_diag_en)
        begin
            case (addr_op)
            2'd0:
            begin
                case (wr_offset_in)
                2'd0:
                begin
                    data_mem_f[wr_index][30-1:0] <= 
                    data_in[30-1:0];
                end
                2'd1:
                begin
                    data_mem_f[wr_index][30*2-1:30] <= 
                    data_in[30-1:0];
                end
                2'd2:
                begin
                    data_mem_f[wr_index][30*3-1:30*2] <= 
                    data_in[30-1:0];
                end
                2'd3:
                begin
                    data_mem_f[wr_index][30*4-1:30*3] <= 
                    data_in[30-1:0];
                end
                default:
                begin
                    data_mem_f[wr_index] <= data_mem_f[wr_index];
                end
                endcase
            end
            2'd1:
            begin
                data_mem_f[wr_index][123:120] <= data_in[4-1:0];
            end
            2'd2: 
            begin
                data_mem_f[wr_index][137:124] <= data_in[14-1:0];
            end
            default:
            begin
                data_mem_f[wr_index] <= data_mem_f[wr_index];
            end
            endcase
        end
        else
        begin
            data_mem_f[wr_index] <= {wr_tag_in, smc_valid_in, smc_data_in};
        end
    end
end
endmodule
      
 
module l2_state(
    input wire clk,
    input wire rst_n,
    input wire pdout_en,
    input wire deepsleep,
    input wire rd_en,
    input wire wr_en,
    input wire [8-1:0] rd_addr,
    input wire [8-1:0] wr_addr,
    input wire [15*4+2+4-1:0] data_in,
    input wire [15*4+2+4-1:0] data_mask_in,
    output reg [15*4+2+4-1:0] data_out,
    output wire [15*4+2+4-1:0] pdata_out,
    
    output wire [4-1:0] srams_rtap_data,
    input wire  [4-1:0] rtap_srams_bist_command,
    input wire  [4-1:0] rtap_srams_bist_data
);
reg [15*4+2+4-1:0] data_in_buf;
reg [15*4+2+4-1:0] data_mask_in_buf;
wire [15*4+2+4-1:0] data_out_real;
always @ (posedge clk)
begin
    data_in_buf <= data_in;
    data_mask_in_buf <= data_mask_in;
end
reg bypass_f;
reg bypass_next;
always @ *
begin
    if (rd_en && wr_en && (rd_addr == wr_addr))
    begin
        bypass_next = 1'b1;
    end
    else
    begin
        bypass_next = 1'b0;
    end
end
always @ (posedge clk)
begin
    bypass_f <= bypass_next;
end
always @ *
begin
    if (bypass_f)
    begin
        data_out[0] = data_mask_in_buf[0] ? data_in_buf[0] : data_out_real[0];
    
        data_out[1] = data_mask_in_buf[1] ? data_in_buf[1] : data_out_real[1];
    
        data_out[2] = data_mask_in_buf[2] ? data_in_buf[2] : data_out_real[2];
    
        data_out[3] = data_mask_in_buf[3] ? data_in_buf[3] : data_out_real[3];
    
        data_out[4] = data_mask_in_buf[4] ? data_in_buf[4] : data_out_real[4];
    
        data_out[5] = data_mask_in_buf[5] ? data_in_buf[5] : data_out_real[5];
    
        data_out[6] = data_mask_in_buf[6] ? data_in_buf[6] : data_out_real[6];
    
        data_out[7] = data_mask_in_buf[7] ? data_in_buf[7] : data_out_real[7];
    
        data_out[8] = data_mask_in_buf[8] ? data_in_buf[8] : data_out_real[8];
    
        data_out[9] = data_mask_in_buf[9] ? data_in_buf[9] : data_out_real[9];
    
        data_out[10] = data_mask_in_buf[10] ? data_in_buf[10] : data_out_real[10];
    
        data_out[11] = data_mask_in_buf[11] ? data_in_buf[11] : data_out_real[11];
    
        data_out[12] = data_mask_in_buf[12] ? data_in_buf[12] : data_out_real[12];
    
        data_out[13] = data_mask_in_buf[13] ? data_in_buf[13] : data_out_real[13];
    
        data_out[14] = data_mask_in_buf[14] ? data_in_buf[14] : data_out_real[14];
    
        data_out[15] = data_mask_in_buf[15] ? data_in_buf[15] : data_out_real[15];
    
        data_out[16] = data_mask_in_buf[16] ? data_in_buf[16] : data_out_real[16];
    
        data_out[17] = data_mask_in_buf[17] ? data_in_buf[17] : data_out_real[17];
    
        data_out[18] = data_mask_in_buf[18] ? data_in_buf[18] : data_out_real[18];
    
        data_out[19] = data_mask_in_buf[19] ? data_in_buf[19] : data_out_real[19];
    
        data_out[20] = data_mask_in_buf[20] ? data_in_buf[20] : data_out_real[20];
    
        data_out[21] = data_mask_in_buf[21] ? data_in_buf[21] : data_out_real[21];
    
        data_out[22] = data_mask_in_buf[22] ? data_in_buf[22] : data_out_real[22];
    
        data_out[23] = data_mask_in_buf[23] ? data_in_buf[23] : data_out_real[23];
    
        data_out[24] = data_mask_in_buf[24] ? data_in_buf[24] : data_out_real[24];
    
        data_out[25] = data_mask_in_buf[25] ? data_in_buf[25] : data_out_real[25];
    
        data_out[26] = data_mask_in_buf[26] ? data_in_buf[26] : data_out_real[26];
    
        data_out[27] = data_mask_in_buf[27] ? data_in_buf[27] : data_out_real[27];
    
        data_out[28] = data_mask_in_buf[28] ? data_in_buf[28] : data_out_real[28];
    
        data_out[29] = data_mask_in_buf[29] ? data_in_buf[29] : data_out_real[29];
    
        data_out[30] = data_mask_in_buf[30] ? data_in_buf[30] : data_out_real[30];
    
        data_out[31] = data_mask_in_buf[31] ? data_in_buf[31] : data_out_real[31];
    
        data_out[32] = data_mask_in_buf[32] ? data_in_buf[32] : data_out_real[32];
    
        data_out[33] = data_mask_in_buf[33] ? data_in_buf[33] : data_out_real[33];
    
        data_out[34] = data_mask_in_buf[34] ? data_in_buf[34] : data_out_real[34];
    
        data_out[35] = data_mask_in_buf[35] ? data_in_buf[35] : data_out_real[35];
    
        data_out[36] = data_mask_in_buf[36] ? data_in_buf[36] : data_out_real[36];
    
        data_out[37] = data_mask_in_buf[37] ? data_in_buf[37] : data_out_real[37];
    
        data_out[38] = data_mask_in_buf[38] ? data_in_buf[38] : data_out_real[38];
    
        data_out[39] = data_mask_in_buf[39] ? data_in_buf[39] : data_out_real[39];
    
        data_out[40] = data_mask_in_buf[40] ? data_in_buf[40] : data_out_real[40];
    
        data_out[41] = data_mask_in_buf[41] ? data_in_buf[41] : data_out_real[41];
    
        data_out[42] = data_mask_in_buf[42] ? data_in_buf[42] : data_out_real[42];
    
        data_out[43] = data_mask_in_buf[43] ? data_in_buf[43] : data_out_real[43];
    
        data_out[44] = data_mask_in_buf[44] ? data_in_buf[44] : data_out_real[44];
    
        data_out[45] = data_mask_in_buf[45] ? data_in_buf[45] : data_out_real[45];
    
        data_out[46] = data_mask_in_buf[46] ? data_in_buf[46] : data_out_real[46];
    
        data_out[47] = data_mask_in_buf[47] ? data_in_buf[47] : data_out_real[47];
    
        data_out[48] = data_mask_in_buf[48] ? data_in_buf[48] : data_out_real[48];
    
        data_out[49] = data_mask_in_buf[49] ? data_in_buf[49] : data_out_real[49];
    
        data_out[50] = data_mask_in_buf[50] ? data_in_buf[50] : data_out_real[50];
    
        data_out[51] = data_mask_in_buf[51] ? data_in_buf[51] : data_out_real[51];
    
        data_out[52] = data_mask_in_buf[52] ? data_in_buf[52] : data_out_real[52];
    
        data_out[53] = data_mask_in_buf[53] ? data_in_buf[53] : data_out_real[53];
    
        data_out[54] = data_mask_in_buf[54] ? data_in_buf[54] : data_out_real[54];
    
        data_out[55] = data_mask_in_buf[55] ? data_in_buf[55] : data_out_real[55];
    
        data_out[56] = data_mask_in_buf[56] ? data_in_buf[56] : data_out_real[56];
    
        data_out[57] = data_mask_in_buf[57] ? data_in_buf[57] : data_out_real[57];
    
        data_out[58] = data_mask_in_buf[58] ? data_in_buf[58] : data_out_real[58];
    
        data_out[59] = data_mask_in_buf[59] ? data_in_buf[59] : data_out_real[59];
    
        data_out[60] = data_mask_in_buf[60] ? data_in_buf[60] : data_out_real[60];
    
        data_out[61] = data_mask_in_buf[61] ? data_in_buf[61] : data_out_real[61];
    
        data_out[62] = data_mask_in_buf[62] ? data_in_buf[62] : data_out_real[62];
    
        data_out[63] = data_mask_in_buf[63] ? data_in_buf[63] : data_out_real[63];
    
        data_out[64] = data_mask_in_buf[64] ? data_in_buf[64] : data_out_real[64];
    
        data_out[65] = data_mask_in_buf[65] ? data_in_buf[65] : data_out_real[65];
    
    end
    else
    begin
        data_out = data_out_real;
    end
end
 
 sram_l2_state l2_state_array (
     .RESET_N(rst_n),
     .MEMCLK         (clk),
     .CEA            (rd_en),
     .RDWENA          (1'b1),
     .AA             (rd_addr),
     .BWA             (),
     .DINA            (),
     .DOUTA           (data_out_real),
     .CEB            (wr_en),
     .RDWENB            (1'b0),
     .AB             (wr_addr),
     .BWB             (data_mask_in),
     .DINB            (data_in),
     .DOUTB           (),
    .BIST_COMMAND(rtap_srams_bist_command),
    .BIST_DIN(rtap_srams_bist_data),
    .BIST_DOUT(srams_rtap_data),
    .SRAMID(8'd15)
 );
endmodule
module cpx_arbitrator(
   clk,
   rst_n,
   uncore_spc_data_ready,
   uncore_spc_data,
   uncore_spc_grant,
   rtap_arb_req_val,
   rtap_arb_req_data,
   rtap_arb_req_threadid,
   fpu_arb_data_rdy,
   fpu_arb_data,
   fpu_arb_grant,
   cpx_arb_spc_data_rdy,
   cpx_arb_spc_data,
   cpx_arb_spc_grant
   );
   input clk;
   input rst_n;
   input               uncore_spc_data_ready;
   input [144:0]       uncore_spc_data;
   input [4:0]         uncore_spc_grant;
   input               fpu_arb_data_rdy;
   input [144:0]       fpu_arb_data;
   input               fpu_arb_grant;
   input               rtap_arb_req_val;
   input [63:0]        rtap_arb_req_data;
   input [1:0]         rtap_arb_req_threadid;
   output reg          cpx_arb_spc_data_rdy;
   output reg [144:0]  cpx_arb_spc_data;
   output reg [4:0]    cpx_arb_spc_grant;
   reg [144:0]         rtap_interrupt_packet;
   always @ *
   begin
      
      rtap_interrupt_packet = 0;
      rtap_interrupt_packet[144] = 1'b1;
      rtap_interrupt_packet[143:140] = 4'b0111;
      rtap_interrupt_packet[135:134] = rtap_arb_req_threadid;
      rtap_interrupt_packet[63:0] = rtap_arb_req_data;
   end
   always @*
   begin
      cpx_arb_spc_data_rdy = uncore_spc_data_ready | fpu_arb_data_rdy | rtap_arb_req_val;
      
      cpx_arb_spc_data = 0;
      if (uncore_spc_data_ready)
         cpx_arb_spc_data = uncore_spc_data;
      else if (fpu_arb_data_rdy)
         cpx_arb_spc_data = fpu_arb_data;
      else if (rtap_arb_req_val)
         cpx_arb_spc_data = rtap_interrupt_packet;
      cpx_arb_spc_grant[4:1] = uncore_spc_grant;
      cpx_arb_spc_grant[0] = fpu_arb_grant | uncore_spc_grant;
   end
endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
module ccx_l15_transducer (
    input                           clk,
    input                           rst_n,
    
    input                           pcx_transducer_req_0,
    input                           pcx_transducer_atomic_req,
    input  [123:117]                pcx_transducer_data_123_117,
    input  [112:0]                  pcx_transducer_data_112_0,
    
    input  [33-1:0]     pcx_transducer_csm,
    
    output [4:0]                    transducer_pcx_grant,
    input                           l15_transducer_ack,
    input                           l15_transducer_header_ack,
    output [4:0]                    transducer_l15_rqtype,
    output [4-1:0]  transducer_l15_amo_op,
    output                          transducer_l15_nc,
    output [2:0]                    transducer_l15_size,
    output [0:0]     transducer_l15_threadid,
    output                          transducer_l15_prefetch,
    output                          transducer_l15_invalidate_cacheline,
    output                          transducer_l15_blockstore,
    output                          transducer_l15_blockinitstore,
    output [1:0]                    transducer_l15_l1rplway,
    output                          transducer_l15_val,
    output [39:0]                   transducer_l15_address,
    output [63:0]                   transducer_l15_data,
    output [63:0]                   transducer_l15_data_next_entry,
    output [33-1:0]     transducer_l15_csm_data,
    
    output reg                      transducer_cpx_data_ready,
    output reg  [144:0]             transducer_cpx_data,
    input                           l15_transducer_val,
    input  [3:0]                    l15_transducer_returntype,
    input                           l15_transducer_l2miss,
    input  [1:0]                    l15_transducer_error,
    input                           l15_transducer_noncacheable,
    input                           l15_transducer_atomic,
    input  [0:0]     l15_transducer_threadid,
    input                           l15_transducer_prefetch,
    input                           l15_transducer_f4b,
    input  [63:0]                   l15_transducer_data_0,
    input  [63:0]                   l15_transducer_data_1,
    input  [63:0]                   l15_transducer_data_2,
    input  [63:0]                   l15_transducer_data_3,
    input                           l15_transducer_inval_icache_all_way,
    input                           l15_transducer_inval_dcache_all_way,
    input  [15:4]                   l15_transducer_inval_address_15_4,
    input                           l15_transducer_cross_invalidate,
    input  [1:0]                    l15_transducer_cross_invalidate_way,
    input                           l15_transducer_inval_dcache_inval,
    input                           l15_transducer_inval_icache_inval,
    input  [1:0]                    l15_transducer_inval_way,
    input                           l15_transducer_blockinitstore,
    output                          transducer_l15_req_ack
);
wire pcxdecoder_pcxbuf_ack;
wire [33-1:0] pcxbuf_pcxdecoder_csm_data;
wire [124-1:0] pcxbuf_pcxdecoder_data;
wire [124-1:0] pcxbuf_pcxdecoder_data_buf1;
wire pcxbuf_pcxdecoder_valid;
wire [4:0] pcx_transducer_req = {4'bx, pcx_transducer_req_0};
wire [123:0] pcx_transducer_data = {pcx_transducer_data_123_117, 4'bx, pcx_transducer_data_112_0};
pcx_buffer pcx_buffer(
    .clk                        (clk),
    .rst_n                      (rst_n),
    .spc_uncore_req             (pcx_transducer_req),
    .spc_uncore_atomic_req      (pcx_transducer_atomic_req),
    .spc_uncore_data            (pcx_transducer_data),
     
    .spc_uncore_csm_data        (pcx_transducer_csm),
     
     
    .pcxdecoder_pcxbuf_ack      (pcxdecoder_pcxbuf_ack),
    .uncore_spc_grant           (transducer_pcx_grant),
    .pcxbuf_pcxdecoder_data     (pcxbuf_pcxdecoder_data),
    .pcxbuf_pcxdecoder_csm_data (pcxbuf_pcxdecoder_csm_data),
    .pcxbuf_pcxdecoder_data_buf1(pcxbuf_pcxdecoder_data_buf1),
    .pcxbuf_pcxdecoder_valid    (pcxbuf_pcxdecoder_valid)
);
pcx_decoder pcx_decoder(
   .clk                                 ( clk                                 ),
   .rst_n                               ( rst_n                               ),
   .pcxbuf_pcxdecoder_data              ( pcxbuf_pcxdecoder_data              ),
   .pcxbuf_pcxdecoder_data_buf1         ( pcxbuf_pcxdecoder_data_buf1         ),
   .pcxbuf_pcxdecoder_csm_data          ( pcxbuf_pcxdecoder_csm_data          ),
   .pcxbuf_pcxdecoder_valid             ( pcxbuf_pcxdecoder_valid             ),
   .l15_pcxdecoder_ack                  ( l15_transducer_ack                  ),
   .l15_pcxdecoder_header_ack           ( l15_transducer_header_ack           ),
   .pcxdecoder_pcxbuf_ack               ( pcxdecoder_pcxbuf_ack               ),
   .pcxdecoder_l15_rqtype               ( transducer_l15_rqtype               ),
   .pcxdecoder_l15_amo_op               ( transducer_l15_amo_op               ),
   .pcxdecoder_l15_nc                   ( transducer_l15_nc                   ),
   .pcxdecoder_l15_size                 ( transducer_l15_size                 ),
   
   .pcxdecoder_l15_threadid             ( transducer_l15_threadid             ),
   .pcxdecoder_l15_prefetch             ( transducer_l15_prefetch             ),
   .pcxdecoder_l15_blockstore           ( transducer_l15_blockstore           ),
   .pcxdecoder_l15_blockinitstore       ( transducer_l15_blockinitstore       ),
   .pcxdecoder_l15_l1rplway             ( transducer_l15_l1rplway             ),
   .pcxdecoder_l15_val                  ( transducer_l15_val                  ),
   .pcxdecoder_l15_invalidate_cacheline ( transducer_l15_invalidate_cacheline ),
   .pcxdecoder_l15_address              ( transducer_l15_address              ),
   .pcxdecoder_l15_csm_data             ( transducer_l15_csm_data             ),
   .pcxdecoder_l15_data                 ( transducer_l15_data                 ),
   .pcxdecoder_l15_data_next_entry      ( transducer_l15_data_next_entry      )
);
wire cpx_data_ready_e;
wire [144:0] cpx_data_e;
always @ (posedge clk)
begin
   if (!rst_n)
   begin
       transducer_cpx_data_ready <= 0;
      
   end
   else
   begin
       transducer_cpx_data_ready <= cpx_data_ready_e;
       transducer_cpx_data <= cpx_data_e;
   end
end
l15_cpxencoder l15_cpxencoder(
    .clk                                (clk),
    .rst_n                              (rst_n),
    .l15_cpxencoder_val                 (l15_transducer_val),
    .l15_cpxencoder_returntype          (l15_transducer_returntype),
    .l15_cpxencoder_l2miss              (l15_transducer_l2miss),
    .l15_cpxencoder_error               (l15_transducer_error),
    .l15_cpxencoder_noncacheable        (l15_transducer_noncacheable),
    .l15_cpxencoder_atomic              (l15_transducer_atomic),
    .l15_cpxencoder_threadid            (l15_transducer_threadid),
    .l15_cpxencoder_prefetch            (l15_transducer_prefetch),
    .l15_cpxencoder_f4b                 (l15_transducer_f4b),
    .l15_cpxencoder_data_0              (l15_transducer_data_0),
    .l15_cpxencoder_data_1              (l15_transducer_data_1),
    .l15_cpxencoder_data_2              (l15_transducer_data_2),
    .l15_cpxencoder_data_3              (l15_transducer_data_3),
    .l15_cpxencoder_inval_icache_all_way(l15_transducer_inval_icache_all_way),
    .l15_cpxencoder_inval_dcache_all_way(l15_transducer_inval_dcache_all_way),
    .l15_cpxencoder_inval_address_15_4  (l15_transducer_inval_address_15_4),
    .l15_cpxencoder_cross_invalidate    (l15_transducer_cross_invalidate),
    .l15_cpxencoder_cross_invalidate_way(l15_transducer_cross_invalidate_way),
    .l15_cpxencoder_inval_dcache_inval  (l15_transducer_inval_dcache_inval),
    .l15_cpxencoder_inval_icache_inval  (l15_transducer_inval_icache_inval),
    .l15_cpxencoder_inval_way           (l15_transducer_inval_way),
    .l15_cpxencoder_blockinitstore      (l15_transducer_blockinitstore),
    .uncore_spc_data_ready              (cpx_data_ready_e),
    .uncore_spc_data                    (cpx_data_e),
    .cpxencoder_l15_req_ack             (transducer_l15_req_ack)
);
endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
  
          
      
    
         
module tile #(
     parameter TILE_TYPE = 0
) (
    input                               clk,
    input                               rst_n,    
    input                               clk_en,   
    input wire [14-1:0]  default_chipid,
    input wire [8-1:0]       default_coreid_x,
    input wire [8-1:0]       default_coreid_y,
    input wire [8-1:0] flat_tileid,
    
    input                               jtag_tiles_ucb_val,
    input [4-1:0]          jtag_tiles_ucb_data,
    output                              tile_jtag_ucb_val,
    output [4-1:0]         tile_jtag_ucb_data,
    
    input [64-1:0]         dyn0_dataIn_N,
    input [64-1:0]         dyn0_dataIn_E,
    input [64-1:0]         dyn0_dataIn_W,
    input [64-1:0]         dyn0_dataIn_S,
    input                               dyn0_validIn_N,
    input                               dyn0_validIn_E,
    input                               dyn0_validIn_W,
    input                               dyn0_validIn_S,
    input                               dyn0_dNo_yummy,
    input                               dyn0_dEo_yummy,
    input                               dyn0_dWo_yummy,
    input                               dyn0_dSo_yummy,
    
    input [64-1:0]         dyn1_dataIn_N,
    input [64-1:0]         dyn1_dataIn_E,
    input [64-1:0]         dyn1_dataIn_W,
    input [64-1:0]         dyn1_dataIn_S,
    input                               dyn1_validIn_N,
    input                               dyn1_validIn_E,
    input                               dyn1_validIn_W,
    input                               dyn1_validIn_S,
    input                               dyn1_dNo_yummy,
    input                               dyn1_dEo_yummy,
    input                               dyn1_dWo_yummy,
    input                               dyn1_dSo_yummy,
    
    input [64-1:0]         dyn2_dataIn_N,
    input [64-1:0]         dyn2_dataIn_E,
    input [64-1:0]         dyn2_dataIn_W,
    input [64-1:0]         dyn2_dataIn_S,
    input                               dyn2_validIn_N,
    input                               dyn2_validIn_E,
    input                               dyn2_validIn_W,
    input                               dyn2_validIn_S,
    input                               dyn2_dNo_yummy,
    input                               dyn2_dEo_yummy,
    input                               dyn2_dWo_yummy,
    input                               dyn2_dSo_yummy,
    
    output [64-1:0]        dyn0_dNo,
    output [64-1:0]        dyn0_dEo,
    output [64-1:0]        dyn0_dWo,
    output [64-1:0]        dyn0_dSo,
    output                              dyn0_dNo_valid,
    output                              dyn0_dEo_valid,
    output                              dyn0_dWo_valid,
    output                              dyn0_dSo_valid,
    output                              dyn0_yummyOut_N,
    output                              dyn0_yummyOut_E,
    output                              dyn0_yummyOut_W,
    output                              dyn0_yummyOut_S,
    
    
    output [64-1:0]        dyn1_dNo,
    output [64-1:0]        dyn1_dEo,
    output [64-1:0]        dyn1_dWo,
    output [64-1:0]        dyn1_dSo,
    output                              dyn1_dNo_valid,
    output                              dyn1_dEo_valid,
    output                              dyn1_dWo_valid,
    output                              dyn1_dSo_valid,
    output                              dyn1_yummyOut_N,
    output                              dyn1_yummyOut_E,
    output                              dyn1_yummyOut_W,
    output                              dyn1_yummyOut_S,
    
    
    output [64-1:0]        dyn2_dNo,
    output [64-1:0]        dyn2_dEo,
    output [64-1:0]        dyn2_dWo,
    output [64-1:0]        dyn2_dSo,
    output                              dyn2_dNo_valid,
    output                              dyn2_dEo_valid,
    output                              dyn2_dWo_valid,
    output                              dyn2_dSo_valid,
    output                              dyn2_yummyOut_N,
    output                              dyn2_yummyOut_E,
    output                              dyn2_yummyOut_W,
    output                              dyn2_yummyOut_S
    
    ,
    
    input                               debug_req_i,   
    output                              unavailable_o, 
    
    input                               timer_irq_i,   
    input                               ipi_i,         
    
    input   [1:0]                       irq_i          
);
    
    wire clk_gated;
    clk_gating_latch clk_gating_latch(
        .clk(clk),
        .clk_en(clk_en),
        .clk_out(clk_gated)
    );
    
    reg rst_n_f;
    always @ (posedge clk)
    begin
      rst_n_f <= rst_n;
    end
    
    wire [14-1:0]        config_chipid;
    wire [8-1:0]             config_coreid_x;
    wire [8-1:0]             config_coreid_y;
    wire [64-1:0]              buffer_processor_data_noc1;
    wire [64-1:0]              buffer_processor_data_noc2;
    wire [64-1:0]              buffer_processor_data_noc3;
    wire                                buffer_processor_valid_noc1;
    wire                                buffer_processor_valid_noc2;
    wire                                buffer_processor_valid_noc3;
    wire                                processor_router_ready_noc1;
    wire                                processor_router_ready_noc2;
    wire                                processor_router_ready_noc3;
    wire                                router_processor_ready_noc1;
    wire                                router_processor_ready_noc2;
    wire                                router_processor_ready_noc3;
    
    wire [64-1:0]          processor_router_data_noc1;
    wire                                processor_router_valid_noc1;
    wire                                buffer_router_yummy_noc1;
    wire [64-1:0]          buffer_router_data_noc1;
    wire                                buffer_router_valid_noc1;
    wire [64-1:0]          processor_router_data_noc2;
    wire                                processor_router_valid_noc2;
    wire                                buffer_router_yummy_noc2;
    wire [64-1:0]          buffer_router_data_noc2;
    wire                                buffer_router_valid_noc2;
    wire [64-1:0]          processor_router_data_noc3;
    wire                                processor_router_valid_noc3;
    wire                                buffer_router_yummy_noc3;
    wire [64-1:0]          buffer_router_data_noc3;
    wire                                buffer_router_valid_noc3;
    wire [64-1:0]          router_buffer_data_noc1;
    wire                                router_buffer_data_val_noc1;
    wire                                router_buffer_consumed_noc1;
    wire                                thanksIn_CGNO0;
    wire [64-1:0]          router_buffer_data_noc2;
    wire                                router_buffer_data_val_noc2;
    wire                                router_buffer_consumed_noc2;
    wire                                thanksIn_CGNO1;
    wire [64-1:0]          router_buffer_data_noc3;
    wire                                router_buffer_data_val_noc3;
    wire                                router_buffer_consumed_noc3;
    wire                                thanksIn_CGNO2;
    wire   [4:0]                        pcx_transducer_req;
    wire                                pcx_transducer_atomic_req;
    wire   [123:0]                      pcx_transducer_data;
    
    wire   [32:0]                   pcx_transducer_csm;
    
    wire [4:0]                          transducer_pcx_grant;
    
    wire                                transducer_cpx_data_ready;
    wire [144:0]                        transducer_cpx_data;
    wire                                spc_grst_l;
    wire                                cpx_arb_spc_data_rdy;
    wire [144:0]                        cpx_arb_spc_data;
    wire [4:0]                          cpx_arb_spc_grant;
    wire [5-1:0]       transducer_l15_rqtype;
    wire [4-1:0]        transducer_l15_amo_op;
    wire                                transducer_l15_nc;
    wire [3-1:0]    transducer_l15_size;
    wire [0:0]           transducer_l15_threadid;
    wire                                transducer_l15_prefetch;
    wire                                transducer_l15_invalidate_cacheline;
    wire                                transducer_l15_blockstore;
    wire                                transducer_l15_blockinitstore;
    wire [1:0]                          transducer_l15_l1rplway;
    wire                                transducer_l15_val;
    wire [39:0]              transducer_l15_address;
    wire [63:0]                         transducer_l15_data;
    wire [63:0]                         transducer_l15_data_next_entry;
    wire [33-1:0]           transducer_l15_csm_data;
    wire                                l15_transducer_ack;
    wire                                l15_transducer_header_ack;
    wire                                l15_transducer_val;
    wire [3:0]                          l15_transducer_returntype;
    wire                                l15_transducer_l2miss;
    wire [1:0]                          l15_transducer_error;
    wire                                l15_transducer_noncacheable;
    wire                                l15_transducer_atomic;
    wire [0:0]           l15_transducer_threadid;
    wire                                l15_transducer_prefetch;
    wire                                l15_transducer_f4b;
    wire [63:0]                         l15_transducer_data_0;
    wire [63:0]                         l15_transducer_data_1;
    wire [63:0]                         l15_transducer_data_2;
    wire [63:0]                         l15_transducer_data_3;
    wire                                l15_transducer_inval_icache_all_way;
    wire                                l15_transducer_inval_dcache_all_way;
    wire [15:4]                         l15_transducer_inval_address_15_4;
    wire                                l15_transducer_cross_invalidate;
    wire [1:0]                          l15_transducer_cross_invalidate_way;
    wire                                l15_transducer_inval_dcache_inval;
    wire                                l15_transducer_inval_icache_inval;
    wire [1:0]                          l15_transducer_inval_way;
    wire                                l15_transducer_blockinitstore;
    wire                                transducer_l15_req_ack;
    wire [94-1:0] core_rtap_data;
    wire rtap_core_val;
    wire [1:0] rtap_core_threadid;
    wire [4-1:0]  rtap_core_id;
    wire [94-1:0] rtap_core_data;
    
    
    wire [144:0]                        fpu_arb_data;
    wire                                fpu_arb_data_rdy;
    wire                                fpu_arb_grant;
    wire                                l15_dmbr_l1missIn;
    wire [4-1:0]          l15_dmbr_l1missTag;
    wire                                l15_dmbr_l2responseIn;
    wire                                l15_dmbr_l2missIn;
    wire [4-1:0]          l15_dmbr_l2missTag;
    wire                                dmbr_l15_stall; 
    wire                                l15_config_req_val_s2;
    wire                                l15_config_req_rw_s2;
    wire [63:0]                         l15_config_write_req_data_s2;
    wire [15:8]     l15_config_req_address_s2;
    wire [63:0]                         config_l15_read_res_data_s3;
    wire                                config_dmbr_func_en;
    wire                                config_dmbr_stall_en;
    wire                                config_dmbr_proc_ld;
    wire [16-1:0]         config_dmbr_replenish_cycles;
    wire [10-1:0]             config_dmbr_bin_scale;
    wire [6-1:0] config_dmbr_cred_bin_0;
wire [6-1:0] config_dmbr_cred_bin_1;
wire [6-1:0] config_dmbr_cred_bin_2;
wire [6-1:0] config_dmbr_cred_bin_3;
wire [6-1:0] config_dmbr_cred_bin_4;
wire [6-1:0] config_dmbr_cred_bin_5;
wire [6-1:0] config_dmbr_cred_bin_6;
wire [6-1:0] config_dmbr_cred_bin_7;
wire [6-1:0] config_dmbr_cred_bin_8;
wire [6-1:0] config_dmbr_cred_bin_9;
    wire [6-1:0] from_dmbr_cred_bin_0;
wire [6-1:0] from_dmbr_cred_bin_1;
wire [6-1:0] from_dmbr_cred_bin_2;
wire [6-1:0] from_dmbr_cred_bin_3;
wire [6-1:0] from_dmbr_cred_bin_4;
wire [6-1:0] from_dmbr_cred_bin_5;
wire [6-1:0] from_dmbr_cred_bin_6;
wire [6-1:0] from_dmbr_cred_bin_7;
wire [6-1:0] from_dmbr_cred_bin_8;
wire [6-1:0] from_dmbr_cred_bin_9;
    wire                                config_csm_en;
    wire [31:0]                         config_system_tile_count;
    wire [2-1:0] config_home_alloc_method;
    wire [22-1:0] config_hmt_base;
    
    wire [4-1:0] srams_rtap_data;
    wire [4-1:0] rtap_srams_bist_command;
    wire [4-1:0] rtap_srams_bist_data;
    wire [4-1:0] l15_rtap_data;
    wire [4-1:0] sparc_rtap_data;
    wire [4-1:0] l2_rtap_data;
    wire [3:0] rtap_lsu_ctlbits_wr_en;
    wire [13:0] rtap_lsu_ctlbits_data;
    wire        rtap_arb_req_val;
    wire [63:0] rtap_arb_req_data;
    wire [1:0]  rtap_arb_req_threadid;
    
    wire rtap_config_req_val;
    wire rtap_config_req_rw;
    wire [63:0] rtap_config_write_req_data;
    wire [15:8] rtap_config_req_address;
    wire [63:0] config_rtap_read_res_data;
    
    
    
    
    
    
    dynamic_node_top_wrap user_dynamic_network0
      (.clk(clk_gated),
       .reset_in(~rst_n_f),
       
       .dataIn_N(dyn0_dataIn_N),
       .dataIn_E(dyn0_dataIn_E),
       .dataIn_S(dyn0_dataIn_S),
       .dataIn_W(dyn0_dataIn_W),
       .dataIn_P(buffer_router_data_noc1),
       
       .validIn_N(dyn0_validIn_N),
       .validIn_E(dyn0_validIn_E),
       .validIn_S(dyn0_validIn_S),
       .validIn_W(dyn0_validIn_W),
       .validIn_P(buffer_router_valid_noc1),
       
       .yummyIn_N(dyn0_dNo_yummy),
       .yummyIn_E(dyn0_dEo_yummy),
       .yummyIn_S(dyn0_dSo_yummy),
       .yummyIn_W(dyn0_dWo_yummy),
       .yummyIn_P(buffer_router_yummy_noc1),
       
       .myLocX(config_coreid_x),
       .myLocY(config_coreid_y),
       .myChipID(config_chipid),
       
       
       
       
       .dataOut_N(dyn0_dNo),
       .dataOut_E(dyn0_dEo),
       .dataOut_S(dyn0_dSo),
       .dataOut_W(dyn0_dWo),
       .dataOut_P(router_buffer_data_noc1), 
       
       .validOut_N(dyn0_dNo_valid),
       .validOut_E(dyn0_dEo_valid),
       .validOut_S(dyn0_dSo_valid),
       .validOut_W(dyn0_dWo_valid),
       .validOut_P(router_buffer_data_val_noc1), 
       
       .yummyOut_N(dyn0_yummyOut_N),
       .yummyOut_E(dyn0_yummyOut_E),
       .yummyOut_W(dyn0_yummyOut_W),
       .yummyOut_S(dyn0_yummyOut_S),
       .yummyOut_P(router_buffer_consumed_noc1), 
       
       .thanksIn_P(thanksIn_CGNO0));
       
       
       
       
    dynamic_node_top_wrap user_dynamic_network1
      (.clk(clk_gated),
       .reset_in(~rst_n_f),
       
       .dataIn_N(dyn1_dataIn_N),
       .dataIn_E(dyn1_dataIn_E),
       .dataIn_S(dyn1_dataIn_S),
       .dataIn_W(dyn1_dataIn_W),
       .dataIn_P(buffer_router_data_noc2),
       
       .validIn_N(dyn1_validIn_N),
       .validIn_E(dyn1_validIn_E),
       .validIn_S(dyn1_validIn_S),
       .validIn_W(dyn1_validIn_W),
       .validIn_P(buffer_router_valid_noc2),
       
       .yummyIn_N(dyn1_dNo_yummy),
       .yummyIn_E(dyn1_dEo_yummy),
       .yummyIn_S(dyn1_dSo_yummy),
       .yummyIn_W(dyn1_dWo_yummy),
       .yummyIn_P(buffer_router_yummy_noc2),
       
       .myLocX(config_coreid_x),
       .myLocY(config_coreid_y),
       .myChipID(config_chipid),
       
       
       
       
       .dataOut_N(dyn1_dNo),
       .dataOut_E(dyn1_dEo),
       .dataOut_S(dyn1_dSo),
       .dataOut_W(dyn1_dWo),
       .dataOut_P(router_buffer_data_noc2), 
       
       .validOut_N(dyn1_dNo_valid),
       .validOut_E(dyn1_dEo_valid),
       .validOut_S(dyn1_dSo_valid),
       .validOut_W(dyn1_dWo_valid),
       .validOut_P(router_buffer_data_val_noc2), 
       
       .yummyOut_N(dyn1_yummyOut_N),
       .yummyOut_E(dyn1_yummyOut_E),
       .yummyOut_W(dyn1_yummyOut_W),
       .yummyOut_S(dyn1_yummyOut_S),
       .yummyOut_P(router_buffer_consumed_noc2), 
       
       .thanksIn_P(thanksIn_CGNO1));
       
       
       
       
    dynamic_node_top_wrap user_dynamic_network2
      (.clk(clk_gated),
       .reset_in(~rst_n_f),
       
       .dataIn_N(dyn2_dataIn_N),
       .dataIn_E(dyn2_dataIn_E),
       .dataIn_S(dyn2_dataIn_S),
       .dataIn_W(dyn2_dataIn_W),
       .dataIn_P(buffer_router_data_noc3),
       
       .validIn_N(dyn2_validIn_N),
       .validIn_E(dyn2_validIn_E),
       .validIn_S(dyn2_validIn_S),
       .validIn_W(dyn2_validIn_W),
       .validIn_P(buffer_router_valid_noc3),
       
       .yummyIn_N(dyn2_dNo_yummy),
       .yummyIn_E(dyn2_dEo_yummy),
       .yummyIn_S(dyn2_dSo_yummy),
       .yummyIn_W(dyn2_dWo_yummy),
       .yummyIn_P(buffer_router_yummy_noc3),
       
       .myLocX(config_coreid_x),
       .myLocY(config_coreid_y),
       .myChipID(config_chipid),
       
       
       
       
       .dataOut_N(dyn2_dNo),
       .dataOut_E(dyn2_dEo),
       .dataOut_S(dyn2_dSo),
       .dataOut_W(dyn2_dWo),
       .dataOut_P(router_buffer_data_noc3), 
       
       .validOut_N(dyn2_dNo_valid),
       .validOut_E(dyn2_dEo_valid),
       .validOut_S(dyn2_dSo_valid),
       .validOut_W(dyn2_dWo_valid),
       .validOut_P(router_buffer_data_val_noc3), 
       
       .yummyOut_N(dyn2_yummyOut_N),
       .yummyOut_E(dyn2_yummyOut_E),
       .yummyOut_W(dyn2_yummyOut_W),
       .yummyOut_S(dyn2_yummyOut_S),
       .yummyOut_P(router_buffer_consumed_noc3), 
       
       .thanksIn_P(thanksIn_CGNO2));
       
       
       
       
    
    
    
    valrdy_to_credit #(16, 5) cgno_blk1(
        .clk(clk_gated),
        .reset(~rst_n_f),
        .data_in(processor_router_data_noc1),
        .valid_in(processor_router_valid_noc1),
        .ready_in(router_processor_ready_noc1),
        .data_out(buffer_router_data_noc1),           
        .valid_out(buffer_router_valid_noc1),       
        .yummy_out(router_buffer_consumed_noc1)    
    );
    valrdy_to_credit #(16, 5) cgno_blk2(
        .clk(clk_gated),
        .reset(~rst_n_f),
        .data_in(processor_router_data_noc2),
        .valid_in(processor_router_valid_noc2),
        .ready_in(router_processor_ready_noc2),
        .data_out(buffer_router_data_noc2),           
        .valid_out(buffer_router_valid_noc2),       
        .yummy_out(router_buffer_consumed_noc2)    
    );
    valrdy_to_credit #(16, 5) cgno_blk3(
        .clk(clk_gated),
        .reset(~rst_n_f),
        .data_in(processor_router_data_noc3),
        .valid_in(processor_router_valid_noc3),
        .ready_in(router_processor_ready_noc3),
        .data_out(buffer_router_data_noc3),           
        .valid_out(buffer_router_valid_noc3),       
        .yummy_out(router_buffer_consumed_noc3)    
    );
    credit_to_valrdy cgni_blk1(
        .clk(clk_gated),
        .reset(~rst_n_f),
        .data_in(router_buffer_data_noc1),
        .valid_in(router_buffer_data_val_noc1),
        .yummy_in(buffer_router_yummy_noc1),
        .data_out(buffer_processor_data_noc1),           
        .valid_out(buffer_processor_valid_noc1),       
        .ready_out(processor_router_ready_noc1)    
    );
    credit_to_valrdy cgni_blk2(
        .clk(clk_gated),
        .reset(~rst_n_f),
        .data_in(router_buffer_data_noc2),
        .valid_in(router_buffer_data_val_noc2),
        .yummy_in(buffer_router_yummy_noc2),
        .data_out(buffer_processor_data_noc2),           
        .valid_out(buffer_processor_valid_noc2),       
        .ready_out(processor_router_ready_noc2)    
    );
    credit_to_valrdy cgni_blk3(
        .clk(clk_gated),
        .reset(~rst_n_f),
        .data_in(router_buffer_data_noc3),
        .valid_in(router_buffer_data_val_noc3),
        .yummy_in(buffer_router_yummy_noc3),
        .data_out(buffer_processor_data_noc3),           
        .valid_out(buffer_processor_valid_noc3),       
        .ready_out(processor_router_ready_noc3)    
    );
generate
if (TILE_TYPE == 0) begin : g_sparc_core
       
       
        
        
 
end
endgenerate
generate
if (TILE_TYPE == 1) begin : g_picorv32_core
 
end
endgenerate
generate
if (TILE_TYPE == 2) begin : g_ariane_core
    
    
    
    
    
    wire [(14 + 40 + 2*64 +      
                        5  + 
                        1 + 
                        2      + 
                        33 )-1:0]  l15_req;
    wire [(16 + 4*64 + (15 - 4 + 1) + 
                        4  +      
                        1 +      
                        2 * 2)-1:0] l15_rtrn;
    
    
    assign l15_rtrn = { l15_transducer_ack,
                        l15_transducer_header_ack,
                        l15_transducer_val,
                        l15_transducer_returntype,
                        l15_transducer_l2miss,
                        l15_transducer_error,
                        l15_transducer_noncacheable,
                        l15_transducer_atomic,
                        l15_transducer_threadid,
                        l15_transducer_prefetch,
                        l15_transducer_f4b,
                        l15_transducer_data_0,
                        l15_transducer_data_1,
                        l15_transducer_data_2,
                        l15_transducer_data_3,
                        l15_transducer_inval_icache_all_way,
                        l15_transducer_inval_dcache_all_way,
                        l15_transducer_inval_address_15_4,
                        l15_transducer_cross_invalidate,
                        l15_transducer_cross_invalidate_way,
                        l15_transducer_inval_dcache_inval,
                        l15_transducer_inval_icache_inval,
                        l15_transducer_inval_way,
                        l15_transducer_blockinitstore };
    wire [2:0] transducer_l15_size_pcx_standard;
    
    
    assign { transducer_l15_val,
             transducer_l15_req_ack,
             transducer_l15_rqtype,
             transducer_l15_nc,
             transducer_l15_size_pcx_standard,
             transducer_l15_threadid,
             transducer_l15_prefetch,
             transducer_l15_invalidate_cacheline,
             transducer_l15_blockstore,
             transducer_l15_blockinitstore,
             transducer_l15_l1rplway,
             transducer_l15_address,
             transducer_l15_data,
             transducer_l15_data_next_entry,
             transducer_l15_csm_data,
             transducer_l15_amo_op} = l15_req;
    
    
    assign transducer_l15_size = (transducer_l15_size_pcx_standard == 3'b000) ? 3'b001 :
                                    (transducer_l15_size_pcx_standard == 3'b001) ? 3'b010 : 
                                    (transducer_l15_size_pcx_standard == 3'b010) ? 3'b011 : 
                                    (transducer_l15_size_pcx_standard == 3'b011) ? 3'b100 : 
                                    (transducer_l15_size_pcx_standard == 3'b111 && 
                                     transducer_l15_rqtype == 5'b10000 && 
                                    ~transducer_l15_invalidate_cacheline) ? 3'b110 : 3'b101; 
    wire [63:0] ariane_bootaddr;
    assign ariane_bootaddr  =  64'h0;
    ariane_verilog_wrap #(
        .DmBaseAddress          ( 64'h0 ),
        .SwapEndianess          ( 1'b1 ),
        .NrExecuteRegionRules   ( 0   ),
        .ExecuteRegionAddrBase  (    ),
        .ExecuteRegionLength    (    ),
        .NrCachedRegionRules    (  1   ),
        .CachedRegionAddrBase   ( {64'h0} ),
        .CachedRegionLength     ( {64'h0} )
    ) core (
        .clk_i       ( clk_gated              ),
        .reset_l     ( rst_n_f                ),
        .spc_grst_l  ( spc_grst_l             ),
        .boot_addr_i ( ariane_bootaddr        ),
        .hart_id_i   ( {{64-8{1'b0}}, flat_tileid} ),
        .irq_i       ( irq_i                  ),
        .ipi_i       ( ipi_i                  ),
        .time_irq_i  ( timer_irq_i            ),
        .debug_req_i ( debug_req_i            ),
        .l15_req_o   ( l15_req                ),
        .l15_rtrn_i  ( l15_rtrn               )
    );
    assign unavailable_o = 1'b0;
 
  end
  endgenerate
    
    
    
    l15_wrap l15(
        .clk(clk_gated),
        .rst_n(spc_grst_l),
        .transducer_l15_rqtype              (transducer_l15_rqtype),
        .transducer_l15_amo_op              (transducer_l15_amo_op),
        .transducer_l15_nc                  (transducer_l15_nc),
        .transducer_l15_size                (transducer_l15_size),
        
        .transducer_l15_threadid            (transducer_l15_threadid),
        .transducer_l15_prefetch            (transducer_l15_prefetch),
        .transducer_l15_blockstore          (transducer_l15_blockstore),
        .transducer_l15_blockinitstore      (transducer_l15_blockinitstore),
        .transducer_l15_l1rplway            (transducer_l15_l1rplway),
        .transducer_l15_val                 (transducer_l15_val),
        .transducer_l15_invalidate_cacheline(transducer_l15_invalidate_cacheline),
        .transducer_l15_address             (transducer_l15_address),
        .transducer_l15_csm_data            (transducer_l15_csm_data),
        .transducer_l15_data                (transducer_l15_data),
        .transducer_l15_data_next_entry     (transducer_l15_data_next_entry),
        .l15_transducer_ack                 (l15_transducer_ack),
        .l15_transducer_header_ack          (l15_transducer_header_ack),
        .l15_transducer_val                 (l15_transducer_val),
        .l15_transducer_returntype          (l15_transducer_returntype),
        .l15_transducer_l2miss              (l15_transducer_l2miss),
        .l15_transducer_error               (l15_transducer_error),
        .l15_transducer_noncacheable        (l15_transducer_noncacheable),
        .l15_transducer_atomic              (l15_transducer_atomic),
        .l15_transducer_threadid            (l15_transducer_threadid),
        .l15_transducer_prefetch            (l15_transducer_prefetch),
        .l15_transducer_f4b                 (l15_transducer_f4b),
        .l15_transducer_data_0              (l15_transducer_data_0),
        .l15_transducer_data_1              (l15_transducer_data_1),
        .l15_transducer_data_2              (l15_transducer_data_2),
        .l15_transducer_data_3              (l15_transducer_data_3),
        .l15_transducer_inval_icache_all_way(l15_transducer_inval_icache_all_way),
        .l15_transducer_inval_dcache_all_way(l15_transducer_inval_dcache_all_way),
        .l15_transducer_inval_address_15_4  (l15_transducer_inval_address_15_4),
        .l15_transducer_cross_invalidate    (l15_transducer_cross_invalidate),
        .l15_transducer_cross_invalidate_way(l15_transducer_cross_invalidate_way),
        .l15_transducer_inval_dcache_inval  (l15_transducer_inval_dcache_inval),
        .l15_transducer_inval_icache_inval  (l15_transducer_inval_icache_inval),
        .l15_transducer_inval_way           (l15_transducer_inval_way),
        .l15_transducer_blockinitstore      (l15_transducer_blockinitstore),
        .transducer_l15_req_ack             (transducer_l15_req_ack),
        .noc1_out_rdy(router_processor_ready_noc1),
        .noc2_in_val(buffer_processor_valid_noc2),
        .noc2_in_data(buffer_processor_data_noc2),
        .noc3_out_rdy(router_processor_ready_noc3),
        .dmbr_l15_stall(dmbr_l15_stall),
        .chipid(config_chipid),
        .coreid_x(config_coreid_x),
        .coreid_y(config_coreid_y),
        .noc1_out_val(processor_router_valid_noc1),
        .noc1_out_data(processor_router_data_noc1),
        .noc2_in_rdy(processor_router_ready_noc2),
        .noc3_out_val(processor_router_valid_noc3),
        .noc3_out_data(processor_router_data_noc3),
        .l15_dmbr_l1missIn(l15_dmbr_l1missIn),
        .l15_dmbr_l1missTag(l15_dmbr_l1missTag),
        .l15_dmbr_l2missIn(l15_dmbr_l2missIn),
        .l15_dmbr_l2missTag(l15_dmbr_l2missTag),
        .l15_dmbr_l2responseIn(l15_dmbr_l2responseIn),
        
        .l15_config_req_val_s2(l15_config_req_val_s2),
        .l15_config_req_rw_s2(l15_config_req_rw_s2),
        .l15_config_write_req_data_s2(l15_config_write_req_data_s2),
        .l15_config_req_address_s2(l15_config_req_address_s2),
        .config_l15_read_res_data_s3(config_l15_read_res_data_s3),
        
        .config_csm_en(config_csm_en),
        .config_hmt_base(config_hmt_base),
        .config_system_tile_count_5_0(config_system_tile_count[5:0]),
        .config_home_alloc_method(config_home_alloc_method),
        
        .srams_rtap_data (l15_rtap_data),
        .rtap_srams_bist_command (rtap_srams_bist_command),
        .rtap_srams_bist_data (rtap_srams_bist_data)
    );
    
    
    
    dmbr dmbr_ins (
        .clk                  (clk_gated                      ),
        .rst                  (~spc_grst_l              ),
        .func_en              (config_dmbr_func_en      ),
        .stall_en             (config_dmbr_stall_en     ),
        
        .proc_ld              (config_dmbr_proc_ld      ),
        
        
        
        .creditIn_0		(config_dmbr_cred_bin_0),
.creditIn_1		(config_dmbr_cred_bin_1),
.creditIn_2		(config_dmbr_cred_bin_2),
.creditIn_3		(config_dmbr_cred_bin_3),
.creditIn_4		(config_dmbr_cred_bin_4),
.creditIn_5		(config_dmbr_cred_bin_5),
.creditIn_6		(config_dmbr_cred_bin_6),
.creditIn_7		(config_dmbr_cred_bin_7),
.creditIn_8		(config_dmbr_cred_bin_8),
.creditIn_9		(config_dmbr_cred_bin_9),
        
        .replenishCyclesIn    (config_dmbr_replenish_cycles ),
        
        .binScaleIn           (config_dmbr_bin_scale        ),
        
        .l1missIn             (l15_dmbr_l1missIn            ),
        .l1missTag            (l15_dmbr_l1missTag           ),
        
        .l2missIn             (l15_dmbr_l2missIn            ),
        .l2missTag            (l15_dmbr_l2missTag           ),
        .l2responseIn         (l15_dmbr_l2responseIn        ),
        
        .curr_cred_bin_0			(from_dmbr_cred_bin_0),
.curr_cred_bin_1			(from_dmbr_cred_bin_1),
.curr_cred_bin_2			(from_dmbr_cred_bin_2),
.curr_cred_bin_3			(from_dmbr_cred_bin_3),
.curr_cred_bin_4			(from_dmbr_cred_bin_4),
.curr_cred_bin_5			(from_dmbr_cred_bin_5),
.curr_cred_bin_6			(from_dmbr_cred_bin_6),
.curr_cred_bin_7			(from_dmbr_cred_bin_7),
.curr_cred_bin_8			(from_dmbr_cred_bin_8),
.curr_cred_bin_9			(from_dmbr_cred_bin_9),
        .stallOut             (dmbr_l15_stall           )
    );
    
    
    
    l2 l2(
        .clk(clk_gated),
        .rst_n(rst_n_f),
        .chipid(config_chipid),
        .coreid_x(config_coreid_x),
        .coreid_y(config_coreid_y),
        .noc1_valid_in(buffer_processor_valid_noc1),
        .noc3_valid_in(buffer_processor_valid_noc3),
        .noc1_data_in(buffer_processor_data_noc1),
        .noc3_data_in(buffer_processor_data_noc3),
        .noc2_ready_out(router_processor_ready_noc2),
        .noc1_ready_in(processor_router_ready_noc1),
        .noc3_ready_in(processor_router_ready_noc3),
        .noc2_valid_out(processor_router_valid_noc2),
        .noc2_data_out(processor_router_data_noc2),
        
        .srams_rtap_data (l2_rtap_data),
        .rtap_srams_bist_command (rtap_srams_bist_command),
        .rtap_srams_bist_data (rtap_srams_bist_data)
    );
    
    
    
    config_regs uncore_config(
        .clk                          (clk_gated                          ),
        .rst_n                        (rst_n_f                        ),
        .l15_config_req_val_s2        (l15_config_req_val_s2        ),
        .l15_config_req_rw_s2         (l15_config_req_rw_s2         ),
        .l15_config_write_req_data_s2 (l15_config_write_req_data_s2 ),
        .l15_config_req_address_s2    (l15_config_req_address_s2    ),
        .config_l15_read_res_data_s3  (config_l15_read_res_data_s3  ),
        .default_chipid               (default_chipid               ),
        .default_coreid_x             (default_coreid_x             ),
        .default_coreid_y             (default_coreid_y             ),
        .config_hmt_base              (config_hmt_base              ),
        .config_dmbr_func_en          (config_dmbr_func_en          ),
        .config_dmbr_stall_en         (config_dmbr_stall_en         ),
        .config_dmbr_proc_ld          (config_dmbr_proc_ld          ),
        .config_dmbr_replenish_cycles (config_dmbr_replenish_cycles ),
        .config_dmbr_bin_scale        (config_dmbr_bin_scale        ),
        
        .config_dmbr_cred_bin_0			(config_dmbr_cred_bin_0),
.config_dmbr_cred_bin_1			(config_dmbr_cred_bin_1),
.config_dmbr_cred_bin_2			(config_dmbr_cred_bin_2),
.config_dmbr_cred_bin_3			(config_dmbr_cred_bin_3),
.config_dmbr_cred_bin_4			(config_dmbr_cred_bin_4),
.config_dmbr_cred_bin_5			(config_dmbr_cred_bin_5),
.config_dmbr_cred_bin_6			(config_dmbr_cred_bin_6),
.config_dmbr_cred_bin_7			(config_dmbr_cred_bin_7),
.config_dmbr_cred_bin_8			(config_dmbr_cred_bin_8),
.config_dmbr_cred_bin_9			(config_dmbr_cred_bin_9),
        
        .from_dmbr_cred_bin_0			(from_dmbr_cred_bin_0),
.from_dmbr_cred_bin_1			(from_dmbr_cred_bin_1),
.from_dmbr_cred_bin_2			(from_dmbr_cred_bin_2),
.from_dmbr_cred_bin_3			(from_dmbr_cred_bin_3),
.from_dmbr_cred_bin_4			(from_dmbr_cred_bin_4),
.from_dmbr_cred_bin_5			(from_dmbr_cred_bin_5),
.from_dmbr_cred_bin_6			(from_dmbr_cred_bin_6),
.from_dmbr_cred_bin_7			(from_dmbr_cred_bin_7),
.from_dmbr_cred_bin_8			(from_dmbr_cred_bin_8),
.from_dmbr_cred_bin_9			(from_dmbr_cred_bin_9),
        .config_csm_en                (config_csm_en                ),
        .config_system_tile_count     (config_system_tile_count     ),
        .config_home_alloc_method     (config_home_alloc_method     ),
        .config_chipid                (config_chipid                ),
        .config_coreid_x              (config_coreid_x              ),
        .config_coreid_y              (config_coreid_y              ),
        
        .rtap_config_req_val (rtap_config_req_val),
        .rtap_config_req_rw (rtap_config_req_rw),
        .rtap_config_write_req_data (rtap_config_write_req_data),
        .rtap_config_req_address (rtap_config_req_address),
        .config_rtap_read_res_data (config_rtap_read_res_data)
    );
    
    
    assign srams_rtap_data = l15_rtap_data
                                | sparc_rtap_data
                                | l2_rtap_data;
    rtap rtap(
        .clk(clk_gated),
        .rst_n(rst_n_f),
        .own_tileid(flat_tileid),
        
        .tile_jtag_ucb_val(tile_jtag_ucb_val),
        .tile_jtag_ucb_data(tile_jtag_ucb_data),
        .jtag_tiles_ucb_val(jtag_tiles_ucb_val),
        .jtag_tiles_ucb_data(jtag_tiles_ucb_data),
        
        .srams_rtap_data (srams_rtap_data),
        .rtap_srams_bist_command (rtap_srams_bist_command),
        .rtap_srams_bist_data (rtap_srams_bist_data),
        
        .rtap_arb_req_val (rtap_arb_req_val),
        .rtap_arb_req_data (rtap_arb_req_data),
        .rtap_arb_req_threadid (rtap_arb_req_threadid),
        
        .rtap_config_req_val (rtap_config_req_val),
        .rtap_config_req_rw (rtap_config_req_rw),
        .rtap_config_write_req_data (rtap_config_write_req_data),
        .rtap_config_req_address (rtap_config_req_address),
        .config_rtap_read_res_data (config_rtap_read_res_data),
        .core_rtap_data          (core_rtap_data),
        .rtap_core_val         (rtap_core_val),
        .rtap_core_threadid         (rtap_core_threadid),
        .rtap_core_id         (rtap_core_id),
        .rtap_core_data         (rtap_core_data)
        );
endmodule
 
 
                               
                               
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
	
   
    
 
   
 
   
 
       
       
       
       
 
 
  
  
  
  
  
  
  
 
 
 
  
 
  
  
  
  
   
    
 
 
 
 
 
 
 
 
module config_regs(
   input wire clk,
   input wire rst_n,
   input wire l15_config_req_val_s2,
   input wire l15_config_req_rw_s2,
   input wire [63:0] l15_config_write_req_data_s2,
   input wire [15:8] l15_config_req_address_s2,
   input wire [14-1:0] default_chipid,
   input wire [8-1:0] default_coreid_x,
   input wire [8-1:0] default_coreid_y,
input wire [6-1:0] from_dmbr_cred_bin_0,
input wire [6-1:0] from_dmbr_cred_bin_1,
input wire [6-1:0] from_dmbr_cred_bin_2,
input wire [6-1:0] from_dmbr_cred_bin_3,
input wire [6-1:0] from_dmbr_cred_bin_4,
input wire [6-1:0] from_dmbr_cred_bin_5,
input wire [6-1:0] from_dmbr_cred_bin_6,
input wire [6-1:0] from_dmbr_cred_bin_7,
input wire [6-1:0] from_dmbr_cred_bin_8,
input wire [6-1:0] from_dmbr_cred_bin_9,
   output wire [63:0] config_l15_read_res_data_s3,
   output wire [22-1:0] config_hmt_base,
   output wire                         config_dmbr_func_en,
   output wire                         config_dmbr_stall_en,
   output wire                         config_dmbr_proc_ld,
   output wire [16-1:0]  config_dmbr_replenish_cycles,
   output wire [10-1:0]      config_dmbr_bin_scale,
output wire [6-1:0] config_dmbr_cred_bin_0,
output wire [6-1:0] config_dmbr_cred_bin_1,
output wire [6-1:0] config_dmbr_cred_bin_2,
output wire [6-1:0] config_dmbr_cred_bin_3,
output wire [6-1:0] config_dmbr_cred_bin_4,
output wire [6-1:0] config_dmbr_cred_bin_5,
output wire [6-1:0] config_dmbr_cred_bin_6,
output wire [6-1:0] config_dmbr_cred_bin_7,
output wire [6-1:0] config_dmbr_cred_bin_8,
output wire [6-1:0] config_dmbr_cred_bin_9,
   output wire config_csm_en,
   output wire [31:0] config_system_tile_count,
   output wire [2-1:0] config_home_alloc_method,
   output wire [14-1:0] config_chipid,
   output wire [8-1:0] config_coreid_x,
   output wire [8-1:0] config_coreid_y,
   
   input wire rtap_config_req_val,
   input wire rtap_config_req_rw,
   input wire [63:0] rtap_config_write_req_data,
   input wire [15:8] rtap_config_req_address,
   output wire [63:0] config_rtap_read_res_data
);
reg [63:0] read_data_s3;
reg [63:0] read_data_s3_next;
reg                        dmbr_func_en            , dmbr_func_en_next;
reg                        dmbr_stall_en           , dmbr_stall_en_next;
reg                        dmbr_proc_ld            , dmbr_proc_ld_next;
reg                        dmbr_rd_cur_val         , dmbr_rd_cur_val_next;
reg [16-1:0] dmbr_replenish_cycles   , dmbr_replenish_cycles_next;
reg [10-1:0]     dmbr_bin_scale          , dmbr_bin_scale_next;
reg [6-1:0] dmbr_cred_bin_0, dmbr_cred_bin_0_next;
reg [6-1:0] dmbr_cred_bin_1, dmbr_cred_bin_1_next;
reg [6-1:0] dmbr_cred_bin_2, dmbr_cred_bin_2_next;
reg [6-1:0] dmbr_cred_bin_3, dmbr_cred_bin_3_next;
reg [6-1:0] dmbr_cred_bin_4, dmbr_cred_bin_4_next;
reg [6-1:0] dmbr_cred_bin_5, dmbr_cred_bin_5_next;
reg [6-1:0] dmbr_cred_bin_6, dmbr_cred_bin_6_next;
reg [6-1:0] dmbr_cred_bin_7, dmbr_cred_bin_7_next;
reg [6-1:0] dmbr_cred_bin_8, dmbr_cred_bin_8_next;
reg [6-1:0] dmbr_cred_bin_9, dmbr_cred_bin_9_next;
reg csm_en;
reg [22-1:0] hmt_base;
reg [31:0] system_tile_count;
reg [2-1:0]  home_alloc_method;
reg csm_en_next;
reg [31:0] system_tile_count_next;
reg [22-1:0] hmt_base_next;
reg [2-1:0]  home_alloc_method_next;
reg [14-1:0] chipid;
reg [8-1:0] coreid_x;
reg [8-1:0] coreid_y;
reg [14-1:0] chipid_next;
reg [8-1:0] coreid_x_next;
reg [8-1:0] coreid_y_next;
assign config_l15_read_res_data_s3 = read_data_s3;
assign config_rtap_read_res_data = read_data_s3; 
assign config_dmbr_func_en = dmbr_func_en;
assign config_dmbr_stall_en = dmbr_stall_en;
assign config_dmbr_proc_ld = dmbr_proc_ld;
assign config_dmbr_replenish_cycles = dmbr_replenish_cycles;
assign config_dmbr_bin_scale = dmbr_bin_scale;
assign config_dmbr_cred_bin_0 = dmbr_cred_bin_0;
assign config_dmbr_cred_bin_1 = dmbr_cred_bin_1;
assign config_dmbr_cred_bin_2 = dmbr_cred_bin_2;
assign config_dmbr_cred_bin_3 = dmbr_cred_bin_3;
assign config_dmbr_cred_bin_4 = dmbr_cred_bin_4;
assign config_dmbr_cred_bin_5 = dmbr_cred_bin_5;
assign config_dmbr_cred_bin_6 = dmbr_cred_bin_6;
assign config_dmbr_cred_bin_7 = dmbr_cred_bin_7;
assign config_dmbr_cred_bin_8 = dmbr_cred_bin_8;
assign config_dmbr_cred_bin_9 = dmbr_cred_bin_9;
assign config_hmt_base = hmt_base;
   assign config_csm_en = csm_en;
assign config_system_tile_count = system_tile_count;
assign config_home_alloc_method = home_alloc_method;
assign config_chipid = chipid;
assign config_coreid_x = coreid_x;
assign config_coreid_y = coreid_y;
localparam default_total_num_tile = 1;
always @ (posedge clk)
begin
   if (!rst_n)
   begin
      read_data_s3 <= 0;
      dmbr_func_en            <= 1'b0;
      dmbr_stall_en           <= 1'b0;
      dmbr_proc_ld            <= 1'b0;
      dmbr_replenish_cycles   <= {16{1'b0}};
      dmbr_bin_scale          <= {10{1'b0}};
      dmbr_cred_bin_0 <= {6{1'b0}};
dmbr_cred_bin_1 <= {6{1'b0}};
dmbr_cred_bin_2 <= {6{1'b0}};
dmbr_cred_bin_3 <= {6{1'b0}};
dmbr_cred_bin_4 <= {6{1'b0}};
dmbr_cred_bin_5 <= {6{1'b0}};
dmbr_cred_bin_6 <= {6{1'b0}};
dmbr_cred_bin_7 <= {6{1'b0}};
dmbr_cred_bin_8 <= {6{1'b0}};
dmbr_cred_bin_9 <= {6{1'b0}};
      dmbr_rd_cur_val <= 1'b0;
      hmt_base <= 22'b0;
      csm_en <= 1'b0;
      system_tile_count <= default_total_num_tile;
      home_alloc_method <= 2'd3;
      chipid <= default_chipid;
      coreid_x <= default_coreid_x;
      coreid_y <= default_coreid_y;
   end
   else
   begin
      read_data_s3 <= read_data_s3_next;
      dmbr_func_en <= dmbr_func_en_next;
      dmbr_stall_en <= dmbr_stall_en_next;
      dmbr_proc_ld <= dmbr_proc_ld_next;
      dmbr_replenish_cycles <= dmbr_replenish_cycles_next;
      dmbr_bin_scale <= dmbr_bin_scale_next;
      dmbr_cred_bin_0 <= dmbr_cred_bin_0_next;
dmbr_cred_bin_1 <= dmbr_cred_bin_1_next;
dmbr_cred_bin_2 <= dmbr_cred_bin_2_next;
dmbr_cred_bin_3 <= dmbr_cred_bin_3_next;
dmbr_cred_bin_4 <= dmbr_cred_bin_4_next;
dmbr_cred_bin_5 <= dmbr_cred_bin_5_next;
dmbr_cred_bin_6 <= dmbr_cred_bin_6_next;
dmbr_cred_bin_7 <= dmbr_cred_bin_7_next;
dmbr_cred_bin_8 <= dmbr_cred_bin_8_next;
dmbr_cred_bin_9 <= dmbr_cred_bin_9_next;
      dmbr_rd_cur_val <= dmbr_rd_cur_val_next;
      hmt_base <= hmt_base_next;
      csm_en <= csm_en_next;
      system_tile_count <= system_tile_count_next;
      home_alloc_method <= home_alloc_method_next;
      chipid <= chipid_next;
      coreid_x <= coreid_x_next;
      coreid_y <= coreid_y_next;
   end
end
reg req_val;
reg req_rw;
reg [63:0] req_data;
reg [15:8] req_address;
always @ *
begin
   req_val = rtap_config_req_val || l15_config_req_val_s2;
   req_rw = l15_config_req_rw_s2;
   req_data = l15_config_write_req_data_s2;
   req_address = l15_config_req_address_s2;
   if (rtap_config_req_val)
   begin
      req_rw = rtap_config_req_rw;
      req_data = rtap_config_write_req_data;
      req_address = rtap_config_req_address;
   end
end
always @ *
begin
   dmbr_func_en_next = dmbr_func_en;
   dmbr_stall_en_next = dmbr_stall_en;
   dmbr_proc_ld_next = dmbr_proc_ld;
   dmbr_replenish_cycles_next = dmbr_replenish_cycles;
   dmbr_bin_scale_next = dmbr_bin_scale;
   dmbr_cred_bin_0_next = dmbr_cred_bin_0;
dmbr_cred_bin_1_next = dmbr_cred_bin_1;
dmbr_cred_bin_2_next = dmbr_cred_bin_2;
dmbr_cred_bin_3_next = dmbr_cred_bin_3;
dmbr_cred_bin_4_next = dmbr_cred_bin_4;
dmbr_cred_bin_5_next = dmbr_cred_bin_5;
dmbr_cred_bin_6_next = dmbr_cred_bin_6;
dmbr_cred_bin_7_next = dmbr_cred_bin_7;
dmbr_cred_bin_8_next = dmbr_cred_bin_8;
dmbr_cred_bin_9_next = dmbr_cred_bin_9;
   dmbr_rd_cur_val_next = dmbr_rd_cur_val;
   hmt_base_next = hmt_base;
   csm_en_next = csm_en;
   system_tile_count_next = system_tile_count;
   home_alloc_method_next = home_alloc_method;
   chipid_next = chipid;
   coreid_x_next = coreid_x;
   coreid_y_next = coreid_y;
   if (req_val && req_rw == 1'b1)
   begin
      case (req_address[15:8])
         8'd0:
         begin
            {chipid_next, coreid_y_next, coreid_x_next} = req_data;
         end
         8'd1:
         begin
            csm_en_next = req_data[0];
         end
         8'd2:
         begin
            dmbr_func_en_next    = req_data[8'h0];
            dmbr_stall_en_next   = req_data[8'h1];
            dmbr_proc_ld_next    = req_data[8'h2];
            dmbr_rd_cur_val_next = req_data[8'h3];
            dmbr_cred_bin_0_next = req_data[9:4];
dmbr_cred_bin_1_next = req_data[15:10];
dmbr_cred_bin_2_next = req_data[21:16];
dmbr_cred_bin_3_next = req_data[27:22];
dmbr_cred_bin_4_next = req_data[33:28];
dmbr_cred_bin_5_next = req_data[39:34];
dmbr_cred_bin_6_next = req_data[45:40];
dmbr_cred_bin_7_next = req_data[51:46];
dmbr_cred_bin_8_next = req_data[57:52];
dmbr_cred_bin_9_next = req_data[63:58];
         end
         8'd5:
         begin
            dmbr_replenish_cycles_next = req_data[15:0];
            dmbr_bin_scale_next        = req_data[25:16];
         end
         8'd3:
         begin
            hmt_base_next = req_data[22-1:0];
         end
         8'd4:
         begin
            system_tile_count_next = req_data[31:0];
         end
         8'd6:
         begin
            home_alloc_method_next = req_data[2-1:0];
         end
      endcase
   end
end
always @ *
begin
   read_data_s3_next = read_data_s3;
   if (req_val && req_rw == 1'b0)
   begin
      case (req_address[15:8])
         8'd0:
         begin
               read_data_s3_next = {chipid, coreid_y, coreid_x};
         end
         8'd1:
         begin
               read_data_s3_next = config_csm_en;
         end
         8'd2:
         begin
            read_data_s3_next[3:0] = {dmbr_rd_cur_val, dmbr_proc_ld, dmbr_stall_en, dmbr_func_en};
            if (dmbr_rd_cur_val)
            begin
            read_data_s3_next[9:4] = from_dmbr_cred_bin_0;
read_data_s3_next[15:10] = from_dmbr_cred_bin_1;
read_data_s3_next[21:16] = from_dmbr_cred_bin_2;
read_data_s3_next[27:22] = from_dmbr_cred_bin_3;
read_data_s3_next[33:28] = from_dmbr_cred_bin_4;
read_data_s3_next[39:34] = from_dmbr_cred_bin_5;
read_data_s3_next[45:40] = from_dmbr_cred_bin_6;
read_data_s3_next[51:46] = from_dmbr_cred_bin_7;
read_data_s3_next[57:52] = from_dmbr_cred_bin_8;
read_data_s3_next[63:58] = from_dmbr_cred_bin_9;
            end
            else
            begin
            read_data_s3_next[9:4] = dmbr_cred_bin_0;
read_data_s3_next[15:10] = dmbr_cred_bin_1;
read_data_s3_next[21:16] = dmbr_cred_bin_2;
read_data_s3_next[27:22] = dmbr_cred_bin_3;
read_data_s3_next[33:28] = dmbr_cred_bin_4;
read_data_s3_next[39:34] = dmbr_cred_bin_5;
read_data_s3_next[45:40] = dmbr_cred_bin_6;
read_data_s3_next[51:46] = dmbr_cred_bin_7;
read_data_s3_next[57:52] = dmbr_cred_bin_8;
read_data_s3_next[63:58] = dmbr_cred_bin_9;
            end
         end
         8'd5:
         begin
            read_data_s3_next = {{64-16-10{1'b0}}, {dmbr_bin_scale, dmbr_replenish_cycles}};
         end
         8'd3:
         begin
            read_data_s3_next = config_hmt_base;
         end
         8'd4:
         begin
            read_data_s3_next = system_tile_count;
         end
         8'd6:
         begin
            read_data_s3_next = home_alloc_method;
         end
      endcase
   end
end
endmodule
module OCI (
   
   input slew,
   input impsel1,
   input impsel2,
   input core_ref_clk,
   input io_clk,
   input rst_n,
   input pll_rst_n,
   input [4:0] pll_rangea,
   input [1:0] clk_mux_sel,
   input clk_en,
   input pll_bypass,
   input async_mux,
   input oram_on,
   input oram_traffic_gen,
   input oram_dummy_gen,
   output pll_lock,
   input  wire jtag_clk,
   input  wire jtag_rst_l,
   input  wire jtag_modesel,
   input  wire jtag_datain,
   output wire jtag_dataout,
   input  [31:0]                 intf_chip_data,
   input  [1:0]                  intf_chip_channel,
   output [2:0]                  intf_chip_credit_back,
   output [31:0]                 chip_intf_data,
   output [1:0]                  chip_intf_channel,
   input  [2:0]                  chip_intf_credit_back,
   
   output core_ref_clk_inter,
   output io_clk_inter,
   output rst_n_inter,
   output pll_rst_n_inter,
   output [4:0] pll_rangea_inter,
   output [1:0] clk_mux_sel_inter,
   output clk_en_inter,
   output pll_bypass_inter,
   output async_mux_inter,
   output oram_on_inter,
   output oram_traffic_gen_inter,
   output oram_dummy_gen_inter,
   input  pll_lock_inter,
   output wire jtag_clk_inter,
   output wire jtag_rst_l_inter,
   output wire jtag_modesel_inter,
   output wire jtag_datain_inter,
   input  wire jtag_dataout_inter,
   output [31:0]                 intf_chip_data_inter,
   output [1:0]                  intf_chip_channel_inter,
   input  [2:0]                  intf_chip_credit_back_inter,
   input  [31:0]                 chip_intf_data_inter,
   input  [1:0]                  chip_intf_channel_inter,
   output [2:0]                  chip_intf_credit_back_inter
   );
    assign core_ref_clk_inter = core_ref_clk;
    assign io_clk_inter = io_clk;
    assign rst_n_inter = rst_n;
    assign pll_rst_n_inter = pll_rst_n;
    assign pll_rangea_inter = pll_rangea;
    assign clk_mux_sel_inter = clk_mux_sel;
    assign clk_en_inter = clk_en;
    assign pll_bypass_inter = pll_bypass;
    assign async_mux_inter = async_mux;
    assign oram_on_inter = oram_on;
    assign oram_traffic_gen_inter = oram_traffic_gen;
    assign oram_dummy_gen_inter = oram_dummy_gen;
    assign pll_lock = pll_lock_inter;
    assign jtag_clk_inter = jtag_clk;
    assign jtag_rst_l_inter = jtag_rst_l;
    assign jtag_modesel_inter = jtag_modesel;
    assign jtag_datain_inter = jtag_datain;
    assign jtag_dataout = jtag_dataout_inter;
    assign intf_chip_data_inter = intf_chip_data;
    assign intf_chip_channel_inter = intf_chip_channel;
    assign intf_chip_credit_back = intf_chip_credit_back_inter;
    assign chip_intf_data = chip_intf_data_inter;
    assign chip_intf_channel = chip_intf_channel_inter;
    assign chip_intf_credit_back_inter = chip_intf_credit_back;
 
   
   endmodule
   
 
    
    
 
    
    
    
    
    
    
 
 
 
  
    
 
 
    
    
    
    
    
    
    
 
 
  
          
      
    
         
module chip(
   
   input                                        slew,
   input                                        impsel1,
   input                                        impsel2,
 
 
   
   input                                        core_ref_clk,
   input                                        io_clk,
 
   
   
   input                                        rst_n,
   input                                        pll_rst_n,
   
   input                                        clk_en,
   
   output                                       pll_lock,
   input                                        pll_bypass,
   input  [4:0]                                 pll_rangea,
   
   
   input  [1:0]                                 clk_mux_sel,
   
   input                                        jtag_clk,
   input                                        jtag_rst_l,
   input                                        jtag_modesel,
   input                                        jtag_datain,
   output                                       jtag_dataout,
   
   input                                        async_mux,
   
   input                                        oram_on,
   input                                        oram_traffic_gen,
   input                                        oram_dummy_gen,
 
   
 
   
   input  [31:0]                                intf_chip_data,
   input  [1:0]                                 intf_chip_channel,
   output [2:0]                                 intf_chip_credit_back,
   output [31:0]                                chip_intf_data,
   output [1:0]                                 chip_intf_channel,
   input  [2:0]                                 chip_intf_credit_back
 
 
    ,
    
    input                                       ndmreset_i,    
    input   [1-1:0]                    debug_req_i,   
    output  [1-1:0]                    unavailable_o, 
    
    input   [1-1:0]                    timer_irq_i,   
    input   [1-1:0]                    ipi_i,         
    
    input   [1*2-1:0]                  irq_i          
);
   
   
   
   
   
 
   
 
   
 
 
   
   wire                                         core_ref_clk_inter;
   wire                                         io_clk_inter;
   wire                                         rst_n_inter;
   wire                                         pll_rst_n_inter;
   wire                                         clk_en_inter;
   wire                                         pll_lock_inter;
   wire                                         pll_bypass_inter;
   wire [4:0]                                   pll_rangea_inter;
   wire [1:0]                                   clk_mux_sel_inter;
   wire                                         jtag_clk_inter;
   wire                                         jtag_rst_l_inter;
   wire                                         jtag_rst_l_inter_sync;
   wire                                         jtag_modesel_inter;
   wire                                         jtag_datain_inter;
   wire                                         jtag_dataout_inter;
   wire                                         async_mux_inter;
   wire                                         oram_on_inter;
   wire                                         oram_traffic_gen_inter;
   wire                                         oram_dummy_gen_inter;
   wire [31:0]                              intf_chip_data_inter;
   wire [1:0]                                   intf_chip_channel_inter;
   wire [2:0]                                   intf_chip_credit_back_inter;
   wire [31:0]                                  chip_intf_data_inter;
   wire [1:0]                                   chip_intf_channel_inter;
   wire [2:0]                                   chip_intf_credit_back_inter;
   
   wire                                         rst_n_inter_sync;
   reg                                          rst_n_inter_sync_f;
   wire                                         io_clk_rst_n_inter_sync;
   reg                                          io_clk_rst_n_inter_sync_f;
   
   wire                                         core_ref_clk_inter_c;
   wire                                         core_ref_clk_inter_t;
   wire                                         clk_muxed;
   wire                                         pll_clk;
   
   reg  [31:0]                                  intf_chip_data_inter_buf_f ;
   reg  [1:0]                                   intf_chip_channel_inter_buf_f ;
   reg  [2:0]                                   chip_intf_credit_back_inter_buf_f ;
   
   wire                                         chip_intf_noc1_valid;
   wire [64-1:0]                   chip_intf_noc1_data;
   wire                                         chip_intf_noc1_rdy;
   wire                                         chip_intf_noc2_valid;
   wire [64-1:0]                   chip_intf_noc2_data;
   wire                                         chip_intf_noc2_rdy;
   wire                                         chip_intf_noc3_valid;
   wire [64-1:0]                   chip_intf_noc3_data;
   wire                                         chip_intf_noc3_rdy;
   wire                                         intf_chip_noc1_valid;
   wire [64-1:0]                   intf_chip_noc1_data;
   wire                                         intf_chip_noc1_rdy;
   wire                                         intf_chip_noc2_valid;
   wire [64-1:0]                   intf_chip_noc2_data;
   wire                                         intf_chip_noc2_rdy;
   wire                                         intf_chip_noc3_valid;
   wire [64-1:0]                   intf_chip_noc3_data;
   wire                                         intf_chip_noc3_rdy;
   
   
   wire                                         processor_offchip_noc1_valid;
   wire [64-1:0]                   processor_offchip_noc1_data;
   wire                                         processor_offchip_noc1_yummy;
   wire                                         processor_offchip_noc2_valid;
   wire [64-1:0]                   processor_offchip_noc2_data;
   wire                                         processor_offchip_noc2_yummy;
   wire                                         processor_offchip_noc3_valid;
   wire [64-1:0]                   processor_offchip_noc3_data;
   wire                                         processor_offchip_noc3_yummy;
   wire                                         offchip_processor_noc1_valid;
   wire [64-1:0]                   offchip_processor_noc1_data;
   wire                                         offchip_processor_noc1_yummy;
   wire                                         offchip_processor_noc2_valid;
   wire [64-1:0]                   offchip_processor_noc2_data;
   wire                                         offchip_processor_noc2_yummy;
   wire                                         offchip_processor_noc3_valid;
   wire [64-1:0]                   offchip_processor_noc3_data;
   wire                                         offchip_processor_noc3_yummy;
 
   
   reg                                          proc_oram_yummy;
   reg                                          oram_proc_valid;
   reg  [64-1:0]                   oram_proc_data;
   reg                                          offchip_oram_yummy;
   reg                                          oram_offchip_valid;
   reg  [64-1:0]                   oram_offchip_data;
   
   wire                                         proc_oram_valid;
   wire [64-1:0]                   proc_oram_data;
   wire                                         proc_oram_yummy_oram;
   wire                                         oram_proc_valid_oram;
   wire [64-1:0]                   oram_proc_data_oram;
   wire                                         oram_proc_yummy;
   wire                                         offchip_oram_valid;
   wire [64-1:0]                   offchip_oram_data;
   wire                                         offchip_oram_yummy_oram;
   wire                                         oram_offchip_valid_oram;
   wire [64-1:0]                   oram_offchip_data_oram;
   wire                                         oram_offchip_yummy;
   
   wire                                         ctap_oram_clk_en;
   wire                                         ctap_oram_req_val;
   wire [4-1:0]             ctap_oram_req_misc;
   wire [64-1:0]             oram_ctap_res_data;
   
   
   
   
   wire                                         tiles_jtag_ucb_val;
   wire [4-1:0]                    tiles_jtag_ucb_data;
   
   wire                                         jtag_tiles_ucb_val;
   wire [4-1:0]                    jtag_tiles_ucb_data;
   wire [127:0]                                 ctap_clk_en_inter; 
   wire tile0_jtag_ucb_val;
wire [4-1:0] tile0_jtag_ucb_data;
   
wire [64-1:0] tile_0_0_out_N_noc1_data;
wire [64-1:0] tile_0_0_out_S_noc1_data;
wire [64-1:0] tile_0_0_out_E_noc1_data;
wire [64-1:0] tile_0_0_out_W_noc1_data;
wire tile_0_0_out_N_noc1_valid;
wire tile_0_0_out_S_noc1_valid;
wire tile_0_0_out_E_noc1_valid;
wire tile_0_0_out_W_noc1_valid;
wire tile_0_0_out_N_noc1_yummy;
wire tile_0_0_out_S_noc1_yummy;
wire tile_0_0_out_E_noc1_yummy;
wire tile_0_0_out_W_noc1_yummy;
wire [64-1:0] tile_0_0_out_N_noc2_data;
wire [64-1:0] tile_0_0_out_S_noc2_data;
wire [64-1:0] tile_0_0_out_E_noc2_data;
wire [64-1:0] tile_0_0_out_W_noc2_data;
wire tile_0_0_out_N_noc2_valid;
wire tile_0_0_out_S_noc2_valid;
wire tile_0_0_out_E_noc2_valid;
wire tile_0_0_out_W_noc2_valid;
wire tile_0_0_out_N_noc2_yummy;
wire tile_0_0_out_S_noc2_yummy;
wire tile_0_0_out_E_noc2_yummy;
wire tile_0_0_out_W_noc2_yummy;
wire [64-1:0] tile_0_0_out_N_noc3_data;
wire [64-1:0] tile_0_0_out_S_noc3_data;
wire [64-1:0] tile_0_0_out_E_noc3_data;
wire [64-1:0] tile_0_0_out_W_noc3_data;
wire tile_0_0_out_N_noc3_valid;
wire tile_0_0_out_S_noc3_valid;
wire tile_0_0_out_E_noc3_valid;
wire tile_0_0_out_W_noc3_valid;
wire tile_0_0_out_N_noc3_yummy;
wire tile_0_0_out_S_noc3_yummy;
wire tile_0_0_out_E_noc3_yummy;
wire tile_0_0_out_W_noc3_yummy;
wire [64-1:0] dummy_out_N_noc1_data = 64'b0;
wire [64-1:0] dummy_out_S_noc1_data = 64'b0;
wire [64-1:0] dummy_out_E_noc1_data = 64'b0;
wire [64-1:0] dummy_out_W_noc1_data = 64'b0;
wire dummy_out_N_noc1_valid = 1'b0;
wire dummy_out_S_noc1_valid = 1'b0;
wire dummy_out_E_noc1_valid = 1'b0;
wire dummy_out_W_noc1_valid = 1'b0;
wire dummy_out_N_noc1_yummy = 1'b0;
wire dummy_out_S_noc1_yummy = 1'b0;
wire dummy_out_E_noc1_yummy = 1'b0;
wire dummy_out_W_noc1_yummy = 1'b0;
wire [64-1:0] dummy_out_N_noc2_data = 64'b0;
wire [64-1:0] dummy_out_S_noc2_data = 64'b0;
wire [64-1:0] dummy_out_E_noc2_data = 64'b0;
wire [64-1:0] dummy_out_W_noc2_data = 64'b0;
wire dummy_out_N_noc2_valid = 1'b0;
wire dummy_out_S_noc2_valid = 1'b0;
wire dummy_out_E_noc2_valid = 1'b0;
wire dummy_out_W_noc2_valid = 1'b0;
wire dummy_out_N_noc2_yummy = 1'b0;
wire dummy_out_S_noc2_yummy = 1'b0;
wire dummy_out_E_noc2_yummy = 1'b0;
wire dummy_out_W_noc2_yummy = 1'b0;
wire [64-1:0] dummy_out_N_noc3_data = 64'b0;
wire [64-1:0] dummy_out_S_noc3_data = 64'b0;
wire [64-1:0] dummy_out_E_noc3_data = 64'b0;
wire [64-1:0] dummy_out_W_noc3_data = 64'b0;
wire dummy_out_N_noc3_valid = 1'b0;
wire dummy_out_S_noc3_valid = 1'b0;
wire dummy_out_E_noc3_valid = 1'b0;
wire dummy_out_W_noc3_valid = 1'b0;
wire dummy_out_N_noc3_yummy = 1'b0;
wire dummy_out_S_noc3_yummy = 1'b0;
wire dummy_out_E_noc3_yummy = 1'b0;
wire dummy_out_W_noc3_yummy = 1'b0;
wire [64-1:0] offchip_out_E_noc1_data;
wire offchip_out_E_noc1_valid;
wire offchip_out_E_noc1_yummy;
wire [64-1:0] offchip_out_E_noc2_data;
wire offchip_out_E_noc2_valid;
wire offchip_out_E_noc2_yummy;
wire [64-1:0] offchip_out_E_noc3_data;
wire offchip_out_E_noc3_valid;
wire offchip_out_E_noc3_yummy;
   
   
   
   
   
   
   always @ (posedge clk_muxed)
      rst_n_inter_sync_f <= rst_n_inter_sync;
   always @ (posedge io_clk_inter)
      io_clk_rst_n_inter_sync_f <= io_clk_rst_n_inter_sync;
   
   always @(posedge io_clk_inter)
   begin
 
       if(~rst_n_inter_sync_f)
       begin
           intf_chip_data_inter_buf_f <= 0;
           intf_chip_channel_inter_buf_f <= 0;
           chip_intf_credit_back_inter_buf_f <= 0;
       end
       else
       begin
           intf_chip_data_inter_buf_f <= intf_chip_data_inter;
           intf_chip_channel_inter_buf_f <= intf_chip_channel_inter;
           chip_intf_credit_back_inter_buf_f <= chip_intf_credit_back_inter;
       end
   end
 
   
   
   
   
   
 
   
assign proc_oram_valid = tile_0_0_out_W_noc2_valid;
assign proc_oram_data = tile_0_0_out_W_noc2_data;
assign oram_proc_yummy = tile_0_0_out_W_noc3_yummy;
   assign offchip_oram_valid = offchip_processor_noc3_valid;
   assign offchip_oram_data = offchip_processor_noc3_data;
   assign oram_offchip_yummy = processor_offchip_noc2_yummy;
assign processor_offchip_noc1_valid = tile_0_0_out_W_noc1_valid;
assign processor_offchip_noc1_data = tile_0_0_out_W_noc1_data;
assign offchip_processor_noc1_yummy = tile_0_0_out_W_noc1_yummy;
   assign processor_offchip_noc2_valid = oram_offchip_valid;
   assign processor_offchip_noc2_data = oram_offchip_data;
assign offchip_processor_noc2_yummy = tile_0_0_out_W_noc2_yummy;
assign processor_offchip_noc3_valid = tile_0_0_out_W_noc3_valid;
assign processor_offchip_noc3_data = tile_0_0_out_W_noc3_data;
   assign offchip_processor_noc3_yummy = offchip_oram_yummy;
assign offchip_out_E_noc1_data = offchip_processor_noc1_data;
assign offchip_out_E_noc1_valid = offchip_processor_noc1_valid;
assign offchip_out_E_noc1_yummy = processor_offchip_noc1_yummy;
assign offchip_out_E_noc2_data = offchip_processor_noc2_data;
assign offchip_out_E_noc2_valid = offchip_processor_noc2_valid;
assign offchip_out_E_noc2_yummy = proc_oram_yummy; 
assign offchip_out_E_noc3_data = oram_proc_data;
assign offchip_out_E_noc3_valid = oram_proc_valid;
assign offchip_out_E_noc3_yummy = processor_offchip_noc3_yummy;
   
   always @ *
   begin
     
     oram_offchip_valid = proc_oram_valid;
     oram_offchip_data = proc_oram_data;
     proc_oram_yummy = oram_offchip_yummy;
     oram_proc_valid = offchip_oram_valid;
     oram_proc_data = offchip_oram_data;
     offchip_oram_yummy = oram_proc_yummy;
     if (oram_on_inter)
     begin
       oram_offchip_valid = oram_offchip_valid_oram;
       oram_offchip_data = oram_offchip_data_oram;
       proc_oram_yummy = proc_oram_yummy_oram;
       oram_proc_valid = oram_proc_valid_oram;
       oram_proc_data = oram_proc_data_oram;
       offchip_oram_yummy = offchip_oram_yummy_oram;
     end
   end
   
assign tiles_jtag_ucb_val = tile0_jtag_ucb_val;
assign tiles_jtag_ucb_data = tile0_jtag_ucb_data;
   
   
   
   
 
 
 
   
   OCI oci_inst (
   
   .slew                (slew),
   .impsel1                (impsel1),
   .impsel2                (impsel2),
   .core_ref_clk           (core_ref_clk),
   .io_clk                 (io_clk),
   .rst_n                  (rst_n),
   .pll_rst_n              (pll_rst_n),
   .pll_rangea             (pll_rangea),
   .clk_mux_sel               (clk_mux_sel),
   .clk_en                 (clk_en),
   .pll_bypass             (pll_bypass),
   .async_mux              (async_mux),
   .oram_on                (oram_on),
   .oram_traffic_gen       (oram_traffic_gen),
   .oram_dummy_gen            (oram_dummy_gen),
   .pll_lock               (pll_lock),
   .jtag_clk               (jtag_clk),
   .jtag_rst_l             (jtag_rst_l),
   .jtag_modesel           (jtag_modesel),
   .jtag_datain               (jtag_datain),
   .jtag_dataout           (jtag_dataout),
   .intf_chip_data            (intf_chip_data),
   .intf_chip_channel         (intf_chip_channel),
   .intf_chip_credit_back     (intf_chip_credit_back),
   .chip_intf_data            (chip_intf_data),
   .chip_intf_channel         (chip_intf_channel),
   .chip_intf_credit_back     (chip_intf_credit_back),
 
   
   .core_ref_clk_inter        (core_ref_clk_inter),
   .io_clk_inter           (io_clk_inter),
   .rst_n_inter               (rst_n_inter),
   .pll_rst_n_inter           (pll_rst_n_inter),
   .pll_rangea_inter       (pll_rangea_inter),
   .clk_mux_sel_inter         (clk_mux_sel_inter),
   .clk_en_inter           (clk_en_inter),
   .pll_bypass_inter       (pll_bypass_inter),
   .async_mux_inter           (async_mux_inter),
   .oram_on_inter          (oram_on_inter),
   .oram_traffic_gen_inter    (oram_traffic_gen_inter),
   .oram_dummy_gen_inter      (oram_dummy_gen_inter),
   .pll_lock_inter            (pll_lock_inter),
   .jtag_clk_inter            (jtag_clk_inter),
   .jtag_rst_l_inter       (jtag_rst_l_inter),
   .jtag_modesel_inter        (jtag_modesel_inter),
   .jtag_datain_inter         (jtag_datain_inter),
   .jtag_dataout_inter        (jtag_dataout_inter),
   .intf_chip_data_inter      (intf_chip_data_inter),
   .intf_chip_channel_inter      (intf_chip_channel_inter),
   .intf_chip_credit_back_inter  (intf_chip_credit_back_inter),
   .chip_intf_data_inter      (chip_intf_data_inter),
   .chip_intf_channel_inter      (chip_intf_channel_inter),
   .chip_intf_credit_back_inter  (chip_intf_credit_back_inter) );
   
   clk_se_to_diff ref_clk_converter (
       .clk_se  (core_ref_clk_inter),
       .clk_p   (core_ref_clk_inter_t),
       .clk_n   (core_ref_clk_inter_c)
   );
   clk_mux clock_mux (
       .clk0_p(core_ref_clk_inter_t),
       .clk0_n(core_ref_clk_inter_c),
       .clk1_p(1'b1),
       .clk1_n(1'b0),
       .clk2(pll_clk),
       .sel(clk_mux_sel_inter),
       .clk_muxed(clk_muxed)
   );
   pll_top pll_top (
      .clk_locked(pll_lock_inter),
      .clk_out(pll_clk),
      .rangeA(pll_rangea_inter),
      .bypass_en(pll_bypass_inter),
      .ref_clk(core_ref_clk_inter),
      .rst(~pll_rst_n_inter)
   );
   
   
   
   
   
   synchronizer rst_sync (
      .clk(clk_muxed),
      .presyncdata(rst_n_inter),
      .syncdata(rst_n_inter_sync)
   );
   synchronizer io_clk_rst_sync (
      .clk(io_clk_inter),
      .presyncdata(rst_n_inter),
      .syncdata(io_clk_rst_n_inter_sync)
   );
   synchronizer jtag_rst_sync (
      .clk(clk_muxed),
      .presyncdata(jtag_rst_l_inter),
      .syncdata(jtag_rst_l_inter_sync)
   );
   
   chip_bridge chip_intf(
       
       
 
       .rst_n                  (rst_n_inter_sync_f),
       .chip_clk               (clk_muxed),
       .intcnct_clk            (io_clk_inter),
       .async_mux              (async_mux_inter),
       .network_out_1          (chip_intf_noc1_data),
       .network_out_2          (chip_intf_noc2_data),
       .network_out_3          (chip_intf_noc3_data),
       .data_out_val_1         (chip_intf_noc1_valid),
       .data_out_val_2         (chip_intf_noc2_valid),
       .data_out_val_3         (chip_intf_noc3_valid),
       .data_out_rdy_1         (chip_intf_noc1_rdy),
       .data_out_rdy_2         (chip_intf_noc2_rdy),
       .data_out_rdy_3         (chip_intf_noc3_rdy),
       .intcnct_data_in        (intf_chip_data_inter_buf_f),
       .intcnct_channel_in     (intf_chip_channel_inter_buf_f),
       .intcnct_credit_back_in (intf_chip_credit_back_inter),
       .network_in_1           (intf_chip_noc1_data),
       .network_in_2           (intf_chip_noc2_data),
       .network_in_3           (intf_chip_noc3_data),
       .data_in_val_1          (intf_chip_noc1_valid),
       .data_in_val_2          (intf_chip_noc2_valid),
       .data_in_val_3          (intf_chip_noc3_valid),
       .data_in_rdy_1          (intf_chip_noc1_rdy),
       .data_in_rdy_2          (intf_chip_noc2_rdy),
       .data_in_rdy_3          (intf_chip_noc3_rdy),
       .intcnct_data_out       (chip_intf_data_inter),
       .intcnct_channel_out    (chip_intf_channel_inter),
       .intcnct_credit_back_out(chip_intf_credit_back_inter_buf_f)
   );
   
   valrdy_to_credit #(4, 3) chip_from_intf_noc1_v2c(
      .clk(clk_muxed),
      .reset(~rst_n_inter_sync_f),
      .data_in(intf_chip_noc1_data),
      .valid_in(intf_chip_noc1_valid),
      .ready_in(intf_chip_noc1_rdy),
      .data_out(offchip_processor_noc1_data),           
      .valid_out(offchip_processor_noc1_valid),       
      .yummy_out(offchip_processor_noc1_yummy)    
   );
   credit_to_valrdy chip_to_intf_noc1_c2v(
      .clk(clk_muxed),
      .reset(~rst_n_inter_sync_f),
      .data_in(processor_offchip_noc1_data),
      .valid_in(processor_offchip_noc1_valid),
      .yummy_in(processor_offchip_noc1_yummy),
      .data_out(chip_intf_noc1_data),           
      .valid_out(chip_intf_noc1_valid),       
      .ready_out(chip_intf_noc1_rdy)    
   );
   valrdy_to_credit #(4, 3) chip_from_intf_noc2_v2c(
      .clk(clk_muxed),
      .reset(~rst_n_inter_sync_f),
      .data_in(intf_chip_noc2_data),
      .valid_in(intf_chip_noc2_valid),
      .ready_in(intf_chip_noc2_rdy),
      .data_out(offchip_processor_noc2_data),           
      .valid_out(offchip_processor_noc2_valid),       
      .yummy_out(offchip_processor_noc2_yummy)    
   );
   credit_to_valrdy chip_to_intf_noc2_c2v(
      .clk(clk_muxed),
      .reset(~rst_n_inter_sync_f),
      .data_in(processor_offchip_noc2_data),
      .valid_in(processor_offchip_noc2_valid),
      .yummy_in(processor_offchip_noc2_yummy),
      .data_out(chip_intf_noc2_data),           
      .valid_out(chip_intf_noc2_valid),       
      .ready_out(chip_intf_noc2_rdy)    
   );
   valrdy_to_credit #(4, 3) chip_from_intf_noc3_v2c(
      .clk(clk_muxed),
      .reset(~rst_n_inter_sync_f),
      .data_in(intf_chip_noc3_data),
      .valid_in(intf_chip_noc3_valid),
      .ready_in(intf_chip_noc3_rdy),
      .data_out(offchip_processor_noc3_data),           
      .valid_out(offchip_processor_noc3_valid),       
      .yummy_out(offchip_processor_noc3_yummy)    
   );
   credit_to_valrdy chip_to_intf_noc3_c2v(
      .clk(clk_muxed),
      .reset(~rst_n_inter_sync_f),
      .data_in(processor_offchip_noc3_data),
      .valid_in(processor_offchip_noc3_valid),
      .yummy_in(processor_offchip_noc3_yummy),
      .data_out(chip_intf_noc3_data),           
      .valid_out(chip_intf_noc3_valid),       
      .ready_out(chip_intf_noc3_rdy)    
   );
 
 
   
   jtag jtag_port(
      .clk(clk_muxed),
      .rst_n(rst_n_inter_sync_f),
      .jtag_clk(jtag_clk_inter),
      .jtag_rst_l(jtag_rst_l_inter_sync),
      .jtag_modesel(jtag_modesel_inter),
      .jtag_datain(jtag_datain_inter),
      .jtag_dataout(jtag_dataout_inter),
      .jtag_dataout_en(),
      .jtag_tiles_ucb_val(jtag_tiles_ucb_val),
      .jtag_tiles_ucb_data(jtag_tiles_ucb_data),
      .tiles_jtag_ucb_val(tiles_jtag_ucb_val),
      .tiles_jtag_ucb_data(tiles_jtag_ucb_data),
      .ctap_oram_req_val(ctap_oram_req_val),
      .ctap_oram_req_misc(ctap_oram_req_misc),
      .oram_ctap_res_data(oram_ctap_res_data),
      
      
      
      .ctap_clk_en(ctap_clk_en_inter),
      .ctap_oram_clk_en(ctap_oram_clk_en)
   );
   
    
tile #(.TILE_TYPE(0))
tile0 (
    .clk                (clk_muxed),
    .rst_n              (rst_n_inter_sync),
    .clk_en             (ctap_clk_en_inter[0] && clk_en_inter),
    .default_chipid             (14'b0),    
    .default_coreid_x           (8'd0),
    .default_coreid_y           (8'd0),
    .flat_tileid                (8'd0),
    .debug_req_i         ( debug_req_i[0]   ),
    .unavailable_o       ( unavailable_o[0] ),
    .timer_irq_i         ( timer_irq_i[0]   ),
    .ipi_i               ( ipi_i[0]         ),
    .irq_i               ( irq_i[0*2 +: 2]  ),
    
    .tile_jtag_ucb_val   ( tile0_jtag_ucb_val      ),
    .tile_jtag_ucb_data  ( tile0_jtag_ucb_data     ),
    
    .jtag_tiles_ucb_val  ( jtag_tiles_ucb_val      ),
    .jtag_tiles_ucb_data ( jtag_tiles_ucb_data     ),
    .dyn0_dataIn_N       ( dummy_out_S_noc1_data   ),
    .dyn0_dataIn_E       ( dummy_out_W_noc1_data   ),
    .dyn0_dataIn_W       ( offchip_out_E_noc1_data   ),
    .dyn0_dataIn_S       ( dummy_out_N_noc1_data   ),
    .dyn0_validIn_N      ( dummy_out_S_noc1_valid  ),
    .dyn0_validIn_E      ( dummy_out_W_noc1_valid  ),
    .dyn0_validIn_W      ( offchip_out_E_noc1_valid  ),
    .dyn0_validIn_S      ( dummy_out_N_noc1_valid  ),
    .dyn0_dNo_yummy      ( dummy_out_S_noc1_yummy  ),
    .dyn0_dEo_yummy      ( dummy_out_W_noc1_yummy  ),
    .dyn0_dWo_yummy      ( offchip_out_E_noc1_yummy  ),
    .dyn0_dSo_yummy      ( dummy_out_N_noc1_yummy  ),
    .dyn0_dNo            ( tile_0_0_out_N_noc1_data  ),
    .dyn0_dEo            ( tile_0_0_out_E_noc1_data  ),
    .dyn0_dWo            ( tile_0_0_out_W_noc1_data  ),
    .dyn0_dSo            ( tile_0_0_out_S_noc1_data  ),
    .dyn0_dNo_valid      ( tile_0_0_out_N_noc1_valid ),
    .dyn0_dEo_valid      ( tile_0_0_out_E_noc1_valid ),
    .dyn0_dWo_valid      ( tile_0_0_out_W_noc1_valid ),
    .dyn0_dSo_valid      ( tile_0_0_out_S_noc1_valid ),
    .dyn0_yummyOut_N     ( tile_0_0_out_N_noc1_yummy ),
    .dyn0_yummyOut_E     ( tile_0_0_out_E_noc1_yummy ),
    .dyn0_yummyOut_W     ( tile_0_0_out_W_noc1_yummy ),
    .dyn0_yummyOut_S     ( tile_0_0_out_S_noc1_yummy ),
    .dyn1_dataIn_N       ( dummy_out_S_noc2_data   ),
    .dyn1_dataIn_E       ( dummy_out_W_noc2_data   ),
    .dyn1_dataIn_W       ( offchip_out_E_noc2_data   ),
    .dyn1_dataIn_S       ( dummy_out_N_noc2_data   ),
    .dyn1_validIn_N      ( dummy_out_S_noc2_valid  ),
    .dyn1_validIn_E      ( dummy_out_W_noc2_valid  ),
    .dyn1_validIn_W      ( offchip_out_E_noc2_valid  ),
    .dyn1_validIn_S      ( dummy_out_N_noc2_valid  ),
    .dyn1_dNo_yummy      ( dummy_out_S_noc2_yummy  ),
    .dyn1_dEo_yummy      ( dummy_out_W_noc2_yummy  ),
    .dyn1_dWo_yummy      ( offchip_out_E_noc2_yummy  ),
    .dyn1_dSo_yummy      ( dummy_out_N_noc2_yummy  ),
    .dyn1_dNo            ( tile_0_0_out_N_noc2_data  ),
    .dyn1_dEo            ( tile_0_0_out_E_noc2_data  ),
    .dyn1_dWo            ( tile_0_0_out_W_noc2_data  ),
    .dyn1_dSo            ( tile_0_0_out_S_noc2_data  ),
    .dyn1_dNo_valid      ( tile_0_0_out_N_noc2_valid ),
    .dyn1_dEo_valid      ( tile_0_0_out_E_noc2_valid ),
    .dyn1_dWo_valid      ( tile_0_0_out_W_noc2_valid ),
    .dyn1_dSo_valid      ( tile_0_0_out_S_noc2_valid ),
    .dyn1_yummyOut_N     ( tile_0_0_out_N_noc2_yummy ),
    .dyn1_yummyOut_E     ( tile_0_0_out_E_noc2_yummy ),
    .dyn1_yummyOut_W     ( tile_0_0_out_W_noc2_yummy ),
    .dyn1_yummyOut_S     ( tile_0_0_out_S_noc2_yummy ),
    .dyn2_dataIn_N       ( dummy_out_S_noc3_data   ),
    .dyn2_dataIn_E       ( dummy_out_W_noc3_data   ),
    .dyn2_dataIn_W       ( offchip_out_E_noc3_data   ),
    .dyn2_dataIn_S       ( dummy_out_N_noc3_data   ),
    .dyn2_validIn_N      ( dummy_out_S_noc3_valid  ),
    .dyn2_validIn_E      ( dummy_out_W_noc3_valid  ),
    .dyn2_validIn_W      ( offchip_out_E_noc3_valid  ),
    .dyn2_validIn_S      ( dummy_out_N_noc3_valid  ),
    .dyn2_dNo_yummy      ( dummy_out_S_noc3_yummy  ),
    .dyn2_dEo_yummy      ( dummy_out_W_noc3_yummy  ),
    .dyn2_dWo_yummy      ( offchip_out_E_noc3_yummy  ),
    .dyn2_dSo_yummy      ( dummy_out_N_noc3_yummy  ),
    .dyn2_dNo            ( tile_0_0_out_N_noc3_data  ),
    .dyn2_dEo            ( tile_0_0_out_E_noc3_data  ),
    .dyn2_dWo            ( tile_0_0_out_W_noc3_data  ),
    .dyn2_dSo            ( tile_0_0_out_S_noc3_data  ),
    .dyn2_dNo_valid      ( tile_0_0_out_N_noc3_valid ),
    .dyn2_dEo_valid      ( tile_0_0_out_E_noc3_valid ),
    .dyn2_dWo_valid      ( tile_0_0_out_W_noc3_valid ),
    .dyn2_dSo_valid      ( tile_0_0_out_S_noc3_valid ),
    .dyn2_yummyOut_N     ( tile_0_0_out_N_noc3_yummy ),
    .dyn2_yummyOut_E     ( tile_0_0_out_E_noc3_yummy ),
    .dyn2_yummyOut_W     ( tile_0_0_out_W_noc3_yummy ),
    .dyn2_yummyOut_S     ( tile_0_0_out_S_noc3_yummy )
);
endmodule
    
    
 
    
    
    
    
    
    
 
 
 
  
    
 
 
    
    
    
    
    
    
    
 
 
module OpenPitonRV64(
 
    
 
 
 
 
 
 
 
 
 
 
 
 
    input sys_clk,
    input                                       sys_rst_n,
 
    
 
    
 
    
 
    
  
 
 
 
  
 
 
 
    
    
 
 
    
    
    
    
    
    
    
     
    
    
    
     
    
    
 
    input                                        mc_clk,
    
    output wire [6     -1:0]    m_axi_awid,
    output wire [64   -1:0]    m_axi_awaddr,
    output wire [8    -1:0]    m_axi_awlen,
    output wire [3   -1:0]    m_axi_awsize,
    output wire [2  -1:0]    m_axi_awburst,
    output wire                                  m_axi_awlock,
    output wire [4  -1:0]    m_axi_awcache,
    output wire [3   -1:0]    m_axi_awprot,
    output wire [4    -1:0]    m_axi_awqos,
    output wire [4 -1:0]    m_axi_awregion,
    output wire [11   -1:0]    m_axi_awuser,
    output wire                                  m_axi_awvalid,
    input  wire                                  m_axi_awready,
    
    output wire  [6     -1:0]    m_axi_wid,
    output wire  [512   -1:0]    m_axi_wdata,
    output wire  [64   -1:0]    m_axi_wstrb,
    output wire                                   m_axi_wlast,
    output wire  [11   -1:0]    m_axi_wuser,
    output wire                                   m_axi_wvalid,
    input  wire                                   m_axi_wready,
    
    output wire  [6     -1:0]    m_axi_arid,
    output wire  [64   -1:0]    m_axi_araddr,
    output wire  [8    -1:0]    m_axi_arlen,
    output wire  [3   -1:0]    m_axi_arsize,
    output wire  [2  -1:0]    m_axi_arburst,
    output wire                                   m_axi_arlock,
    output wire  [4  -1:0]    m_axi_arcache,
    output wire  [3   -1:0]    m_axi_arprot,
    output wire  [4    -1:0]    m_axi_arqos,
    output wire  [4 -1:0]    m_axi_arregion,
    output wire  [11   -1:0]    m_axi_aruser,
    output wire                                   m_axi_arvalid,
    input  wire                                   m_axi_arready,
    
    input  wire  [6     -1:0]    m_axi_rid,
    input  wire  [512   -1:0]    m_axi_rdata,
    input  wire  [2   -1:0]    m_axi_rresp,
    input  wire                                   m_axi_rlast,
    input  wire  [11   -1:0]    m_axi_ruser,
    input  wire                                   m_axi_rvalid,
    output wire                                   m_axi_rready,
    
    input  wire  [6     -1:0]    m_axi_bid,
    input  wire  [2   -1:0]    m_axi_bresp,
    input  wire  [11   -1:0]    m_axi_buser,
    input  wire                                   m_axi_bvalid,
    output wire                                   m_axi_bready,
    input  wire                                   ddr_ready,
 
 
 
 
 
    
    
    
    
    
    
 
    
    
    
    
 
 
    
 
 
 
    input [31:0]                                       ext_irq,
    input [31:0]                                      ext_irq_trigger
 
);
wire                core_ref_clk;
wire                io_clk;
 
wire                io_clk_loopback;
reg                 sys_rst_n_rect;
reg                 chip_rst_n;
reg                 jtag_rst_n_full;
reg                 pll_rst_n_full;
reg                 passthru_rst_n;
wire                passthru_chip_rst_n;
wire                passthru_jtag_rst_n;
wire                passthru_pll_rst_n;
reg                 chipset_rst_n;
wire                pll_lock;
 
wire                piton_prsnt_n;
wire                piton_ready_n;
wire [31:0]         intf_chip_data;
wire [1:0]          intf_chip_channel;
wire [2:0]          intf_chip_credit_back;
wire [31:0]         chip_intf_data;
wire [1:0]          chip_intf_channel;
wire [2:0]          chip_intf_credit_back;
wire                         processor_offchip_noc1_valid;
wire [64-1:0]   processor_offchip_noc1_data;
wire                         processor_offchip_noc1_yummy;
wire                         processor_offchip_noc2_valid;
wire [64-1:0]   processor_offchip_noc2_data;
wire                         processor_offchip_noc2_yummy;
wire                         processor_offchip_noc3_valid;
wire [64-1:0]   processor_offchip_noc3_data;
wire                         processor_offchip_noc3_yummy;
wire                         offchip_processor_noc1_valid;
wire [64-1:0]   offchip_processor_noc1_data;
wire                         offchip_processor_noc1_yummy;
wire                         offchip_processor_noc2_valid;
wire [64-1:0]   offchip_processor_noc2_data;
wire                         offchip_processor_noc2_yummy;
wire                         offchip_processor_noc3_valid;
wire [64-1:0]   offchip_processor_noc3_data;
wire                         offchip_processor_noc3_yummy;
 
 
wire [31:0]         chipset_passthru_data_p;
wire [31:0]         chipset_passthru_data_n;
wire [1:0]          chipset_passthru_channel_p;
wire [1:0]          chipset_passthru_channel_n;
wire [2:0]          chipset_passthru_credit_back_p;
wire [2:0]          chipset_passthru_credit_back_n;
wire [31:0]         passthru_chipset_data_p;
wire [31:0]         passthru_chipset_data_n;
wire [1:0]          passthru_chipset_channel_p;
wire [1:0]          passthru_chipset_channel_n;
wire [2:0]          passthru_chipset_credit_back_p;
wire [2:0]          passthru_chipset_credit_back_n;
wire                     ndmreset;    
wire                     dmactive;    
wire  [1-1:0]   debug_req;   
wire  [1-1:0]   unavailable; 
wire                     rtc;         
wire  [1-1:0]   timer_irq;   
wire  [1-1:0]   ipi;         
wire  [1*2-1:0] irq;         
 
 
reg [6:0] rtc_div;
always @(posedge core_ref_clk or negedge chip_rst_n) begin : p_rtc_div
  if(~chip_rst_n) begin
    rtc_div <= 7'h0;
  end else begin
    rtc_div <= rtc_div + 7'h1;
  end
end
assign rtc = rtc_div[6];
 
always @ *
begin
 
    sys_rst_n_rect = sys_rst_n;
end
always @ *
begin
    chip_rst_n = sys_rst_n_rect & passthru_chip_rst_n;
    jtag_rst_n_full = passthru_jtag_rst_n;
 
    pll_rst_n_full = passthru_pll_rst_n;
 
    
    
    passthru_rst_n = sys_rst_n_rect;
    
    
    
    
    
    
    chipset_rst_n = sys_rst_n;
end
assign passthru_chip_rst_n = 1'b1;
assign passthru_jtag_rst_n = 1'b1;
assign passthru_pll_rst_n = 1'b1;
chip chip(
    
    
    .slew (1'b1),
    .impsel1(1'b1),
    .impsel2(1'b1),
 
    
    .core_ref_clk(core_ref_clk),
    .io_clk(io_clk),
    .rst_n(chip_rst_n),
    .pll_rst_n(pll_rst_n_full),
    
    
    .clk_en(1'b1),
    
    .pll_lock (pll_lock),
    
    .pll_bypass (1'b1),
    .pll_rangea (5'b0),
 
    
    
    
    .clk_mux_sel (2'b0),
 
    
    
    .jtag_clk(1'b0),
    .jtag_rst_l(1'b1),
    .jtag_modesel(1'b1),
    .jtag_datain(1'b0),
    .jtag_dataout(),
 
    
    
 
    
    .async_mux (1'b1),
 
 
    
    .intf_chip_data(intf_chip_data),
    .intf_chip_channel(intf_chip_channel),
    .intf_chip_credit_back(intf_chip_credit_back),
    
    .chip_intf_data(chip_intf_data),
    .chip_intf_channel(chip_intf_channel),
    .chip_intf_credit_back(chip_intf_credit_back)
 
    ,
    
    .ndmreset_i                     ( ndmreset                   ), 
    .debug_req_i                    ( debug_req                  ), 
    .unavailable_o                  ( unavailable                ), 
    
    .timer_irq_i                    ( timer_irq                  ), 
    .ipi_i                          ( ipi                        ), 
    
    .irq_i                          ( irq                        )  
);
    
    
    
 
 
chipset chipset(
    
    
    .sys_clk(sys_clk),
 
 
 
 
 
 
 
 
 
    .io_clk(io_clk),
 
 
 
    
    .rst_n(chipset_rst_n),
    
    
    
    
    
 
    .piton_prsnt_n(1'b0),
    .piton_ready_n(1'b0),
 
    
    
    
    
 
    
    .intf_chip_data(intf_chip_data),
    .intf_chip_channel(intf_chip_channel),
    .intf_chip_credit_back(intf_chip_credit_back),
    .chip_intf_data(chip_intf_data),
    .chip_intf_channel(chip_intf_channel),
    .chip_intf_credit_back(chip_intf_credit_back),
 
    
 
 
    .mc_clk(mc_clk),
    
    .m_axi_awid(m_axi_awid),
    .m_axi_awaddr(m_axi_awaddr),
    .m_axi_awlen(m_axi_awlen),
    .m_axi_awsize(m_axi_awsize),
    .m_axi_awburst(m_axi_awburst),
    .m_axi_awlock(m_axi_awlock),
    .m_axi_awcache(m_axi_awcache),
    .m_axi_awprot(m_axi_awprot),
    .m_axi_awqos(m_axi_awqos),
    .m_axi_awregion(m_axi_awregion),
    .m_axi_awuser(m_axi_awuser),
    .m_axi_awvalid(m_axi_awvalid),
    .m_axi_awready(m_axi_awready),
    
    .m_axi_wid(m_axi_wid),
    .m_axi_wdata(m_axi_wdata),
    .m_axi_wstrb(m_axi_wstrb),
    .m_axi_wlast(m_axi_wlast),
    .m_axi_wuser(m_axi_wuser),
    .m_axi_wvalid(m_axi_wvalid),
    .m_axi_wready(m_axi_wready),
    
    .m_axi_arid(m_axi_arid),
    .m_axi_araddr(m_axi_araddr),
    .m_axi_arlen(m_axi_arlen),
    .m_axi_arsize(m_axi_arsize),
    .m_axi_arburst(m_axi_arburst),
    .m_axi_arlock(m_axi_arlock),
    .m_axi_arcache(m_axi_arcache),
    .m_axi_arprot(m_axi_arprot),
    .m_axi_arqos(m_axi_arqos),
    .m_axi_arregion(m_axi_arregion),
    .m_axi_aruser(m_axi_aruser),
    .m_axi_arvalid(m_axi_arvalid),
    .m_axi_arready(m_axi_arready),
    
    .m_axi_rid(m_axi_rid),
    .m_axi_rdata(m_axi_rdata),
    .m_axi_rresp(m_axi_rresp),
    .m_axi_rlast(m_axi_rlast),
    .m_axi_ruser(m_axi_ruser),
    .m_axi_rvalid(m_axi_rvalid),
    .m_axi_rready(m_axi_rready),
    
    .m_axi_bid(m_axi_bid),
    .m_axi_bresp(m_axi_bresp),
    .m_axi_buser(m_axi_buser),
    .m_axi_bvalid(m_axi_bvalid),
    .m_axi_bready(m_axi_bready),
    .ddr_ready(ddr_ready),
 
 
 
 
 
    
    
    
    
    
    
 
    
     
 
    .ext_irq(ext_irq),
    .ext_irq_trigger(ext_irq_trigger)
    ,
    
    .ndmreset_o                     ( ndmreset                   ), 
    .dmactive_o                     ( dmactive                   ), 
    .debug_req_o                    ( debug_req                  ), 
    .unavailable_i                  ( unavailable                ), 
    
    .tck_i                          ( tck_i                      ),
    .tms_i                          ( tms_i                      ),
    .trst_ni                        ( trst_ni                    ),
    .td_i                           ( td_i                       ),
    .td_o                           ( td_o                       ),
    .tdo_oe_o                       (                            ),
    
    .rtc_i                          ( rtc                        ), 
    .timer_irq_o                    ( timer_irq                  ), 
    .ipi_o                          ( ipi                        ), 
    
    .irq_o                          ( irq                        )  
);
endmodule


